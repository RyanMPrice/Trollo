magic
tech gf180mcuC
magscale 1 10
timestamp 1670260711
<< metal1 >>
rect 1344 60394 59024 60428
rect 1344 60342 4478 60394
rect 4530 60342 4582 60394
rect 4634 60342 4686 60394
rect 4738 60342 35198 60394
rect 35250 60342 35302 60394
rect 35354 60342 35406 60394
rect 35458 60342 59024 60394
rect 1344 60308 59024 60342
rect 22878 60226 22930 60238
rect 21970 60174 21982 60226
rect 22034 60223 22046 60226
rect 22530 60223 22542 60226
rect 22034 60177 22542 60223
rect 22034 60174 22046 60177
rect 22530 60174 22542 60177
rect 22594 60174 22606 60226
rect 22878 60162 22930 60174
rect 10434 60062 10446 60114
rect 10498 60062 10510 60114
rect 31042 60062 31054 60114
rect 31106 60062 31118 60114
rect 51090 60062 51102 60114
rect 51154 60062 51166 60114
rect 4622 60002 4674 60014
rect 4622 59938 4674 59950
rect 9774 60002 9826 60014
rect 14590 60002 14642 60014
rect 11330 59950 11342 60002
rect 11394 59950 11406 60002
rect 9774 59938 9826 59950
rect 14590 59938 14642 59950
rect 23326 60002 23378 60014
rect 23326 59938 23378 59950
rect 23550 60002 23602 60014
rect 30370 59950 30382 60002
rect 30434 59950 30446 60002
rect 33954 59950 33966 60002
rect 34018 59950 34030 60002
rect 50418 59950 50430 60002
rect 50482 59950 50494 60002
rect 23550 59938 23602 59950
rect 5070 59890 5122 59902
rect 5070 59826 5122 59838
rect 6302 59890 6354 59902
rect 6302 59826 6354 59838
rect 14702 59890 14754 59902
rect 14702 59826 14754 59838
rect 15038 59890 15090 59902
rect 15038 59826 15090 59838
rect 22766 59890 22818 59902
rect 22766 59826 22818 59838
rect 22990 59890 23042 59902
rect 22990 59826 23042 59838
rect 26910 59890 26962 59902
rect 26910 59826 26962 59838
rect 33630 59890 33682 59902
rect 33630 59826 33682 59838
rect 43710 59890 43762 59902
rect 43710 59826 43762 59838
rect 3726 59778 3778 59790
rect 3726 59714 3778 59726
rect 4174 59778 4226 59790
rect 4174 59714 4226 59726
rect 5854 59778 5906 59790
rect 5854 59714 5906 59726
rect 6750 59778 6802 59790
rect 6750 59714 6802 59726
rect 7198 59778 7250 59790
rect 7198 59714 7250 59726
rect 7646 59778 7698 59790
rect 7646 59714 7698 59726
rect 8094 59778 8146 59790
rect 8094 59714 8146 59726
rect 8542 59778 8594 59790
rect 8542 59714 8594 59726
rect 8990 59778 9042 59790
rect 8990 59714 9042 59726
rect 12350 59778 12402 59790
rect 12350 59714 12402 59726
rect 12910 59778 12962 59790
rect 12910 59714 12962 59726
rect 13582 59778 13634 59790
rect 13582 59714 13634 59726
rect 14030 59778 14082 59790
rect 14030 59714 14082 59726
rect 14926 59778 14978 59790
rect 14926 59714 14978 59726
rect 15710 59778 15762 59790
rect 15710 59714 15762 59726
rect 16158 59778 16210 59790
rect 16158 59714 16210 59726
rect 16606 59778 16658 59790
rect 16606 59714 16658 59726
rect 17614 59778 17666 59790
rect 17614 59714 17666 59726
rect 18062 59778 18114 59790
rect 18062 59714 18114 59726
rect 18734 59778 18786 59790
rect 18734 59714 18786 59726
rect 19182 59778 19234 59790
rect 19182 59714 19234 59726
rect 19742 59778 19794 59790
rect 19742 59714 19794 59726
rect 20190 59778 20242 59790
rect 20190 59714 20242 59726
rect 20638 59778 20690 59790
rect 20638 59714 20690 59726
rect 21422 59778 21474 59790
rect 21422 59714 21474 59726
rect 21870 59778 21922 59790
rect 21870 59714 21922 59726
rect 22318 59778 22370 59790
rect 22318 59714 22370 59726
rect 24222 59778 24274 59790
rect 24222 59714 24274 59726
rect 24558 59778 24610 59790
rect 24558 59714 24610 59726
rect 25230 59778 25282 59790
rect 25230 59714 25282 59726
rect 27022 59778 27074 59790
rect 27022 59714 27074 59726
rect 29822 59778 29874 59790
rect 29822 59714 29874 59726
rect 33182 59778 33234 59790
rect 33182 59714 33234 59726
rect 33742 59778 33794 59790
rect 33742 59714 33794 59726
rect 34750 59778 34802 59790
rect 34750 59714 34802 59726
rect 35534 59778 35586 59790
rect 35534 59714 35586 59726
rect 42926 59778 42978 59790
rect 42926 59714 42978 59726
rect 43822 59778 43874 59790
rect 43822 59714 43874 59726
rect 44942 59778 44994 59790
rect 44942 59714 44994 59726
rect 49870 59778 49922 59790
rect 49870 59714 49922 59726
rect 1344 59610 59024 59644
rect 1344 59558 19838 59610
rect 19890 59558 19942 59610
rect 19994 59558 20046 59610
rect 20098 59558 50558 59610
rect 50610 59558 50662 59610
rect 50714 59558 50766 59610
rect 50818 59558 59024 59610
rect 1344 59524 59024 59558
rect 4622 59442 4674 59454
rect 4622 59378 4674 59390
rect 8990 59442 9042 59454
rect 8990 59378 9042 59390
rect 10110 59442 10162 59454
rect 10110 59378 10162 59390
rect 11006 59442 11058 59454
rect 11006 59378 11058 59390
rect 12798 59442 12850 59454
rect 12798 59378 12850 59390
rect 15934 59442 15986 59454
rect 15934 59378 15986 59390
rect 17950 59442 18002 59454
rect 17950 59378 18002 59390
rect 24894 59442 24946 59454
rect 24894 59378 24946 59390
rect 25678 59442 25730 59454
rect 25678 59378 25730 59390
rect 27918 59442 27970 59454
rect 27918 59378 27970 59390
rect 34190 59442 34242 59454
rect 34190 59378 34242 59390
rect 36990 59442 37042 59454
rect 36990 59378 37042 59390
rect 5070 59330 5122 59342
rect 5070 59266 5122 59278
rect 6414 59330 6466 59342
rect 6414 59266 6466 59278
rect 8654 59330 8706 59342
rect 8654 59266 8706 59278
rect 10670 59330 10722 59342
rect 10670 59266 10722 59278
rect 19518 59330 19570 59342
rect 19518 59266 19570 59278
rect 20078 59330 20130 59342
rect 20078 59266 20130 59278
rect 29934 59330 29986 59342
rect 29934 59266 29986 59278
rect 30158 59330 30210 59342
rect 30158 59266 30210 59278
rect 30718 59330 30770 59342
rect 30718 59266 30770 59278
rect 32622 59330 32674 59342
rect 32622 59266 32674 59278
rect 34414 59330 34466 59342
rect 34414 59266 34466 59278
rect 36430 59330 36482 59342
rect 36430 59266 36482 59278
rect 38222 59330 38274 59342
rect 38222 59266 38274 59278
rect 42030 59330 42082 59342
rect 42030 59266 42082 59278
rect 42254 59330 42306 59342
rect 42254 59266 42306 59278
rect 45502 59330 45554 59342
rect 45502 59266 45554 59278
rect 14590 59218 14642 59230
rect 14354 59166 14366 59218
rect 14418 59166 14430 59218
rect 14590 59154 14642 59166
rect 14702 59218 14754 59230
rect 20302 59218 20354 59230
rect 19058 59166 19070 59218
rect 19122 59166 19134 59218
rect 14702 59154 14754 59166
rect 20302 59154 20354 59166
rect 20526 59218 20578 59230
rect 28030 59218 28082 59230
rect 21746 59166 21758 59218
rect 21810 59166 21822 59218
rect 23874 59166 23886 59218
rect 23938 59166 23950 59218
rect 24098 59166 24110 59218
rect 24162 59166 24174 59218
rect 24322 59166 24334 59218
rect 24386 59166 24398 59218
rect 26674 59166 26686 59218
rect 26738 59166 26750 59218
rect 20526 59154 20578 59166
rect 28030 59154 28082 59166
rect 28142 59218 28194 59230
rect 28142 59154 28194 59166
rect 29822 59218 29874 59230
rect 29822 59154 29874 59166
rect 30830 59218 30882 59230
rect 30830 59154 30882 59166
rect 32510 59218 32562 59230
rect 32510 59154 32562 59166
rect 32846 59218 32898 59230
rect 35198 59218 35250 59230
rect 33954 59166 33966 59218
rect 34018 59166 34030 59218
rect 32846 59154 32898 59166
rect 35198 59154 35250 59166
rect 36318 59218 36370 59230
rect 36318 59154 36370 59166
rect 36654 59218 36706 59230
rect 36654 59154 36706 59166
rect 38110 59218 38162 59230
rect 38110 59154 38162 59166
rect 38446 59218 38498 59230
rect 38446 59154 38498 59166
rect 40574 59218 40626 59230
rect 40574 59154 40626 59166
rect 41470 59218 41522 59230
rect 41470 59154 41522 59166
rect 42702 59218 42754 59230
rect 42702 59154 42754 59166
rect 43038 59218 43090 59230
rect 43038 59154 43090 59166
rect 43486 59218 43538 59230
rect 43486 59154 43538 59166
rect 43710 59218 43762 59230
rect 43710 59154 43762 59166
rect 44270 59218 44322 59230
rect 44270 59154 44322 59166
rect 44494 59218 44546 59230
rect 44494 59154 44546 59166
rect 44942 59218 44994 59230
rect 44942 59154 44994 59166
rect 45390 59218 45442 59230
rect 45390 59154 45442 59166
rect 2718 59106 2770 59118
rect 2718 59042 2770 59054
rect 3278 59106 3330 59118
rect 3278 59042 3330 59054
rect 3614 59106 3666 59118
rect 3614 59042 3666 59054
rect 4174 59106 4226 59118
rect 4174 59042 4226 59054
rect 5406 59106 5458 59118
rect 5406 59042 5458 59054
rect 5966 59106 6018 59118
rect 5966 59042 6018 59054
rect 6862 59106 6914 59118
rect 6862 59042 6914 59054
rect 7310 59106 7362 59118
rect 7310 59042 7362 59054
rect 7758 59106 7810 59118
rect 7758 59042 7810 59054
rect 8094 59106 8146 59118
rect 8094 59042 8146 59054
rect 9662 59106 9714 59118
rect 9662 59042 9714 59054
rect 11902 59106 11954 59118
rect 11902 59042 11954 59054
rect 12350 59106 12402 59118
rect 12350 59042 12402 59054
rect 13246 59106 13298 59118
rect 13246 59042 13298 59054
rect 13694 59106 13746 59118
rect 16606 59106 16658 59118
rect 16034 59054 16046 59106
rect 16098 59054 16110 59106
rect 13694 59042 13746 59054
rect 16606 59042 16658 59054
rect 17054 59106 17106 59118
rect 20190 59106 20242 59118
rect 27246 59106 27298 59118
rect 18610 59054 18622 59106
rect 18674 59054 18686 59106
rect 22082 59054 22094 59106
rect 22146 59054 22158 59106
rect 26786 59054 26798 59106
rect 26850 59054 26862 59106
rect 17054 59042 17106 59054
rect 20190 59042 20242 59054
rect 27246 59042 27298 59054
rect 28366 59106 28418 59118
rect 28366 59042 28418 59054
rect 29374 59106 29426 59118
rect 29374 59042 29426 59054
rect 31278 59106 31330 59118
rect 31278 59042 31330 59054
rect 39454 59106 39506 59118
rect 39454 59042 39506 59054
rect 42478 59106 42530 59118
rect 42478 59042 42530 59054
rect 43262 59106 43314 59118
rect 43262 59042 43314 59054
rect 44382 59106 44434 59118
rect 44382 59042 44434 59054
rect 45950 59106 46002 59118
rect 45950 59042 46002 59054
rect 15710 58994 15762 59006
rect 28590 58994 28642 59006
rect 15138 58942 15150 58994
rect 15202 58942 15214 58994
rect 22418 58942 22430 58994
rect 22482 58942 22494 58994
rect 23538 58942 23550 58994
rect 23602 58942 23614 58994
rect 15710 58930 15762 58942
rect 28590 58930 28642 58942
rect 30718 58994 30770 59006
rect 30718 58930 30770 58942
rect 34078 58994 34130 59006
rect 34078 58930 34130 58942
rect 35086 58994 35138 59006
rect 35086 58930 35138 58942
rect 35422 58994 35474 59006
rect 35422 58930 35474 58942
rect 35534 58994 35586 59006
rect 35534 58930 35586 58942
rect 38894 58994 38946 59006
rect 38894 58930 38946 58942
rect 39230 58994 39282 59006
rect 40350 58994 40402 59006
rect 40002 58942 40014 58994
rect 40066 58942 40078 58994
rect 39230 58930 39282 58942
rect 40350 58930 40402 58942
rect 1344 58826 59024 58860
rect 1344 58774 4478 58826
rect 4530 58774 4582 58826
rect 4634 58774 4686 58826
rect 4738 58774 35198 58826
rect 35250 58774 35302 58826
rect 35354 58774 35406 58826
rect 35458 58774 59024 58826
rect 1344 58740 59024 58774
rect 30158 58658 30210 58670
rect 11218 58606 11230 58658
rect 11282 58655 11294 58658
rect 11890 58655 11902 58658
rect 11282 58609 11902 58655
rect 11282 58606 11294 58609
rect 11890 58606 11902 58609
rect 11954 58606 11966 58658
rect 30158 58594 30210 58606
rect 37662 58658 37714 58670
rect 44382 58658 44434 58670
rect 40562 58606 40574 58658
rect 40626 58606 40638 58658
rect 37662 58594 37714 58606
rect 44382 58594 44434 58606
rect 12126 58546 12178 58558
rect 12126 58482 12178 58494
rect 16606 58546 16658 58558
rect 16606 58482 16658 58494
rect 18174 58546 18226 58558
rect 24558 58546 24610 58558
rect 19058 58494 19070 58546
rect 19122 58494 19134 58546
rect 22082 58494 22094 58546
rect 22146 58494 22158 58546
rect 18174 58482 18226 58494
rect 24558 58482 24610 58494
rect 27358 58546 27410 58558
rect 27358 58482 27410 58494
rect 28702 58546 28754 58558
rect 28702 58482 28754 58494
rect 29934 58546 29986 58558
rect 29934 58482 29986 58494
rect 32958 58546 33010 58558
rect 36766 58546 36818 58558
rect 36418 58494 36430 58546
rect 36482 58494 36494 58546
rect 32958 58482 33010 58494
rect 36766 58482 36818 58494
rect 41246 58546 41298 58558
rect 41246 58482 41298 58494
rect 42814 58546 42866 58558
rect 42814 58482 42866 58494
rect 46398 58546 46450 58558
rect 46398 58482 46450 58494
rect 47182 58546 47234 58558
rect 47182 58482 47234 58494
rect 50654 58546 50706 58558
rect 51202 58494 51214 58546
rect 51266 58494 51278 58546
rect 50654 58482 50706 58494
rect 13022 58434 13074 58446
rect 13022 58370 13074 58382
rect 13806 58434 13858 58446
rect 15150 58434 15202 58446
rect 18062 58434 18114 58446
rect 25454 58434 25506 58446
rect 26910 58434 26962 58446
rect 31502 58434 31554 58446
rect 33182 58434 33234 58446
rect 34750 58434 34802 58446
rect 14018 58382 14030 58434
rect 14082 58382 14094 58434
rect 16258 58382 16270 58434
rect 16322 58382 16334 58434
rect 17490 58382 17502 58434
rect 17554 58382 17566 58434
rect 19170 58382 19182 58434
rect 19234 58382 19246 58434
rect 22306 58382 22318 58434
rect 22370 58382 22382 58434
rect 23762 58382 23774 58434
rect 23826 58382 23838 58434
rect 24770 58382 24782 58434
rect 24834 58382 24846 58434
rect 25890 58382 25902 58434
rect 25954 58382 25966 58434
rect 30482 58382 30494 58434
rect 30546 58382 30558 58434
rect 32050 58382 32062 58434
rect 32114 58382 32126 58434
rect 33506 58382 33518 58434
rect 33570 58382 33582 58434
rect 34402 58382 34414 58434
rect 34466 58382 34478 58434
rect 13806 58370 13858 58382
rect 15150 58370 15202 58382
rect 18062 58370 18114 58382
rect 25454 58370 25506 58382
rect 26910 58370 26962 58382
rect 31502 58370 31554 58382
rect 33182 58370 33234 58382
rect 34750 58370 34802 58382
rect 34974 58434 35026 58446
rect 37550 58434 37602 58446
rect 36082 58382 36094 58434
rect 36146 58382 36158 58434
rect 34974 58370 35026 58382
rect 37550 58370 37602 58382
rect 38670 58434 38722 58446
rect 40014 58434 40066 58446
rect 44606 58434 44658 58446
rect 39106 58382 39118 58434
rect 39170 58382 39182 58434
rect 39442 58382 39454 58434
rect 39506 58382 39518 58434
rect 40562 58382 40574 58434
rect 40626 58382 40638 58434
rect 42018 58382 42030 58434
rect 42082 58382 42094 58434
rect 42354 58382 42366 58434
rect 42418 58382 42430 58434
rect 43474 58382 43486 58434
rect 43538 58382 43550 58434
rect 44146 58382 44158 58434
rect 44210 58382 44222 58434
rect 38670 58370 38722 58382
rect 40014 58370 40066 58382
rect 44606 58370 44658 58382
rect 46622 58434 46674 58446
rect 50430 58434 50482 58446
rect 47506 58382 47518 58434
rect 47570 58382 47582 58434
rect 50082 58382 50094 58434
rect 50146 58382 50158 58434
rect 46622 58370 46674 58382
rect 50430 58370 50482 58382
rect 7310 58322 7362 58334
rect 7310 58258 7362 58270
rect 9102 58322 9154 58334
rect 9102 58258 9154 58270
rect 9886 58322 9938 58334
rect 9886 58258 9938 58270
rect 12686 58322 12738 58334
rect 12686 58258 12738 58270
rect 14702 58322 14754 58334
rect 14702 58258 14754 58270
rect 15486 58322 15538 58334
rect 15486 58258 15538 58270
rect 19854 58322 19906 58334
rect 19854 58258 19906 58270
rect 22878 58322 22930 58334
rect 22878 58258 22930 58270
rect 23438 58322 23490 58334
rect 23438 58258 23490 58270
rect 24446 58322 24498 58334
rect 24446 58258 24498 58270
rect 26350 58322 26402 58334
rect 26350 58258 26402 58270
rect 27134 58322 27186 58334
rect 27134 58258 27186 58270
rect 27470 58322 27522 58334
rect 27470 58258 27522 58270
rect 28814 58322 28866 58334
rect 37662 58322 37714 58334
rect 51550 58322 51602 58334
rect 32274 58270 32286 58322
rect 32338 58270 32350 58322
rect 40226 58270 40238 58322
rect 40290 58270 40302 58322
rect 43138 58270 43150 58322
rect 43202 58270 43214 58322
rect 28814 58258 28866 58270
rect 37662 58258 37714 58270
rect 51550 58258 51602 58270
rect 1934 58210 1986 58222
rect 1934 58146 1986 58158
rect 2494 58210 2546 58222
rect 2494 58146 2546 58158
rect 2942 58210 2994 58222
rect 2942 58146 2994 58158
rect 3390 58210 3442 58222
rect 3390 58146 3442 58158
rect 3950 58210 4002 58222
rect 3950 58146 4002 58158
rect 4510 58210 4562 58222
rect 4510 58146 4562 58158
rect 4958 58210 5010 58222
rect 4958 58146 5010 58158
rect 5966 58210 6018 58222
rect 5966 58146 6018 58158
rect 6302 58210 6354 58222
rect 6302 58146 6354 58158
rect 6750 58210 6802 58222
rect 6750 58146 6802 58158
rect 7758 58210 7810 58222
rect 7758 58146 7810 58158
rect 8206 58210 8258 58222
rect 8206 58146 8258 58158
rect 8654 58210 8706 58222
rect 8654 58146 8706 58158
rect 9438 58210 9490 58222
rect 9438 58146 9490 58158
rect 10446 58210 10498 58222
rect 10446 58146 10498 58158
rect 10782 58210 10834 58222
rect 10782 58146 10834 58158
rect 11342 58210 11394 58222
rect 11342 58146 11394 58158
rect 11678 58210 11730 58222
rect 11678 58146 11730 58158
rect 12798 58210 12850 58222
rect 12798 58146 12850 58158
rect 15374 58210 15426 58222
rect 15374 58146 15426 58158
rect 16494 58210 16546 58222
rect 16494 58146 16546 58158
rect 20526 58210 20578 58222
rect 20526 58146 20578 58158
rect 20974 58210 21026 58222
rect 20974 58146 21026 58158
rect 23550 58210 23602 58222
rect 23550 58146 23602 58158
rect 28590 58210 28642 58222
rect 28590 58146 28642 58158
rect 31166 58210 31218 58222
rect 31166 58146 31218 58158
rect 34862 58210 34914 58222
rect 34862 58146 34914 58158
rect 38782 58210 38834 58222
rect 38782 58146 38834 58158
rect 38894 58210 38946 58222
rect 38894 58146 38946 58158
rect 40126 58210 40178 58222
rect 40126 58146 40178 58158
rect 44270 58210 44322 58222
rect 44270 58146 44322 58158
rect 45390 58210 45442 58222
rect 47294 58210 47346 58222
rect 46050 58158 46062 58210
rect 46114 58158 46126 58210
rect 45390 58146 45442 58158
rect 47294 58146 47346 58158
rect 51326 58210 51378 58222
rect 51326 58146 51378 58158
rect 1344 58042 59024 58076
rect 1344 57990 19838 58042
rect 19890 57990 19942 58042
rect 19994 57990 20046 58042
rect 20098 57990 50558 58042
rect 50610 57990 50662 58042
rect 50714 57990 50766 58042
rect 50818 57990 59024 58042
rect 1344 57956 59024 57990
rect 3166 57874 3218 57886
rect 3166 57810 3218 57822
rect 4062 57874 4114 57886
rect 4062 57810 4114 57822
rect 8990 57874 9042 57886
rect 8990 57810 9042 57822
rect 16382 57874 16434 57886
rect 27918 57874 27970 57886
rect 19282 57822 19294 57874
rect 19346 57822 19358 57874
rect 20402 57822 20414 57874
rect 20466 57822 20478 57874
rect 16382 57810 16434 57822
rect 27918 57810 27970 57822
rect 28142 57874 28194 57886
rect 28142 57810 28194 57822
rect 29486 57874 29538 57886
rect 29486 57810 29538 57822
rect 29822 57874 29874 57886
rect 29822 57810 29874 57822
rect 33742 57874 33794 57886
rect 33742 57810 33794 57822
rect 33966 57874 34018 57886
rect 33966 57810 34018 57822
rect 35646 57874 35698 57886
rect 35646 57810 35698 57822
rect 36430 57874 36482 57886
rect 36430 57810 36482 57822
rect 38110 57874 38162 57886
rect 38110 57810 38162 57822
rect 39678 57874 39730 57886
rect 39678 57810 39730 57822
rect 40462 57874 40514 57886
rect 43262 57874 43314 57886
rect 42130 57822 42142 57874
rect 42194 57822 42206 57874
rect 40462 57810 40514 57822
rect 43262 57810 43314 57822
rect 43486 57874 43538 57886
rect 43486 57810 43538 57822
rect 44158 57874 44210 57886
rect 44158 57810 44210 57822
rect 44494 57874 44546 57886
rect 44494 57810 44546 57822
rect 44606 57874 44658 57886
rect 44606 57810 44658 57822
rect 46734 57874 46786 57886
rect 46734 57810 46786 57822
rect 14366 57762 14418 57774
rect 14366 57698 14418 57710
rect 23102 57762 23154 57774
rect 23102 57698 23154 57710
rect 27806 57762 27858 57774
rect 27806 57698 27858 57710
rect 28590 57762 28642 57774
rect 28590 57698 28642 57710
rect 29710 57762 29762 57774
rect 29710 57698 29762 57710
rect 31278 57762 31330 57774
rect 31278 57698 31330 57710
rect 33630 57762 33682 57774
rect 33630 57698 33682 57710
rect 34526 57762 34578 57774
rect 34526 57698 34578 57710
rect 36318 57762 36370 57774
rect 36318 57698 36370 57710
rect 36990 57762 37042 57774
rect 36990 57698 37042 57710
rect 40350 57762 40402 57774
rect 40350 57698 40402 57710
rect 51214 57762 51266 57774
rect 51214 57698 51266 57710
rect 9998 57650 10050 57662
rect 9998 57586 10050 57598
rect 10446 57650 10498 57662
rect 14254 57650 14306 57662
rect 13794 57598 13806 57650
rect 13858 57598 13870 57650
rect 10446 57586 10498 57598
rect 14254 57586 14306 57598
rect 18958 57650 19010 57662
rect 18958 57586 19010 57598
rect 19854 57650 19906 57662
rect 19854 57586 19906 57598
rect 20078 57650 20130 57662
rect 20078 57586 20130 57598
rect 21982 57650 22034 57662
rect 21982 57586 22034 57598
rect 23438 57650 23490 57662
rect 23438 57586 23490 57598
rect 23662 57650 23714 57662
rect 23662 57586 23714 57598
rect 28702 57650 28754 57662
rect 28702 57586 28754 57598
rect 29150 57650 29202 57662
rect 31166 57650 31218 57662
rect 30594 57598 30606 57650
rect 30658 57598 30670 57650
rect 29150 57586 29202 57598
rect 31166 57586 31218 57598
rect 32062 57650 32114 57662
rect 32062 57586 32114 57598
rect 32398 57650 32450 57662
rect 32398 57586 32450 57598
rect 32734 57650 32786 57662
rect 32734 57586 32786 57598
rect 34750 57650 34802 57662
rect 34750 57586 34802 57598
rect 35086 57650 35138 57662
rect 35086 57586 35138 57598
rect 38222 57650 38274 57662
rect 38222 57586 38274 57598
rect 38446 57650 38498 57662
rect 39230 57650 39282 57662
rect 38658 57598 38670 57650
rect 38722 57598 38734 57650
rect 38446 57586 38498 57598
rect 39230 57586 39282 57598
rect 39454 57650 39506 57662
rect 39454 57586 39506 57598
rect 39790 57650 39842 57662
rect 39790 57586 39842 57598
rect 41806 57650 41858 57662
rect 41806 57586 41858 57598
rect 42814 57650 42866 57662
rect 42814 57586 42866 57598
rect 44382 57650 44434 57662
rect 44382 57586 44434 57598
rect 46286 57650 46338 57662
rect 46286 57586 46338 57598
rect 46510 57650 46562 57662
rect 46510 57586 46562 57598
rect 46958 57650 47010 57662
rect 46958 57586 47010 57598
rect 47518 57650 47570 57662
rect 47518 57586 47570 57598
rect 47742 57650 47794 57662
rect 47742 57586 47794 57598
rect 48078 57650 48130 57662
rect 51886 57650 51938 57662
rect 50194 57598 50206 57650
rect 50258 57598 50270 57650
rect 48078 57586 48130 57598
rect 51886 57586 51938 57598
rect 52110 57650 52162 57662
rect 52110 57586 52162 57598
rect 52334 57650 52386 57662
rect 52334 57586 52386 57598
rect 2158 57538 2210 57550
rect 2158 57474 2210 57486
rect 2830 57538 2882 57550
rect 2830 57474 2882 57486
rect 3726 57538 3778 57550
rect 3726 57474 3778 57486
rect 4622 57538 4674 57550
rect 4622 57474 4674 57486
rect 5070 57538 5122 57550
rect 5070 57474 5122 57486
rect 5518 57538 5570 57550
rect 5518 57474 5570 57486
rect 5854 57538 5906 57550
rect 5854 57474 5906 57486
rect 6414 57538 6466 57550
rect 6414 57474 6466 57486
rect 6862 57538 6914 57550
rect 6862 57474 6914 57486
rect 7198 57538 7250 57550
rect 7198 57474 7250 57486
rect 7646 57538 7698 57550
rect 7646 57474 7698 57486
rect 8094 57538 8146 57550
rect 8094 57474 8146 57486
rect 8542 57538 8594 57550
rect 8542 57474 8594 57486
rect 10894 57538 10946 57550
rect 10894 57474 10946 57486
rect 11230 57538 11282 57550
rect 11230 57474 11282 57486
rect 12014 57538 12066 57550
rect 12014 57474 12066 57486
rect 12350 57538 12402 57550
rect 12350 57474 12402 57486
rect 12798 57538 12850 57550
rect 12798 57474 12850 57486
rect 14926 57538 14978 57550
rect 14926 57474 14978 57486
rect 15374 57538 15426 57550
rect 17614 57538 17666 57550
rect 16258 57486 16270 57538
rect 16322 57486 16334 57538
rect 15374 57474 15426 57486
rect 17614 57474 17666 57486
rect 18174 57538 18226 57550
rect 18174 57474 18226 57486
rect 18734 57538 18786 57550
rect 18734 57474 18786 57486
rect 20974 57538 21026 57550
rect 20974 57474 21026 57486
rect 21422 57538 21474 57550
rect 21422 57474 21474 57486
rect 23214 57538 23266 57550
rect 23214 57474 23266 57486
rect 24110 57538 24162 57550
rect 24110 57474 24162 57486
rect 24558 57538 24610 57550
rect 24558 57474 24610 57486
rect 25566 57538 25618 57550
rect 25566 57474 25618 57486
rect 26014 57538 26066 57550
rect 26014 57474 26066 57486
rect 32510 57538 32562 57550
rect 32510 57474 32562 57486
rect 34974 57538 35026 57550
rect 34974 57474 35026 57486
rect 37438 57538 37490 57550
rect 37438 57474 37490 57486
rect 38334 57538 38386 57550
rect 38334 57474 38386 57486
rect 41582 57538 41634 57550
rect 41582 57474 41634 57486
rect 43374 57538 43426 57550
rect 43374 57474 43426 57486
rect 45054 57538 45106 57550
rect 45054 57474 45106 57486
rect 45502 57538 45554 57550
rect 45502 57474 45554 57486
rect 47854 57538 47906 57550
rect 50542 57538 50594 57550
rect 50306 57486 50318 57538
rect 50370 57486 50382 57538
rect 47854 57474 47906 57486
rect 50542 57474 50594 57486
rect 51998 57538 52050 57550
rect 51998 57474 52050 57486
rect 53118 57538 53170 57550
rect 53118 57474 53170 57486
rect 53566 57538 53618 57550
rect 53566 57474 53618 57486
rect 54014 57538 54066 57550
rect 54014 57474 54066 57486
rect 16606 57426 16658 57438
rect 6738 57374 6750 57426
rect 6802 57423 6814 57426
rect 7858 57423 7870 57426
rect 6802 57377 7870 57423
rect 6802 57374 6814 57377
rect 7858 57374 7870 57377
rect 7922 57374 7934 57426
rect 8082 57374 8094 57426
rect 8146 57423 8158 57426
rect 8530 57423 8542 57426
rect 8146 57377 8542 57423
rect 8146 57374 8158 57377
rect 8530 57374 8542 57377
rect 8594 57374 8606 57426
rect 16606 57362 16658 57374
rect 22206 57426 22258 57438
rect 36542 57426 36594 57438
rect 22530 57374 22542 57426
rect 22594 57374 22606 57426
rect 22206 57362 22258 57374
rect 36542 57362 36594 57374
rect 51326 57426 51378 57438
rect 53106 57374 53118 57426
rect 53170 57423 53182 57426
rect 53890 57423 53902 57426
rect 53170 57377 53902 57423
rect 53170 57374 53182 57377
rect 53890 57374 53902 57377
rect 53954 57374 53966 57426
rect 51326 57362 51378 57374
rect 1344 57258 59024 57292
rect 1344 57206 4478 57258
rect 4530 57206 4582 57258
rect 4634 57206 4686 57258
rect 4738 57206 35198 57258
rect 35250 57206 35302 57258
rect 35354 57206 35406 57258
rect 35458 57206 59024 57258
rect 1344 57172 59024 57206
rect 17726 57090 17778 57102
rect 23550 57090 23602 57102
rect 6962 57038 6974 57090
rect 7026 57087 7038 57090
rect 11106 57087 11118 57090
rect 7026 57041 11118 57087
rect 7026 57038 7038 57041
rect 11106 57038 11118 57041
rect 11170 57038 11182 57090
rect 22754 57038 22766 57090
rect 22818 57038 22830 57090
rect 17726 57026 17778 57038
rect 23550 57026 23602 57038
rect 23998 57090 24050 57102
rect 23998 57026 24050 57038
rect 34638 57090 34690 57102
rect 34638 57026 34690 57038
rect 35646 57090 35698 57102
rect 35646 57026 35698 57038
rect 35870 57090 35922 57102
rect 35870 57026 35922 57038
rect 43486 57090 43538 57102
rect 43486 57026 43538 57038
rect 43822 57090 43874 57102
rect 47058 57038 47070 57090
rect 47122 57038 47134 57090
rect 43822 57026 43874 57038
rect 1934 56978 1986 56990
rect 1934 56914 1986 56926
rect 2382 56978 2434 56990
rect 2382 56914 2434 56926
rect 6974 56978 7026 56990
rect 6974 56914 7026 56926
rect 8206 56978 8258 56990
rect 8206 56914 8258 56926
rect 8766 56978 8818 56990
rect 8766 56914 8818 56926
rect 13582 56978 13634 56990
rect 13582 56914 13634 56926
rect 16718 56978 16770 56990
rect 16718 56914 16770 56926
rect 19070 56978 19122 56990
rect 19070 56914 19122 56926
rect 20190 56978 20242 56990
rect 20190 56914 20242 56926
rect 25790 56978 25842 56990
rect 25790 56914 25842 56926
rect 26126 56978 26178 56990
rect 26126 56914 26178 56926
rect 26574 56978 26626 56990
rect 26574 56914 26626 56926
rect 28702 56978 28754 56990
rect 28702 56914 28754 56926
rect 29598 56978 29650 56990
rect 29598 56914 29650 56926
rect 34750 56978 34802 56990
rect 34750 56914 34802 56926
rect 42590 56978 42642 56990
rect 42590 56914 42642 56926
rect 43262 56978 43314 56990
rect 51998 56978 52050 56990
rect 46274 56926 46286 56978
rect 46338 56926 46350 56978
rect 53778 56926 53790 56978
rect 53842 56926 53854 56978
rect 43262 56914 43314 56926
rect 51998 56914 52050 56926
rect 11118 56866 11170 56878
rect 11118 56802 11170 56814
rect 12350 56866 12402 56878
rect 12350 56802 12402 56814
rect 14142 56866 14194 56878
rect 22206 56866 22258 56878
rect 23774 56866 23826 56878
rect 16034 56814 16046 56866
rect 16098 56814 16110 56866
rect 16482 56814 16494 56866
rect 16546 56814 16558 56866
rect 17490 56814 17502 56866
rect 17554 56814 17566 56866
rect 17826 56814 17838 56866
rect 17890 56814 17902 56866
rect 23314 56814 23326 56866
rect 23378 56814 23390 56866
rect 14142 56802 14194 56814
rect 22206 56802 22258 56814
rect 23774 56802 23826 56814
rect 24558 56866 24610 56878
rect 24558 56802 24610 56814
rect 25006 56866 25058 56878
rect 25006 56802 25058 56814
rect 25118 56866 25170 56878
rect 25118 56802 25170 56814
rect 28814 56866 28866 56878
rect 30494 56866 30546 56878
rect 30034 56814 30046 56866
rect 30098 56814 30110 56866
rect 28814 56802 28866 56814
rect 30494 56802 30546 56814
rect 31054 56866 31106 56878
rect 31054 56802 31106 56814
rect 31726 56866 31778 56878
rect 31726 56802 31778 56814
rect 36094 56866 36146 56878
rect 36094 56802 36146 56814
rect 36318 56866 36370 56878
rect 36318 56802 36370 56814
rect 36542 56866 36594 56878
rect 36542 56802 36594 56814
rect 38670 56866 38722 56878
rect 39342 56866 39394 56878
rect 38770 56814 38782 56866
rect 38834 56814 38846 56866
rect 38670 56802 38722 56814
rect 39342 56802 39394 56814
rect 39454 56866 39506 56878
rect 39454 56802 39506 56814
rect 40014 56866 40066 56878
rect 40014 56802 40066 56814
rect 40686 56866 40738 56878
rect 48190 56866 48242 56878
rect 46386 56814 46398 56866
rect 46450 56814 46462 56866
rect 40686 56802 40738 56814
rect 48190 56802 48242 56814
rect 48302 56866 48354 56878
rect 48302 56802 48354 56814
rect 49982 56866 50034 56878
rect 49982 56802 50034 56814
rect 50094 56866 50146 56878
rect 50094 56802 50146 56814
rect 50654 56866 50706 56878
rect 51202 56814 51214 56866
rect 51266 56814 51278 56866
rect 51650 56814 51662 56866
rect 51714 56814 51726 56866
rect 52210 56814 52222 56866
rect 52274 56814 52286 56866
rect 53330 56814 53342 56866
rect 53394 56814 53406 56866
rect 54114 56814 54126 56866
rect 54178 56814 54190 56866
rect 54674 56814 54686 56866
rect 54738 56814 54750 56866
rect 50654 56802 50706 56814
rect 17278 56754 17330 56766
rect 17278 56690 17330 56702
rect 18958 56754 19010 56766
rect 18958 56690 19010 56702
rect 19182 56754 19234 56766
rect 19182 56690 19234 56702
rect 22094 56754 22146 56766
rect 22094 56690 22146 56702
rect 22318 56754 22370 56766
rect 22318 56690 22370 56702
rect 24110 56754 24162 56766
rect 24110 56690 24162 56702
rect 28590 56754 28642 56766
rect 28590 56690 28642 56702
rect 31502 56754 31554 56766
rect 31502 56690 31554 56702
rect 32174 56754 32226 56766
rect 32174 56690 32226 56702
rect 36430 56754 36482 56766
rect 36430 56690 36482 56702
rect 38558 56754 38610 56766
rect 38558 56690 38610 56702
rect 48414 56754 48466 56766
rect 52322 56702 52334 56754
rect 52386 56702 52398 56754
rect 48414 56690 48466 56702
rect 2830 56642 2882 56654
rect 2830 56578 2882 56590
rect 3502 56642 3554 56654
rect 3502 56578 3554 56590
rect 3950 56642 4002 56654
rect 3950 56578 4002 56590
rect 4286 56642 4338 56654
rect 4286 56578 4338 56590
rect 4846 56642 4898 56654
rect 4846 56578 4898 56590
rect 6078 56642 6130 56654
rect 6078 56578 6130 56590
rect 6414 56642 6466 56654
rect 6414 56578 6466 56590
rect 7422 56642 7474 56654
rect 7422 56578 7474 56590
rect 7870 56642 7922 56654
rect 7870 56578 7922 56590
rect 9214 56642 9266 56654
rect 9214 56578 9266 56590
rect 9774 56642 9826 56654
rect 9774 56578 9826 56590
rect 10222 56642 10274 56654
rect 10222 56578 10274 56590
rect 10670 56642 10722 56654
rect 10670 56578 10722 56590
rect 11566 56642 11618 56654
rect 11566 56578 11618 56590
rect 11902 56642 11954 56654
rect 11902 56578 11954 56590
rect 12686 56642 12738 56654
rect 12686 56578 12738 56590
rect 12910 56642 12962 56654
rect 12910 56578 12962 56590
rect 13022 56642 13074 56654
rect 13022 56578 13074 56590
rect 14590 56642 14642 56654
rect 14590 56578 14642 56590
rect 15038 56642 15090 56654
rect 15038 56578 15090 56590
rect 18062 56642 18114 56654
rect 18062 56578 18114 56590
rect 19854 56642 19906 56654
rect 19854 56578 19906 56590
rect 20750 56642 20802 56654
rect 20750 56578 20802 56590
rect 25230 56642 25282 56654
rect 25230 56578 25282 56590
rect 27022 56642 27074 56654
rect 27022 56578 27074 56590
rect 31390 56642 31442 56654
rect 31390 56578 31442 56590
rect 32622 56642 32674 56654
rect 32622 56578 32674 56590
rect 37662 56642 37714 56654
rect 37662 56578 37714 56590
rect 39006 56642 39058 56654
rect 39006 56578 39058 56590
rect 40126 56642 40178 56654
rect 40126 56578 40178 56590
rect 40238 56642 40290 56654
rect 40238 56578 40290 56590
rect 41022 56642 41074 56654
rect 50206 56642 50258 56654
rect 47730 56590 47742 56642
rect 47794 56590 47806 56642
rect 41022 56578 41074 56590
rect 50206 56578 50258 56590
rect 55246 56642 55298 56654
rect 55246 56578 55298 56590
rect 1344 56474 59024 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 59024 56474
rect 1344 56388 59024 56422
rect 2718 56306 2770 56318
rect 2718 56242 2770 56254
rect 5406 56306 5458 56318
rect 5406 56242 5458 56254
rect 5854 56306 5906 56318
rect 5854 56242 5906 56254
rect 6862 56306 6914 56318
rect 6862 56242 6914 56254
rect 7646 56306 7698 56318
rect 7646 56242 7698 56254
rect 8542 56306 8594 56318
rect 8542 56242 8594 56254
rect 11118 56306 11170 56318
rect 11118 56242 11170 56254
rect 14366 56306 14418 56318
rect 14366 56242 14418 56254
rect 15262 56306 15314 56318
rect 15262 56242 15314 56254
rect 16494 56306 16546 56318
rect 16494 56242 16546 56254
rect 16942 56306 16994 56318
rect 16942 56242 16994 56254
rect 18622 56306 18674 56318
rect 18622 56242 18674 56254
rect 20974 56306 21026 56318
rect 20974 56242 21026 56254
rect 22542 56306 22594 56318
rect 22542 56242 22594 56254
rect 23662 56306 23714 56318
rect 23662 56242 23714 56254
rect 26462 56306 26514 56318
rect 26462 56242 26514 56254
rect 27806 56306 27858 56318
rect 27806 56242 27858 56254
rect 30158 56306 30210 56318
rect 30158 56242 30210 56254
rect 30718 56306 30770 56318
rect 30718 56242 30770 56254
rect 35534 56306 35586 56318
rect 35534 56242 35586 56254
rect 38222 56306 38274 56318
rect 38222 56242 38274 56254
rect 40014 56306 40066 56318
rect 40014 56242 40066 56254
rect 42814 56306 42866 56318
rect 42814 56242 42866 56254
rect 43934 56306 43986 56318
rect 43934 56242 43986 56254
rect 44158 56306 44210 56318
rect 44158 56242 44210 56254
rect 51102 56306 51154 56318
rect 51102 56242 51154 56254
rect 54014 56306 54066 56318
rect 54014 56242 54066 56254
rect 9998 56194 10050 56206
rect 9998 56130 10050 56142
rect 12798 56194 12850 56206
rect 12798 56130 12850 56142
rect 13470 56194 13522 56206
rect 13470 56130 13522 56142
rect 13694 56194 13746 56206
rect 13694 56130 13746 56142
rect 19294 56194 19346 56206
rect 19294 56130 19346 56142
rect 46510 56194 46562 56206
rect 46510 56130 46562 56142
rect 51214 56194 51266 56206
rect 51214 56130 51266 56142
rect 52334 56194 52386 56206
rect 52334 56130 52386 56142
rect 1934 56082 1986 56094
rect 1934 56018 1986 56030
rect 8094 56082 8146 56094
rect 8094 56018 8146 56030
rect 11006 56082 11058 56094
rect 11006 56018 11058 56030
rect 11342 56082 11394 56094
rect 14254 56082 14306 56094
rect 12114 56030 12126 56082
rect 12178 56030 12190 56082
rect 11342 56018 11394 56030
rect 14254 56018 14306 56030
rect 21422 56082 21474 56094
rect 21422 56018 21474 56030
rect 21982 56082 22034 56094
rect 22430 56082 22482 56094
rect 22306 56030 22318 56082
rect 22370 56030 22382 56082
rect 21982 56018 22034 56030
rect 22430 56018 22482 56030
rect 22654 56082 22706 56094
rect 22654 56018 22706 56030
rect 23886 56082 23938 56094
rect 23886 56018 23938 56030
rect 24334 56082 24386 56094
rect 24334 56018 24386 56030
rect 26238 56082 26290 56094
rect 26238 56018 26290 56030
rect 26574 56082 26626 56094
rect 26574 56018 26626 56030
rect 26798 56082 26850 56094
rect 26798 56018 26850 56030
rect 39118 56082 39170 56094
rect 39118 56018 39170 56030
rect 39342 56082 39394 56094
rect 39342 56018 39394 56030
rect 44606 56082 44658 56094
rect 44606 56018 44658 56030
rect 46734 56082 46786 56094
rect 51998 56082 52050 56094
rect 50194 56030 50206 56082
rect 50258 56030 50270 56082
rect 51762 56030 51774 56082
rect 51826 56030 51838 56082
rect 46734 56018 46786 56030
rect 51998 56018 52050 56030
rect 52222 56082 52274 56094
rect 52222 56018 52274 56030
rect 2382 55970 2434 55982
rect 2382 55906 2434 55918
rect 3166 55970 3218 55982
rect 3166 55906 3218 55918
rect 3614 55970 3666 55982
rect 3614 55906 3666 55918
rect 4062 55970 4114 55982
rect 4062 55906 4114 55918
rect 4622 55970 4674 55982
rect 4622 55906 4674 55918
rect 5070 55970 5122 55982
rect 5070 55906 5122 55918
rect 6302 55970 6354 55982
rect 6302 55906 6354 55918
rect 7310 55970 7362 55982
rect 7310 55906 7362 55918
rect 8990 55970 9042 55982
rect 8990 55906 9042 55918
rect 10446 55970 10498 55982
rect 14030 55970 14082 55982
rect 11890 55918 11902 55970
rect 11954 55918 11966 55970
rect 10446 55906 10498 55918
rect 14030 55906 14082 55918
rect 14926 55970 14978 55982
rect 14926 55906 14978 55918
rect 16046 55970 16098 55982
rect 16046 55906 16098 55918
rect 17614 55970 17666 55982
rect 17614 55906 17666 55918
rect 18174 55970 18226 55982
rect 20190 55970 20242 55982
rect 19170 55918 19182 55970
rect 19234 55918 19246 55970
rect 18174 55906 18226 55918
rect 20190 55906 20242 55918
rect 23774 55970 23826 55982
rect 23774 55906 23826 55918
rect 24670 55970 24722 55982
rect 24670 55906 24722 55918
rect 25566 55970 25618 55982
rect 25566 55906 25618 55918
rect 27358 55970 27410 55982
rect 27358 55906 27410 55918
rect 28254 55970 28306 55982
rect 28254 55906 28306 55918
rect 31278 55970 31330 55982
rect 31278 55906 31330 55918
rect 31838 55970 31890 55982
rect 31838 55906 31890 55918
rect 35086 55970 35138 55982
rect 35086 55906 35138 55918
rect 38558 55970 38610 55982
rect 38558 55906 38610 55918
rect 40350 55970 40402 55982
rect 40350 55906 40402 55918
rect 43374 55970 43426 55982
rect 44382 55970 44434 55982
rect 44034 55918 44046 55970
rect 44098 55918 44110 55970
rect 43374 55906 43426 55918
rect 44382 55906 44434 55918
rect 44830 55970 44882 55982
rect 44830 55906 44882 55918
rect 48302 55970 48354 55982
rect 48302 55906 48354 55918
rect 49534 55970 49586 55982
rect 52894 55970 52946 55982
rect 50306 55918 50318 55970
rect 50370 55918 50382 55970
rect 49534 55906 49586 55918
rect 52894 55906 52946 55918
rect 53902 55970 53954 55982
rect 53902 55906 53954 55918
rect 54462 55970 54514 55982
rect 54462 55906 54514 55918
rect 19518 55858 19570 55870
rect 5954 55806 5966 55858
rect 6018 55855 6030 55858
rect 7858 55855 7870 55858
rect 6018 55809 7870 55855
rect 6018 55806 6030 55809
rect 7858 55806 7870 55809
rect 7922 55806 7934 55858
rect 19518 55794 19570 55806
rect 20078 55858 20130 55870
rect 20078 55794 20130 55806
rect 31390 55858 31442 55870
rect 31390 55794 31442 55806
rect 39566 55858 39618 55870
rect 39566 55794 39618 55806
rect 47070 55858 47122 55870
rect 47070 55794 47122 55806
rect 1344 55690 59024 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 59024 55690
rect 1344 55604 59024 55638
rect 14142 55522 14194 55534
rect 22990 55522 23042 55534
rect 38782 55522 38834 55534
rect 6738 55470 6750 55522
rect 6802 55519 6814 55522
rect 6962 55519 6974 55522
rect 6802 55473 6974 55519
rect 6802 55470 6814 55473
rect 6962 55470 6974 55473
rect 7026 55470 7038 55522
rect 7634 55470 7646 55522
rect 7698 55519 7710 55522
rect 8194 55519 8206 55522
rect 7698 55473 8206 55519
rect 7698 55470 7710 55473
rect 8194 55470 8206 55473
rect 8258 55519 8270 55522
rect 8866 55519 8878 55522
rect 8258 55473 8878 55519
rect 8258 55470 8270 55473
rect 8866 55470 8878 55473
rect 8930 55470 8942 55522
rect 10658 55470 10670 55522
rect 10722 55519 10734 55522
rect 11666 55519 11678 55522
rect 10722 55473 11678 55519
rect 10722 55470 10734 55473
rect 11666 55470 11678 55473
rect 11730 55470 11742 55522
rect 14466 55470 14478 55522
rect 14530 55519 14542 55522
rect 14914 55519 14926 55522
rect 14530 55473 14926 55519
rect 14530 55470 14542 55473
rect 14914 55470 14926 55473
rect 14978 55470 14990 55522
rect 37538 55470 37550 55522
rect 37602 55470 37614 55522
rect 43250 55470 43262 55522
rect 43314 55470 43326 55522
rect 14142 55458 14194 55470
rect 22990 55458 23042 55470
rect 38782 55458 38834 55470
rect 3614 55410 3666 55422
rect 3614 55346 3666 55358
rect 5854 55410 5906 55422
rect 5854 55346 5906 55358
rect 6750 55410 6802 55422
rect 6750 55346 6802 55358
rect 7646 55410 7698 55422
rect 7646 55346 7698 55358
rect 8542 55410 8594 55422
rect 12910 55410 12962 55422
rect 15150 55410 15202 55422
rect 18958 55410 19010 55422
rect 12114 55358 12126 55410
rect 12178 55358 12190 55410
rect 13794 55358 13806 55410
rect 13858 55358 13870 55410
rect 16594 55358 16606 55410
rect 16658 55358 16670 55410
rect 8542 55346 8594 55358
rect 12910 55346 12962 55358
rect 15150 55346 15202 55358
rect 18958 55346 19010 55358
rect 20638 55410 20690 55422
rect 28030 55410 28082 55422
rect 23314 55358 23326 55410
rect 23378 55358 23390 55410
rect 25554 55358 25566 55410
rect 25618 55358 25630 55410
rect 20638 55346 20690 55358
rect 28030 55346 28082 55358
rect 32286 55410 32338 55422
rect 41358 55410 41410 55422
rect 46510 55410 46562 55422
rect 35970 55358 35982 55410
rect 36034 55358 36046 55410
rect 42578 55358 42590 55410
rect 42642 55358 42654 55410
rect 32286 55346 32338 55358
rect 41358 55346 41410 55358
rect 46510 55346 46562 55358
rect 47854 55410 47906 55422
rect 53666 55358 53678 55410
rect 53730 55358 53742 55410
rect 47854 55346 47906 55358
rect 19742 55298 19794 55310
rect 24670 55298 24722 55310
rect 26462 55298 26514 55310
rect 12450 55246 12462 55298
rect 12514 55246 12526 55298
rect 18722 55246 18734 55298
rect 18786 55246 18798 55298
rect 19954 55246 19966 55298
rect 20018 55246 20030 55298
rect 26002 55246 26014 55298
rect 26066 55246 26078 55298
rect 19742 55234 19794 55246
rect 24670 55234 24722 55246
rect 26462 55234 26514 55246
rect 27134 55298 27186 55310
rect 32174 55298 32226 55310
rect 27570 55246 27582 55298
rect 27634 55246 27646 55298
rect 27134 55234 27186 55246
rect 32174 55234 32226 55246
rect 33406 55298 33458 55310
rect 34302 55298 34354 55310
rect 37886 55298 37938 55310
rect 33730 55246 33742 55298
rect 33794 55246 33806 55298
rect 35634 55246 35646 55298
rect 35698 55246 35710 55298
rect 33406 55234 33458 55246
rect 34302 55234 34354 55246
rect 37886 55234 37938 55246
rect 38110 55298 38162 55310
rect 39678 55298 39730 55310
rect 39442 55246 39454 55298
rect 39506 55246 39518 55298
rect 38110 55234 38162 55246
rect 39678 55234 39730 55246
rect 40462 55298 40514 55310
rect 46958 55298 47010 55310
rect 47518 55298 47570 55310
rect 40674 55246 40686 55298
rect 40738 55246 40750 55298
rect 42466 55246 42478 55298
rect 42530 55246 42542 55298
rect 47282 55246 47294 55298
rect 47346 55246 47358 55298
rect 40462 55234 40514 55246
rect 46958 55234 47010 55246
rect 47518 55234 47570 55246
rect 47742 55298 47794 55310
rect 47742 55234 47794 55246
rect 1822 55186 1874 55198
rect 1822 55122 1874 55134
rect 9998 55186 10050 55198
rect 9998 55122 10050 55134
rect 16718 55186 16770 55198
rect 16718 55122 16770 55134
rect 16942 55186 16994 55198
rect 16942 55122 16994 55134
rect 19070 55186 19122 55198
rect 19070 55122 19122 55134
rect 28478 55186 28530 55198
rect 28478 55122 28530 55134
rect 29934 55186 29986 55198
rect 29934 55122 29986 55134
rect 32510 55186 32562 55198
rect 32510 55122 32562 55134
rect 32734 55186 32786 55198
rect 32734 55122 32786 55134
rect 36318 55186 36370 55198
rect 36318 55122 36370 55134
rect 38670 55186 38722 55198
rect 38670 55122 38722 55134
rect 39790 55186 39842 55198
rect 39790 55122 39842 55134
rect 47966 55186 48018 55198
rect 47966 55122 48018 55134
rect 48414 55186 48466 55198
rect 48414 55122 48466 55134
rect 53790 55186 53842 55198
rect 53790 55122 53842 55134
rect 54014 55186 54066 55198
rect 54014 55122 54066 55134
rect 2158 55074 2210 55086
rect 2158 55010 2210 55022
rect 2606 55074 2658 55086
rect 2606 55010 2658 55022
rect 3054 55074 3106 55086
rect 3054 55010 3106 55022
rect 3950 55074 4002 55086
rect 3950 55010 4002 55022
rect 4398 55074 4450 55086
rect 4398 55010 4450 55022
rect 4846 55074 4898 55086
rect 4846 55010 4898 55022
rect 6414 55074 6466 55086
rect 6414 55010 6466 55022
rect 7198 55074 7250 55086
rect 7198 55010 7250 55022
rect 8094 55074 8146 55086
rect 8094 55010 8146 55022
rect 8990 55074 9042 55086
rect 8990 55010 9042 55022
rect 9550 55074 9602 55086
rect 9550 55010 9602 55022
rect 10446 55074 10498 55086
rect 10446 55010 10498 55022
rect 10894 55074 10946 55086
rect 10894 55010 10946 55022
rect 11342 55074 11394 55086
rect 11342 55010 11394 55022
rect 13918 55074 13970 55086
rect 13918 55010 13970 55022
rect 14590 55074 14642 55086
rect 14590 55010 14642 55022
rect 15710 55074 15762 55086
rect 15710 55010 15762 55022
rect 16158 55074 16210 55086
rect 16158 55010 16210 55022
rect 17390 55074 17442 55086
rect 17390 55010 17442 55022
rect 17838 55074 17890 55086
rect 17838 55010 17890 55022
rect 21758 55074 21810 55086
rect 21758 55010 21810 55022
rect 22206 55074 22258 55086
rect 22206 55010 22258 55022
rect 23214 55074 23266 55086
rect 23214 55010 23266 55022
rect 23774 55074 23826 55086
rect 23774 55010 23826 55022
rect 24222 55074 24274 55086
rect 24222 55010 24274 55022
rect 29822 55074 29874 55086
rect 29822 55010 29874 55022
rect 38782 55074 38834 55086
rect 38782 55010 38834 55022
rect 49086 55074 49138 55086
rect 49086 55010 49138 55022
rect 54462 55074 54514 55086
rect 54462 55010 54514 55022
rect 1344 54906 59024 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 59024 54906
rect 1344 54820 59024 54854
rect 2270 54738 2322 54750
rect 2270 54674 2322 54686
rect 2718 54738 2770 54750
rect 2718 54674 2770 54686
rect 7646 54738 7698 54750
rect 7646 54674 7698 54686
rect 8542 54738 8594 54750
rect 8542 54674 8594 54686
rect 8990 54738 9042 54750
rect 8990 54674 9042 54686
rect 10558 54738 10610 54750
rect 10558 54674 10610 54686
rect 11454 54738 11506 54750
rect 11454 54674 11506 54686
rect 12014 54738 12066 54750
rect 12014 54674 12066 54686
rect 13022 54738 13074 54750
rect 21870 54738 21922 54750
rect 16818 54686 16830 54738
rect 16882 54686 16894 54738
rect 13022 54674 13074 54686
rect 21870 54674 21922 54686
rect 22766 54738 22818 54750
rect 22766 54674 22818 54686
rect 23998 54738 24050 54750
rect 23998 54674 24050 54686
rect 24446 54738 24498 54750
rect 35422 54738 35474 54750
rect 26674 54686 26686 54738
rect 26738 54686 26750 54738
rect 24446 54674 24498 54686
rect 35422 54674 35474 54686
rect 35534 54738 35586 54750
rect 35534 54674 35586 54686
rect 41806 54738 41858 54750
rect 41806 54674 41858 54686
rect 46398 54738 46450 54750
rect 46398 54674 46450 54686
rect 47406 54738 47458 54750
rect 47406 54674 47458 54686
rect 48302 54738 48354 54750
rect 48302 54674 48354 54686
rect 48414 54738 48466 54750
rect 48414 54674 48466 54686
rect 51438 54738 51490 54750
rect 51438 54674 51490 54686
rect 52222 54738 52274 54750
rect 52222 54674 52274 54686
rect 53454 54738 53506 54750
rect 53454 54674 53506 54686
rect 1822 54626 1874 54638
rect 1822 54562 1874 54574
rect 13246 54626 13298 54638
rect 13246 54562 13298 54574
rect 14030 54626 14082 54638
rect 14030 54562 14082 54574
rect 14142 54626 14194 54638
rect 19070 54626 19122 54638
rect 15026 54574 15038 54626
rect 15090 54574 15102 54626
rect 16594 54574 16606 54626
rect 16658 54574 16670 54626
rect 14142 54562 14194 54574
rect 19070 54562 19122 54574
rect 27134 54626 27186 54638
rect 27134 54562 27186 54574
rect 32846 54626 32898 54638
rect 32846 54562 32898 54574
rect 39454 54626 39506 54638
rect 39454 54562 39506 54574
rect 41918 54626 41970 54638
rect 41918 54562 41970 54574
rect 42926 54626 42978 54638
rect 42926 54562 42978 54574
rect 46174 54626 46226 54638
rect 46174 54562 46226 54574
rect 47294 54626 47346 54638
rect 47294 54562 47346 54574
rect 48526 54626 48578 54638
rect 48526 54562 48578 54574
rect 50542 54626 50594 54638
rect 50542 54562 50594 54574
rect 52446 54626 52498 54638
rect 52446 54562 52498 54574
rect 54350 54626 54402 54638
rect 54350 54562 54402 54574
rect 4398 54514 4450 54526
rect 4398 54450 4450 54462
rect 4958 54514 5010 54526
rect 19966 54514 20018 54526
rect 13794 54462 13806 54514
rect 13858 54462 13870 54514
rect 15586 54462 15598 54514
rect 15650 54462 15662 54514
rect 19506 54462 19518 54514
rect 19570 54462 19582 54514
rect 4958 54450 5010 54462
rect 19966 54450 20018 54462
rect 27246 54514 27298 54526
rect 28142 54514 28194 54526
rect 29038 54514 29090 54526
rect 46062 54514 46114 54526
rect 51214 54514 51266 54526
rect 27458 54462 27470 54514
rect 27522 54462 27534 54514
rect 28578 54462 28590 54514
rect 28642 54462 28654 54514
rect 30146 54462 30158 54514
rect 30210 54462 30222 54514
rect 32386 54462 32398 54514
rect 32450 54462 32462 54514
rect 35746 54462 35758 54514
rect 35810 54511 35822 54514
rect 35970 54511 35982 54514
rect 35810 54465 35982 54511
rect 35810 54462 35822 54465
rect 35970 54462 35982 54465
rect 36034 54462 36046 54514
rect 36530 54462 36542 54514
rect 36594 54462 36606 54514
rect 41570 54462 41582 54514
rect 41634 54462 41646 54514
rect 48066 54462 48078 54514
rect 48130 54462 48142 54514
rect 48738 54462 48750 54514
rect 48802 54462 48814 54514
rect 49858 54462 49870 54514
rect 49922 54462 49934 54514
rect 27246 54450 27298 54462
rect 28142 54450 28194 54462
rect 29038 54450 29090 54462
rect 46062 54450 46114 54462
rect 51214 54450 51266 54462
rect 51438 54514 51490 54526
rect 51438 54450 51490 54462
rect 51774 54514 51826 54526
rect 51774 54450 51826 54462
rect 52558 54514 52610 54526
rect 52558 54450 52610 54462
rect 53006 54514 53058 54526
rect 53006 54450 53058 54462
rect 53678 54514 53730 54526
rect 53678 54450 53730 54462
rect 54238 54514 54290 54526
rect 54238 54450 54290 54462
rect 3166 54402 3218 54414
rect 3166 54338 3218 54350
rect 3502 54402 3554 54414
rect 3502 54338 3554 54350
rect 3950 54402 4002 54414
rect 3950 54338 4002 54350
rect 5294 54402 5346 54414
rect 5294 54338 5346 54350
rect 5742 54402 5794 54414
rect 5742 54338 5794 54350
rect 6414 54402 6466 54414
rect 6414 54338 6466 54350
rect 6750 54402 6802 54414
rect 6750 54338 6802 54350
rect 7310 54402 7362 54414
rect 7310 54338 7362 54350
rect 8206 54402 8258 54414
rect 8206 54338 8258 54350
rect 9662 54402 9714 54414
rect 9662 54338 9714 54350
rect 10222 54402 10274 54414
rect 10222 54338 10274 54350
rect 11118 54402 11170 54414
rect 11118 54338 11170 54350
rect 12350 54402 12402 54414
rect 17614 54402 17666 54414
rect 12898 54350 12910 54402
rect 12962 54350 12974 54402
rect 12350 54338 12402 54350
rect 17614 54338 17666 54350
rect 18062 54402 18114 54414
rect 18062 54338 18114 54350
rect 18622 54402 18674 54414
rect 18622 54338 18674 54350
rect 20638 54402 20690 54414
rect 20638 54338 20690 54350
rect 21086 54402 21138 54414
rect 21086 54338 21138 54350
rect 22318 54402 22370 54414
rect 22318 54338 22370 54350
rect 23326 54402 23378 54414
rect 23326 54338 23378 54350
rect 25006 54402 25058 54414
rect 25006 54338 25058 54350
rect 25678 54402 25730 54414
rect 25678 54338 25730 54350
rect 26126 54402 26178 54414
rect 30830 54402 30882 54414
rect 33742 54402 33794 54414
rect 29922 54350 29934 54402
rect 29986 54350 29998 54402
rect 32498 54350 32510 54402
rect 32562 54350 32574 54402
rect 26126 54338 26178 54350
rect 30830 54338 30882 54350
rect 33742 54338 33794 54350
rect 35646 54402 35698 54414
rect 43038 54402 43090 54414
rect 53566 54402 53618 54414
rect 36418 54350 36430 54402
rect 36482 54350 36494 54402
rect 39330 54350 39342 54402
rect 39394 54350 39406 54402
rect 50082 54350 50094 54402
rect 50146 54350 50158 54402
rect 35646 54338 35698 54350
rect 43038 54338 43090 54350
rect 53566 54338 53618 54350
rect 33630 54290 33682 54302
rect 2146 54238 2158 54290
rect 2210 54287 2222 54290
rect 2482 54287 2494 54290
rect 2210 54241 2494 54287
rect 2210 54238 2222 54241
rect 2482 54238 2494 54241
rect 2546 54238 2558 54290
rect 10882 54238 10894 54290
rect 10946 54287 10958 54290
rect 12338 54287 12350 54290
rect 10946 54241 12350 54287
rect 10946 54238 10958 54241
rect 12338 54238 12350 54241
rect 12402 54238 12414 54290
rect 33630 54226 33682 54238
rect 36206 54290 36258 54302
rect 36206 54226 36258 54238
rect 39678 54290 39730 54302
rect 39678 54226 39730 54238
rect 43150 54290 43202 54302
rect 43150 54226 43202 54238
rect 47518 54290 47570 54302
rect 47518 54226 47570 54238
rect 1344 54122 59024 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 59024 54122
rect 1344 54036 59024 54070
rect 14030 53954 14082 53966
rect 5842 53902 5854 53954
rect 5906 53951 5918 53954
rect 6290 53951 6302 53954
rect 5906 53905 6302 53951
rect 5906 53902 5918 53905
rect 6290 53902 6302 53905
rect 6354 53902 6366 53954
rect 14030 53890 14082 53902
rect 15822 53954 15874 53966
rect 15822 53890 15874 53902
rect 15934 53954 15986 53966
rect 15934 53890 15986 53902
rect 16382 53954 16434 53966
rect 16382 53890 16434 53902
rect 16606 53954 16658 53966
rect 16606 53890 16658 53902
rect 19070 53954 19122 53966
rect 19070 53890 19122 53902
rect 28702 53954 28754 53966
rect 28702 53890 28754 53902
rect 32510 53954 32562 53966
rect 40338 53902 40350 53954
rect 40402 53902 40414 53954
rect 32510 53890 32562 53902
rect 3278 53842 3330 53854
rect 3278 53778 3330 53790
rect 3726 53842 3778 53854
rect 3726 53778 3778 53790
rect 7086 53842 7138 53854
rect 7086 53778 7138 53790
rect 8766 53842 8818 53854
rect 8766 53778 8818 53790
rect 9662 53842 9714 53854
rect 9662 53778 9714 53790
rect 11902 53842 11954 53854
rect 18510 53842 18562 53854
rect 12226 53790 12238 53842
rect 12290 53790 12302 53842
rect 13682 53790 13694 53842
rect 13746 53790 13758 53842
rect 11902 53778 11954 53790
rect 18510 53778 18562 53790
rect 20414 53842 20466 53854
rect 20414 53778 20466 53790
rect 20526 53842 20578 53854
rect 20526 53778 20578 53790
rect 29710 53842 29762 53854
rect 35982 53842 36034 53854
rect 42702 53842 42754 53854
rect 32722 53790 32734 53842
rect 32786 53790 32798 53842
rect 39666 53790 39678 53842
rect 39730 53790 39742 53842
rect 29710 53778 29762 53790
rect 35982 53778 36034 53790
rect 42702 53778 42754 53790
rect 44718 53842 44770 53854
rect 52222 53842 52274 53854
rect 45938 53790 45950 53842
rect 46002 53790 46014 53842
rect 48178 53790 48190 53842
rect 48242 53790 48254 53842
rect 44718 53778 44770 53790
rect 52222 53778 52274 53790
rect 2382 53730 2434 53742
rect 2382 53666 2434 53678
rect 4174 53730 4226 53742
rect 4174 53666 4226 53678
rect 4958 53730 5010 53742
rect 4958 53666 5010 53678
rect 6526 53730 6578 53742
rect 6526 53666 6578 53678
rect 7534 53730 7586 53742
rect 7534 53666 7586 53678
rect 9214 53730 9266 53742
rect 9214 53666 9266 53678
rect 10110 53730 10162 53742
rect 14590 53730 14642 53742
rect 12562 53678 12574 53730
rect 12626 53678 12638 53730
rect 10110 53666 10162 53678
rect 14590 53666 14642 53678
rect 14926 53730 14978 53742
rect 14926 53666 14978 53678
rect 15934 53730 15986 53742
rect 19630 53730 19682 53742
rect 19394 53678 19406 53730
rect 19458 53678 19470 53730
rect 15934 53666 15986 53678
rect 19630 53666 19682 53678
rect 19742 53730 19794 53742
rect 23998 53730 24050 53742
rect 22418 53678 22430 53730
rect 22482 53678 22494 53730
rect 23650 53678 23662 53730
rect 23714 53678 23726 53730
rect 19742 53666 19794 53678
rect 23998 53666 24050 53678
rect 24222 53730 24274 53742
rect 24222 53666 24274 53678
rect 26238 53730 26290 53742
rect 26238 53666 26290 53678
rect 27246 53730 27298 53742
rect 27246 53666 27298 53678
rect 27582 53730 27634 53742
rect 27582 53666 27634 53678
rect 29598 53730 29650 53742
rect 29598 53666 29650 53678
rect 29822 53730 29874 53742
rect 35422 53730 35474 53742
rect 30146 53678 30158 53730
rect 30210 53678 30222 53730
rect 29822 53666 29874 53678
rect 35422 53666 35474 53678
rect 35758 53730 35810 53742
rect 35758 53666 35810 53678
rect 36430 53730 36482 53742
rect 41694 53730 41746 53742
rect 46846 53730 46898 53742
rect 39554 53678 39566 53730
rect 39618 53678 39630 53730
rect 44034 53678 44046 53730
rect 44098 53678 44110 53730
rect 46162 53678 46174 53730
rect 46226 53678 46238 53730
rect 36430 53666 36482 53678
rect 41694 53666 41746 53678
rect 46846 53666 46898 53678
rect 48526 53730 48578 53742
rect 48526 53666 48578 53678
rect 49422 53730 49474 53742
rect 49422 53666 49474 53678
rect 51326 53730 51378 53742
rect 53454 53730 53506 53742
rect 51762 53678 51774 53730
rect 51826 53678 51838 53730
rect 51326 53666 51378 53678
rect 53454 53666 53506 53678
rect 53566 53730 53618 53742
rect 53890 53678 53902 53730
rect 53954 53678 53966 53730
rect 53566 53666 53618 53678
rect 2046 53618 2098 53630
rect 2046 53554 2098 53566
rect 14702 53618 14754 53630
rect 14702 53554 14754 53566
rect 22990 53618 23042 53630
rect 22990 53554 23042 53566
rect 27358 53618 27410 53630
rect 27358 53554 27410 53566
rect 28814 53618 28866 53630
rect 28814 53554 28866 53566
rect 32734 53618 32786 53630
rect 32734 53554 32786 53566
rect 33406 53618 33458 53630
rect 33406 53554 33458 53566
rect 33518 53618 33570 53630
rect 33518 53554 33570 53566
rect 35086 53618 35138 53630
rect 35086 53554 35138 53566
rect 36206 53618 36258 53630
rect 48190 53618 48242 53630
rect 43026 53566 43038 53618
rect 43090 53566 43102 53618
rect 36206 53554 36258 53566
rect 48190 53554 48242 53566
rect 49086 53618 49138 53630
rect 49086 53554 49138 53566
rect 2830 53506 2882 53518
rect 2830 53442 2882 53454
rect 5630 53506 5682 53518
rect 5630 53442 5682 53454
rect 6078 53506 6130 53518
rect 6078 53442 6130 53454
rect 7982 53506 8034 53518
rect 7982 53442 8034 53454
rect 8318 53506 8370 53518
rect 8318 53442 8370 53454
rect 10894 53506 10946 53518
rect 10894 53442 10946 53454
rect 11342 53506 11394 53518
rect 11342 53442 11394 53454
rect 13806 53506 13858 53518
rect 13806 53442 13858 53454
rect 15374 53506 15426 53518
rect 15374 53442 15426 53454
rect 17166 53506 17218 53518
rect 17166 53442 17218 53454
rect 17614 53506 17666 53518
rect 17614 53442 17666 53454
rect 18062 53506 18114 53518
rect 18062 53442 18114 53454
rect 19518 53506 19570 53518
rect 19518 53442 19570 53454
rect 20638 53506 20690 53518
rect 20638 53442 20690 53454
rect 21982 53506 22034 53518
rect 21982 53442 22034 53454
rect 22654 53506 22706 53518
rect 22654 53442 22706 53454
rect 22766 53506 22818 53518
rect 22766 53442 22818 53454
rect 22878 53506 22930 53518
rect 22878 53442 22930 53454
rect 23886 53506 23938 53518
rect 23886 53442 23938 53454
rect 24110 53506 24162 53518
rect 24110 53442 24162 53454
rect 24894 53506 24946 53518
rect 24894 53442 24946 53454
rect 25342 53506 25394 53518
rect 25342 53442 25394 53454
rect 25678 53506 25730 53518
rect 25678 53442 25730 53454
rect 26798 53506 26850 53518
rect 26798 53442 26850 53454
rect 28030 53506 28082 53518
rect 28030 53442 28082 53454
rect 35198 53506 35250 53518
rect 35198 53442 35250 53454
rect 41806 53506 41858 53518
rect 41806 53442 41858 53454
rect 42030 53506 42082 53518
rect 42030 53442 42082 53454
rect 47294 53506 47346 53518
rect 47294 53442 47346 53454
rect 47966 53506 48018 53518
rect 47966 53442 48018 53454
rect 49198 53506 49250 53518
rect 49198 53442 49250 53454
rect 1344 53338 59024 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 59024 53338
rect 1344 53252 59024 53286
rect 3054 53170 3106 53182
rect 3054 53106 3106 53118
rect 4510 53170 4562 53182
rect 4510 53106 4562 53118
rect 5070 53170 5122 53182
rect 5070 53106 5122 53118
rect 5854 53170 5906 53182
rect 5854 53106 5906 53118
rect 6302 53170 6354 53182
rect 6302 53106 6354 53118
rect 6750 53170 6802 53182
rect 6750 53106 6802 53118
rect 7198 53170 7250 53182
rect 7198 53106 7250 53118
rect 8990 53170 9042 53182
rect 8990 53106 9042 53118
rect 9886 53170 9938 53182
rect 9886 53106 9938 53118
rect 10334 53170 10386 53182
rect 10334 53106 10386 53118
rect 11790 53170 11842 53182
rect 11790 53106 11842 53118
rect 12686 53170 12738 53182
rect 12686 53106 12738 53118
rect 20526 53170 20578 53182
rect 20526 53106 20578 53118
rect 21534 53170 21586 53182
rect 21534 53106 21586 53118
rect 22430 53170 22482 53182
rect 22430 53106 22482 53118
rect 26910 53170 26962 53182
rect 26910 53106 26962 53118
rect 33966 53170 34018 53182
rect 33966 53106 34018 53118
rect 39566 53170 39618 53182
rect 39566 53106 39618 53118
rect 42814 53170 42866 53182
rect 42814 53106 42866 53118
rect 5406 53058 5458 53070
rect 5406 52994 5458 53006
rect 18286 53058 18338 53070
rect 18286 52994 18338 53006
rect 19854 53058 19906 53070
rect 19854 52994 19906 53006
rect 20414 53058 20466 53070
rect 20414 52994 20466 53006
rect 20638 53058 20690 53070
rect 20638 52994 20690 53006
rect 21982 53058 22034 53070
rect 21982 52994 22034 53006
rect 23774 53058 23826 53070
rect 23774 52994 23826 53006
rect 24670 53058 24722 53070
rect 24670 52994 24722 53006
rect 24894 53058 24946 53070
rect 24894 52994 24946 53006
rect 29038 53058 29090 53070
rect 29038 52994 29090 53006
rect 30270 53058 30322 53070
rect 30270 52994 30322 53006
rect 33742 53058 33794 53070
rect 33742 52994 33794 53006
rect 38334 53058 38386 53070
rect 38334 52994 38386 53006
rect 43262 53058 43314 53070
rect 43262 52994 43314 53006
rect 50654 53058 50706 53070
rect 50654 52994 50706 53006
rect 2270 52946 2322 52958
rect 2270 52882 2322 52894
rect 14814 52946 14866 52958
rect 14814 52882 14866 52894
rect 22206 52946 22258 52958
rect 22206 52882 22258 52894
rect 22542 52946 22594 52958
rect 23998 52946 24050 52958
rect 26798 52946 26850 52958
rect 23314 52894 23326 52946
rect 23378 52894 23390 52946
rect 23538 52894 23550 52946
rect 23602 52894 23614 52946
rect 26450 52894 26462 52946
rect 26514 52894 26526 52946
rect 22542 52882 22594 52894
rect 23998 52882 24050 52894
rect 26798 52882 26850 52894
rect 27022 52946 27074 52958
rect 27022 52882 27074 52894
rect 29710 52946 29762 52958
rect 33630 52946 33682 52958
rect 39342 52946 39394 52958
rect 30034 52894 30046 52946
rect 30098 52894 30110 52946
rect 36530 52894 36542 52946
rect 36594 52894 36606 52946
rect 37538 52894 37550 52946
rect 37602 52894 37614 52946
rect 29710 52882 29762 52894
rect 33630 52882 33682 52894
rect 39342 52882 39394 52894
rect 39566 52946 39618 52958
rect 39566 52882 39618 52894
rect 39790 52946 39842 52958
rect 39790 52882 39842 52894
rect 42590 52946 42642 52958
rect 42590 52882 42642 52894
rect 43038 52946 43090 52958
rect 53230 52946 53282 52958
rect 49858 52894 49870 52946
rect 49922 52894 49934 52946
rect 53554 52894 53566 52946
rect 53618 52894 53630 52946
rect 43038 52882 43090 52894
rect 53230 52882 53282 52894
rect 1822 52834 1874 52846
rect 1822 52770 1874 52782
rect 2718 52834 2770 52846
rect 2718 52770 2770 52782
rect 3502 52834 3554 52846
rect 3502 52770 3554 52782
rect 4174 52834 4226 52846
rect 4174 52770 4226 52782
rect 7646 52834 7698 52846
rect 7646 52770 7698 52782
rect 8094 52834 8146 52846
rect 8094 52770 8146 52782
rect 8542 52834 8594 52846
rect 8542 52770 8594 52782
rect 10894 52834 10946 52846
rect 10894 52770 10946 52782
rect 11342 52834 11394 52846
rect 11342 52770 11394 52782
rect 12238 52834 12290 52846
rect 12238 52770 12290 52782
rect 13134 52834 13186 52846
rect 13134 52770 13186 52782
rect 13918 52834 13970 52846
rect 13918 52770 13970 52782
rect 14366 52834 14418 52846
rect 14366 52770 14418 52782
rect 15374 52834 15426 52846
rect 15374 52770 15426 52782
rect 16046 52834 16098 52846
rect 16046 52770 16098 52782
rect 16494 52834 16546 52846
rect 16494 52770 16546 52782
rect 16942 52834 16994 52846
rect 16942 52770 16994 52782
rect 18958 52834 19010 52846
rect 18958 52770 19010 52782
rect 19518 52834 19570 52846
rect 23886 52834 23938 52846
rect 25678 52834 25730 52846
rect 22418 52782 22430 52834
rect 22482 52782 22494 52834
rect 24546 52782 24558 52834
rect 24610 52782 24622 52834
rect 19518 52770 19570 52782
rect 23886 52770 23938 52782
rect 25678 52770 25730 52782
rect 27470 52834 27522 52846
rect 27470 52770 27522 52782
rect 27918 52834 27970 52846
rect 27918 52770 27970 52782
rect 28366 52834 28418 52846
rect 40350 52834 40402 52846
rect 30146 52782 30158 52834
rect 30210 52782 30222 52834
rect 36642 52782 36654 52834
rect 36706 52782 36718 52834
rect 28366 52770 28418 52782
rect 40350 52770 40402 52782
rect 47742 52834 47794 52846
rect 53118 52834 53170 52846
rect 50082 52782 50094 52834
rect 50146 52782 50158 52834
rect 47742 52770 47794 52782
rect 53118 52770 53170 52782
rect 18062 52722 18114 52734
rect 5954 52670 5966 52722
rect 6018 52719 6030 52722
rect 8418 52719 8430 52722
rect 6018 52673 8430 52719
rect 6018 52670 6030 52673
rect 8418 52670 8430 52673
rect 8482 52670 8494 52722
rect 11778 52670 11790 52722
rect 11842 52719 11854 52722
rect 12114 52719 12126 52722
rect 11842 52673 12126 52719
rect 11842 52670 11854 52673
rect 12114 52670 12126 52673
rect 12178 52670 12190 52722
rect 13906 52670 13918 52722
rect 13970 52719 13982 52722
rect 14466 52719 14478 52722
rect 13970 52673 14478 52719
rect 13970 52670 13982 52673
rect 14466 52670 14478 52673
rect 14530 52670 14542 52722
rect 18062 52658 18114 52670
rect 18398 52722 18450 52734
rect 18722 52670 18734 52722
rect 18786 52719 18798 52722
rect 19954 52719 19966 52722
rect 18786 52673 19966 52719
rect 18786 52670 18798 52673
rect 19954 52670 19966 52673
rect 20018 52670 20030 52722
rect 18398 52658 18450 52670
rect 1344 52554 59024 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 59024 52554
rect 1344 52468 59024 52502
rect 25006 52386 25058 52398
rect 2482 52334 2494 52386
rect 2546 52383 2558 52386
rect 2706 52383 2718 52386
rect 2546 52337 2718 52383
rect 2546 52334 2558 52337
rect 2706 52334 2718 52337
rect 2770 52334 2782 52386
rect 40562 52334 40574 52386
rect 40626 52334 40638 52386
rect 25006 52322 25058 52334
rect 1822 52274 1874 52286
rect 1822 52210 1874 52222
rect 2270 52274 2322 52286
rect 2270 52210 2322 52222
rect 3054 52274 3106 52286
rect 3054 52210 3106 52222
rect 4286 52274 4338 52286
rect 4286 52210 4338 52222
rect 6078 52274 6130 52286
rect 6078 52210 6130 52222
rect 6526 52274 6578 52286
rect 6526 52210 6578 52222
rect 6974 52274 7026 52286
rect 6974 52210 7026 52222
rect 8094 52274 8146 52286
rect 8094 52210 8146 52222
rect 8542 52274 8594 52286
rect 8542 52210 8594 52222
rect 9438 52274 9490 52286
rect 9438 52210 9490 52222
rect 13806 52274 13858 52286
rect 13806 52210 13858 52222
rect 14254 52274 14306 52286
rect 19966 52274 20018 52286
rect 17154 52222 17166 52274
rect 17218 52222 17230 52274
rect 18386 52222 18398 52274
rect 18450 52222 18462 52274
rect 19394 52222 19406 52274
rect 19458 52222 19470 52274
rect 14254 52210 14306 52222
rect 19966 52210 20018 52222
rect 20526 52274 20578 52286
rect 20526 52210 20578 52222
rect 22094 52274 22146 52286
rect 22094 52210 22146 52222
rect 22766 52274 22818 52286
rect 22766 52210 22818 52222
rect 24334 52274 24386 52286
rect 24334 52210 24386 52222
rect 26350 52274 26402 52286
rect 26350 52210 26402 52222
rect 30606 52274 30658 52286
rect 30606 52210 30658 52222
rect 33070 52274 33122 52286
rect 33070 52210 33122 52222
rect 35086 52274 35138 52286
rect 46062 52274 46114 52286
rect 39890 52222 39902 52274
rect 39954 52222 39966 52274
rect 35086 52210 35138 52222
rect 46062 52210 46114 52222
rect 53454 52274 53506 52286
rect 53454 52210 53506 52222
rect 4846 52162 4898 52174
rect 4846 52098 4898 52110
rect 9102 52162 9154 52174
rect 12462 52162 12514 52174
rect 10546 52110 10558 52162
rect 10610 52110 10622 52162
rect 11106 52110 11118 52162
rect 11170 52110 11182 52162
rect 11666 52110 11678 52162
rect 11730 52110 11742 52162
rect 9102 52098 9154 52110
rect 12462 52098 12514 52110
rect 13022 52162 13074 52174
rect 13022 52098 13074 52110
rect 15150 52162 15202 52174
rect 20862 52162 20914 52174
rect 15698 52110 15710 52162
rect 15762 52110 15774 52162
rect 16034 52110 16046 52162
rect 16098 52110 16110 52162
rect 18274 52110 18286 52162
rect 18338 52110 18350 52162
rect 15150 52098 15202 52110
rect 20862 52098 20914 52110
rect 21534 52162 21586 52174
rect 21534 52098 21586 52110
rect 22542 52162 22594 52174
rect 22542 52098 22594 52110
rect 22990 52162 23042 52174
rect 22990 52098 23042 52110
rect 23214 52162 23266 52174
rect 23214 52098 23266 52110
rect 23774 52162 23826 52174
rect 23774 52098 23826 52110
rect 24222 52162 24274 52174
rect 28926 52162 28978 52174
rect 24658 52110 24670 52162
rect 24722 52159 24734 52162
rect 24882 52159 24894 52162
rect 24722 52113 24894 52159
rect 24722 52110 24734 52113
rect 24882 52110 24894 52113
rect 24946 52110 24958 52162
rect 24222 52098 24274 52110
rect 28926 52098 28978 52110
rect 29710 52162 29762 52174
rect 31166 52162 31218 52174
rect 41134 52162 41186 52174
rect 30146 52110 30158 52162
rect 30210 52110 30222 52162
rect 34626 52110 34638 52162
rect 34690 52110 34702 52162
rect 39778 52110 39790 52162
rect 39842 52110 39854 52162
rect 29710 52098 29762 52110
rect 31166 52098 31218 52110
rect 41134 52098 41186 52110
rect 46174 52162 46226 52174
rect 46174 52098 46226 52110
rect 46622 52162 46674 52174
rect 46622 52098 46674 52110
rect 52782 52162 52834 52174
rect 52782 52098 52834 52110
rect 53566 52162 53618 52174
rect 53890 52110 53902 52162
rect 53954 52110 53966 52162
rect 53566 52098 53618 52110
rect 14814 52050 14866 52062
rect 10434 51998 10446 52050
rect 10498 51998 10510 52050
rect 10882 51998 10894 52050
rect 10946 51998 10958 52050
rect 14814 51986 14866 51998
rect 14926 52050 14978 52062
rect 14926 51986 14978 51998
rect 26910 52050 26962 52062
rect 26910 51986 26962 51998
rect 27134 52050 27186 52062
rect 27134 51986 27186 51998
rect 27358 52050 27410 52062
rect 27358 51986 27410 51998
rect 27470 52050 27522 52062
rect 45950 52050 46002 52062
rect 33282 51998 33294 52050
rect 33346 51998 33358 52050
rect 27470 51986 27522 51998
rect 45950 51986 46002 51998
rect 52446 52050 52498 52062
rect 52446 51986 52498 51998
rect 2606 51938 2658 51950
rect 2606 51874 2658 51886
rect 3950 51938 4002 51950
rect 3950 51874 4002 51886
rect 5630 51938 5682 51950
rect 5630 51874 5682 51886
rect 7646 51938 7698 51950
rect 7646 51874 7698 51886
rect 23102 51938 23154 51950
rect 23102 51874 23154 51886
rect 24446 51938 24498 51950
rect 24446 51874 24498 51886
rect 25118 51938 25170 51950
rect 25118 51874 25170 51886
rect 25230 51938 25282 51950
rect 25230 51874 25282 51886
rect 26014 51938 26066 51950
rect 26014 51874 26066 51886
rect 27918 51938 27970 51950
rect 27918 51874 27970 51886
rect 28478 51938 28530 51950
rect 28478 51874 28530 51886
rect 32174 51938 32226 51950
rect 32174 51874 32226 51886
rect 52558 51938 52610 51950
rect 52558 51874 52610 51886
rect 1344 51770 59024 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 59024 51770
rect 1344 51684 59024 51718
rect 2270 51602 2322 51614
rect 2270 51538 2322 51550
rect 3166 51602 3218 51614
rect 3166 51538 3218 51550
rect 4846 51602 4898 51614
rect 4846 51538 4898 51550
rect 5294 51602 5346 51614
rect 5294 51538 5346 51550
rect 5742 51602 5794 51614
rect 5742 51538 5794 51550
rect 12462 51602 12514 51614
rect 12462 51538 12514 51550
rect 15710 51602 15762 51614
rect 15710 51538 15762 51550
rect 15822 51602 15874 51614
rect 15822 51538 15874 51550
rect 17838 51602 17890 51614
rect 17838 51538 17890 51550
rect 18846 51602 18898 51614
rect 18846 51538 18898 51550
rect 21198 51602 21250 51614
rect 21198 51538 21250 51550
rect 22094 51602 22146 51614
rect 29150 51602 29202 51614
rect 23538 51550 23550 51602
rect 23602 51550 23614 51602
rect 22094 51538 22146 51550
rect 29150 51538 29202 51550
rect 33854 51602 33906 51614
rect 33854 51538 33906 51550
rect 36654 51602 36706 51614
rect 36654 51538 36706 51550
rect 37550 51602 37602 51614
rect 37550 51538 37602 51550
rect 42142 51602 42194 51614
rect 55122 51550 55134 51602
rect 55186 51550 55198 51602
rect 42142 51538 42194 51550
rect 8878 51490 8930 51502
rect 19406 51490 19458 51502
rect 13010 51438 13022 51490
rect 13074 51438 13086 51490
rect 8878 51426 8930 51438
rect 19406 51426 19458 51438
rect 22990 51490 23042 51502
rect 22990 51426 23042 51438
rect 25902 51490 25954 51502
rect 25902 51426 25954 51438
rect 28254 51490 28306 51502
rect 28254 51426 28306 51438
rect 29374 51490 29426 51502
rect 29374 51426 29426 51438
rect 39454 51490 39506 51502
rect 39454 51426 39506 51438
rect 42254 51490 42306 51502
rect 47854 51490 47906 51502
rect 45938 51438 45950 51490
rect 46002 51438 46014 51490
rect 42254 51426 42306 51438
rect 47854 51426 47906 51438
rect 52334 51490 52386 51502
rect 52334 51426 52386 51438
rect 3614 51378 3666 51390
rect 3614 51314 3666 51326
rect 6190 51378 6242 51390
rect 6190 51314 6242 51326
rect 6638 51378 6690 51390
rect 6638 51314 6690 51326
rect 6862 51378 6914 51390
rect 6862 51314 6914 51326
rect 7534 51378 7586 51390
rect 7534 51314 7586 51326
rect 7758 51378 7810 51390
rect 7758 51314 7810 51326
rect 7982 51378 8034 51390
rect 7982 51314 8034 51326
rect 8654 51378 8706 51390
rect 8654 51314 8706 51326
rect 8990 51378 9042 51390
rect 10894 51378 10946 51390
rect 10434 51326 10446 51378
rect 10498 51326 10510 51378
rect 10658 51326 10670 51378
rect 10722 51326 10734 51378
rect 8990 51314 9042 51326
rect 10894 51314 10946 51326
rect 11118 51378 11170 51390
rect 15598 51378 15650 51390
rect 18286 51378 18338 51390
rect 23214 51378 23266 51390
rect 11330 51326 11342 51378
rect 11394 51326 11406 51378
rect 14242 51326 14254 51378
rect 14306 51326 14318 51378
rect 15922 51326 15934 51378
rect 15986 51326 15998 51378
rect 18610 51326 18622 51378
rect 18674 51326 18686 51378
rect 20066 51326 20078 51378
rect 20130 51326 20142 51378
rect 11118 51314 11170 51326
rect 15598 51314 15650 51326
rect 18286 51314 18338 51326
rect 23214 51314 23266 51326
rect 24334 51378 24386 51390
rect 24334 51314 24386 51326
rect 24558 51378 24610 51390
rect 24558 51314 24610 51326
rect 25006 51378 25058 51390
rect 25006 51314 25058 51326
rect 26126 51378 26178 51390
rect 29486 51378 29538 51390
rect 32622 51378 32674 51390
rect 27794 51326 27806 51378
rect 27858 51326 27870 51378
rect 30258 51326 30270 51378
rect 30322 51326 30334 51378
rect 32386 51326 32398 51378
rect 32450 51326 32462 51378
rect 26126 51314 26178 51326
rect 29486 51314 29538 51326
rect 32622 51314 32674 51326
rect 33742 51378 33794 51390
rect 33742 51314 33794 51326
rect 33966 51378 34018 51390
rect 36206 51378 36258 51390
rect 34066 51326 34078 51378
rect 34130 51326 34142 51378
rect 33966 51314 34018 51326
rect 36206 51314 36258 51326
rect 36542 51378 36594 51390
rect 36542 51314 36594 51326
rect 36878 51378 36930 51390
rect 39342 51378 39394 51390
rect 44046 51378 44098 51390
rect 37314 51326 37326 51378
rect 37378 51326 37390 51378
rect 38994 51326 39006 51378
rect 39058 51326 39070 51378
rect 43138 51326 43150 51378
rect 43202 51326 43214 51378
rect 36878 51314 36930 51326
rect 39342 51314 39394 51326
rect 44046 51314 44098 51326
rect 44942 51378 44994 51390
rect 47170 51326 47182 51378
rect 47234 51326 47246 51378
rect 51874 51326 51886 51378
rect 51938 51326 51950 51378
rect 44942 51314 44994 51326
rect 1934 51266 1986 51278
rect 1934 51202 1986 51214
rect 2718 51266 2770 51278
rect 2718 51202 2770 51214
rect 4062 51266 4114 51278
rect 4062 51202 4114 51214
rect 6750 51266 6802 51278
rect 6750 51202 6802 51214
rect 7870 51266 7922 51278
rect 16942 51266 16994 51278
rect 13906 51214 13918 51266
rect 13970 51214 13982 51266
rect 7870 51202 7922 51214
rect 16942 51202 16994 51214
rect 18958 51266 19010 51278
rect 21646 51266 21698 51278
rect 19730 51214 19742 51266
rect 19794 51214 19806 51266
rect 18958 51202 19010 51214
rect 21646 51202 21698 51214
rect 24446 51266 24498 51278
rect 28702 51266 28754 51278
rect 31054 51266 31106 51278
rect 27458 51214 27470 51266
rect 27522 51214 27534 51266
rect 30706 51214 30718 51266
rect 30770 51214 30782 51266
rect 24446 51202 24498 51214
rect 28702 51202 28754 51214
rect 31054 51202 31106 51214
rect 32734 51266 32786 51278
rect 32734 51202 32786 51214
rect 34638 51266 34690 51278
rect 34638 51202 34690 51214
rect 39902 51266 39954 51278
rect 45838 51266 45890 51278
rect 55694 51266 55746 51278
rect 43250 51214 43262 51266
rect 43314 51214 43326 51266
rect 51538 51214 51550 51266
rect 51602 51214 51614 51266
rect 39902 51202 39954 51214
rect 45838 51202 45890 51214
rect 55694 51202 55746 51214
rect 56254 51266 56306 51278
rect 56254 51202 56306 51214
rect 58046 51266 58098 51278
rect 58046 51202 58098 51214
rect 58382 51266 58434 51278
rect 58382 51202 58434 51214
rect 16270 51154 16322 51166
rect 26462 51154 26514 51166
rect 1698 51102 1710 51154
rect 1762 51151 1774 51154
rect 2706 51151 2718 51154
rect 1762 51105 2718 51151
rect 1762 51102 1774 51105
rect 2706 51102 2718 51105
rect 2770 51102 2782 51154
rect 11554 51102 11566 51154
rect 11618 51102 11630 51154
rect 12114 51102 12126 51154
rect 12178 51151 12190 51154
rect 12786 51151 12798 51154
rect 12178 51105 12798 51151
rect 12178 51102 12190 51105
rect 12786 51102 12798 51105
rect 12850 51102 12862 51154
rect 21186 51102 21198 51154
rect 21250 51151 21262 51154
rect 22194 51151 22206 51154
rect 21250 51105 22206 51151
rect 21250 51102 21262 51105
rect 22194 51102 22206 51105
rect 22258 51102 22270 51154
rect 16270 51090 16322 51102
rect 26462 51090 26514 51102
rect 34414 51154 34466 51166
rect 34414 51090 34466 51102
rect 37662 51154 37714 51166
rect 37662 51090 37714 51102
rect 42030 51154 42082 51166
rect 42030 51090 42082 51102
rect 45054 51154 45106 51166
rect 45054 51090 45106 51102
rect 55470 51154 55522 51166
rect 57698 51102 57710 51154
rect 57762 51151 57774 51154
rect 58370 51151 58382 51154
rect 57762 51105 58382 51151
rect 57762 51102 57774 51105
rect 58370 51102 58382 51105
rect 58434 51102 58446 51154
rect 55470 51090 55522 51102
rect 1344 50986 59024 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 59024 50986
rect 1344 50900 59024 50934
rect 6302 50818 6354 50830
rect 6302 50754 6354 50766
rect 12126 50818 12178 50830
rect 12126 50754 12178 50766
rect 16382 50818 16434 50830
rect 16382 50754 16434 50766
rect 16718 50818 16770 50830
rect 31278 50818 31330 50830
rect 33406 50818 33458 50830
rect 21858 50766 21870 50818
rect 21922 50815 21934 50818
rect 23650 50815 23662 50818
rect 21922 50769 23662 50815
rect 21922 50766 21934 50769
rect 23650 50766 23662 50769
rect 23714 50766 23726 50818
rect 32050 50766 32062 50818
rect 32114 50815 32126 50818
rect 32498 50815 32510 50818
rect 32114 50769 32510 50815
rect 32114 50766 32126 50769
rect 32498 50766 32510 50769
rect 32562 50766 32574 50818
rect 16718 50754 16770 50766
rect 31278 50754 31330 50766
rect 33406 50754 33458 50766
rect 39342 50818 39394 50830
rect 41918 50818 41970 50830
rect 46286 50818 46338 50830
rect 39666 50766 39678 50818
rect 39730 50766 39742 50818
rect 42914 50766 42926 50818
rect 42978 50766 42990 50818
rect 39342 50754 39394 50766
rect 41918 50754 41970 50766
rect 46286 50754 46338 50766
rect 51550 50818 51602 50830
rect 51550 50754 51602 50766
rect 55918 50818 55970 50830
rect 55918 50754 55970 50766
rect 58158 50818 58210 50830
rect 58158 50754 58210 50766
rect 2606 50706 2658 50718
rect 2606 50642 2658 50654
rect 2942 50706 2994 50718
rect 2942 50642 2994 50654
rect 4510 50706 4562 50718
rect 4510 50642 4562 50654
rect 6862 50706 6914 50718
rect 6862 50642 6914 50654
rect 7758 50706 7810 50718
rect 7758 50642 7810 50654
rect 12238 50706 12290 50718
rect 12238 50642 12290 50654
rect 12910 50706 12962 50718
rect 18174 50706 18226 50718
rect 21870 50706 21922 50718
rect 13906 50654 13918 50706
rect 13970 50654 13982 50706
rect 19170 50654 19182 50706
rect 19234 50654 19246 50706
rect 19954 50654 19966 50706
rect 20018 50654 20030 50706
rect 12910 50642 12962 50654
rect 18174 50642 18226 50654
rect 21870 50642 21922 50654
rect 22318 50706 22370 50718
rect 22318 50642 22370 50654
rect 23662 50706 23714 50718
rect 27358 50706 27410 50718
rect 30606 50706 30658 50718
rect 27010 50654 27022 50706
rect 27074 50654 27086 50706
rect 27906 50654 27918 50706
rect 27970 50654 27982 50706
rect 30146 50654 30158 50706
rect 30210 50654 30222 50706
rect 23662 50642 23714 50654
rect 27358 50642 27410 50654
rect 30606 50642 30658 50654
rect 32510 50706 32562 50718
rect 38558 50706 38610 50718
rect 41806 50706 41858 50718
rect 50654 50706 50706 50718
rect 36418 50654 36430 50706
rect 36482 50654 36494 50706
rect 37650 50654 37662 50706
rect 37714 50654 37726 50706
rect 40226 50654 40238 50706
rect 40290 50654 40302 50706
rect 43138 50654 43150 50706
rect 43202 50654 43214 50706
rect 46050 50654 46062 50706
rect 46114 50654 46126 50706
rect 48514 50654 48526 50706
rect 48578 50654 48590 50706
rect 32510 50642 32562 50654
rect 38558 50642 38610 50654
rect 41806 50642 41858 50654
rect 50654 50642 50706 50654
rect 2158 50594 2210 50606
rect 2158 50530 2210 50542
rect 4062 50594 4114 50606
rect 6974 50594 7026 50606
rect 14030 50594 14082 50606
rect 14478 50594 14530 50606
rect 6626 50542 6638 50594
rect 6690 50542 6702 50594
rect 9090 50542 9102 50594
rect 9154 50542 9166 50594
rect 9874 50542 9886 50594
rect 9938 50542 9950 50594
rect 10882 50542 10894 50594
rect 10946 50542 10958 50594
rect 14130 50542 14142 50594
rect 14194 50542 14206 50594
rect 4062 50530 4114 50542
rect 6974 50530 7026 50542
rect 14030 50530 14082 50542
rect 14478 50530 14530 50542
rect 14702 50594 14754 50606
rect 14702 50530 14754 50542
rect 15150 50594 15202 50606
rect 23326 50594 23378 50606
rect 20290 50542 20302 50594
rect 20354 50542 20366 50594
rect 15150 50530 15202 50542
rect 23326 50530 23378 50542
rect 24558 50594 24610 50606
rect 24558 50530 24610 50542
rect 24894 50594 24946 50606
rect 31390 50594 31442 50606
rect 36766 50594 36818 50606
rect 39118 50594 39170 50606
rect 26898 50542 26910 50594
rect 26962 50542 26974 50594
rect 29922 50542 29934 50594
rect 29986 50542 29998 50594
rect 33394 50542 33406 50594
rect 33458 50542 33470 50594
rect 36306 50542 36318 50594
rect 36370 50542 36382 50594
rect 37874 50542 37886 50594
rect 37938 50542 37950 50594
rect 24894 50530 24946 50542
rect 31390 50530 31442 50542
rect 36766 50530 36818 50542
rect 39118 50530 39170 50542
rect 40574 50594 40626 50606
rect 40574 50530 40626 50542
rect 41022 50594 41074 50606
rect 46734 50594 46786 50606
rect 41570 50542 41582 50594
rect 41634 50542 41646 50594
rect 43362 50542 43374 50594
rect 43426 50542 43438 50594
rect 41022 50530 41074 50542
rect 46734 50530 46786 50542
rect 47070 50594 47122 50606
rect 54462 50594 54514 50606
rect 49970 50542 49982 50594
rect 50034 50542 50046 50594
rect 54226 50542 54238 50594
rect 54290 50542 54302 50594
rect 47070 50530 47122 50542
rect 54462 50530 54514 50542
rect 56142 50594 56194 50606
rect 56814 50594 56866 50606
rect 56354 50542 56366 50594
rect 56418 50542 56430 50594
rect 56142 50530 56194 50542
rect 56814 50530 56866 50542
rect 57262 50594 57314 50606
rect 57262 50530 57314 50542
rect 57486 50594 57538 50606
rect 57486 50530 57538 50542
rect 5070 50482 5122 50494
rect 5070 50418 5122 50430
rect 7646 50482 7698 50494
rect 7646 50418 7698 50430
rect 7870 50482 7922 50494
rect 12350 50482 12402 50494
rect 8754 50430 8766 50482
rect 8818 50430 8830 50482
rect 9762 50430 9774 50482
rect 9826 50430 9838 50482
rect 7870 50418 7922 50430
rect 12350 50418 12402 50430
rect 13806 50482 13858 50494
rect 13806 50418 13858 50430
rect 15598 50482 15650 50494
rect 15598 50418 15650 50430
rect 15822 50482 15874 50494
rect 15822 50418 15874 50430
rect 16494 50482 16546 50494
rect 16494 50418 16546 50430
rect 20862 50482 20914 50494
rect 20862 50418 20914 50430
rect 25118 50482 25170 50494
rect 25118 50418 25170 50430
rect 25790 50482 25842 50494
rect 25790 50418 25842 50430
rect 28030 50482 28082 50494
rect 28030 50418 28082 50430
rect 28254 50482 28306 50494
rect 28254 50418 28306 50430
rect 28814 50482 28866 50494
rect 28814 50418 28866 50430
rect 31278 50482 31330 50494
rect 31278 50418 31330 50430
rect 32062 50482 32114 50494
rect 32062 50418 32114 50430
rect 33070 50482 33122 50494
rect 33070 50418 33122 50430
rect 35198 50482 35250 50494
rect 35198 50418 35250 50430
rect 40350 50482 40402 50494
rect 51774 50482 51826 50494
rect 48962 50430 48974 50482
rect 49026 50430 49038 50482
rect 40350 50418 40402 50430
rect 51774 50418 51826 50430
rect 54126 50482 54178 50494
rect 54126 50418 54178 50430
rect 58046 50482 58098 50494
rect 58046 50418 58098 50430
rect 3502 50370 3554 50382
rect 3502 50306 3554 50318
rect 5742 50370 5794 50382
rect 5742 50306 5794 50318
rect 6750 50370 6802 50382
rect 6750 50306 6802 50318
rect 11006 50370 11058 50382
rect 11006 50306 11058 50318
rect 11342 50370 11394 50382
rect 11342 50306 11394 50318
rect 15486 50370 15538 50382
rect 15486 50306 15538 50318
rect 17614 50370 17666 50382
rect 17614 50306 17666 50318
rect 18734 50370 18786 50382
rect 18734 50306 18786 50318
rect 22766 50370 22818 50382
rect 22766 50306 22818 50318
rect 25006 50370 25058 50382
rect 25006 50306 25058 50318
rect 33854 50370 33906 50382
rect 33854 50306 33906 50318
rect 34302 50370 34354 50382
rect 34302 50306 34354 50318
rect 34750 50370 34802 50382
rect 34750 50306 34802 50318
rect 46062 50370 46114 50382
rect 46062 50306 46114 50318
rect 46958 50370 47010 50382
rect 53566 50370 53618 50382
rect 51202 50318 51214 50370
rect 51266 50318 51278 50370
rect 46958 50306 47010 50318
rect 53566 50306 53618 50318
rect 56254 50370 56306 50382
rect 56254 50306 56306 50318
rect 57150 50370 57202 50382
rect 57150 50306 57202 50318
rect 58158 50370 58210 50382
rect 58158 50306 58210 50318
rect 1344 50202 59024 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 59024 50202
rect 1344 50116 59024 50150
rect 3390 50034 3442 50046
rect 3390 49970 3442 49982
rect 4958 50034 5010 50046
rect 4958 49970 5010 49982
rect 5630 50034 5682 50046
rect 5630 49970 5682 49982
rect 8318 50034 8370 50046
rect 8318 49970 8370 49982
rect 10222 50034 10274 50046
rect 10222 49970 10274 49982
rect 10558 50034 10610 50046
rect 10558 49970 10610 49982
rect 11454 50034 11506 50046
rect 11454 49970 11506 49982
rect 11678 50034 11730 50046
rect 11678 49970 11730 49982
rect 12686 50034 12738 50046
rect 15710 50034 15762 50046
rect 14242 49982 14254 50034
rect 14306 49982 14318 50034
rect 12686 49970 12738 49982
rect 15710 49970 15762 49982
rect 17838 50034 17890 50046
rect 17838 49970 17890 49982
rect 18062 50034 18114 50046
rect 18062 49970 18114 49982
rect 19294 50034 19346 50046
rect 19294 49970 19346 49982
rect 25678 50034 25730 50046
rect 29598 50034 29650 50046
rect 26674 49982 26686 50034
rect 26738 49982 26750 50034
rect 25678 49970 25730 49982
rect 29598 49970 29650 49982
rect 30382 50034 30434 50046
rect 30382 49970 30434 49982
rect 30494 50034 30546 50046
rect 30494 49970 30546 49982
rect 31950 50034 32002 50046
rect 31950 49970 32002 49982
rect 32622 50034 32674 50046
rect 39790 50034 39842 50046
rect 45950 50034 46002 50046
rect 36082 49982 36094 50034
rect 36146 49982 36158 50034
rect 43250 49982 43262 50034
rect 43314 49982 43326 50034
rect 32622 49970 32674 49982
rect 39790 49970 39842 49982
rect 45950 49970 46002 49982
rect 52558 50034 52610 50046
rect 52558 49970 52610 49982
rect 53118 50034 53170 50046
rect 53118 49970 53170 49982
rect 57598 50034 57650 50046
rect 57598 49970 57650 49982
rect 57822 50034 57874 50046
rect 57822 49970 57874 49982
rect 4734 49922 4786 49934
rect 4734 49858 4786 49870
rect 7982 49922 8034 49934
rect 7982 49858 8034 49870
rect 12462 49922 12514 49934
rect 12462 49858 12514 49870
rect 17726 49922 17778 49934
rect 17726 49858 17778 49870
rect 19854 49922 19906 49934
rect 19854 49858 19906 49870
rect 29486 49922 29538 49934
rect 29486 49858 29538 49870
rect 31726 49922 31778 49934
rect 31726 49858 31778 49870
rect 39678 49922 39730 49934
rect 39678 49858 39730 49870
rect 39902 49922 39954 49934
rect 39902 49858 39954 49870
rect 40350 49922 40402 49934
rect 40350 49858 40402 49870
rect 58382 49922 58434 49934
rect 58382 49858 58434 49870
rect 58494 49922 58546 49934
rect 58494 49858 58546 49870
rect 2382 49810 2434 49822
rect 2382 49746 2434 49758
rect 3950 49810 4002 49822
rect 8318 49810 8370 49822
rect 6962 49758 6974 49810
rect 7026 49758 7038 49810
rect 3950 49746 4002 49758
rect 8318 49746 8370 49758
rect 8542 49810 8594 49822
rect 8542 49746 8594 49758
rect 10110 49810 10162 49822
rect 11790 49810 11842 49822
rect 10322 49758 10334 49810
rect 10386 49758 10398 49810
rect 10110 49746 10162 49758
rect 11790 49746 11842 49758
rect 12350 49810 12402 49822
rect 12350 49746 12402 49758
rect 13134 49810 13186 49822
rect 13134 49746 13186 49758
rect 13358 49810 13410 49822
rect 13358 49746 13410 49758
rect 13806 49810 13858 49822
rect 13806 49746 13858 49758
rect 18510 49810 18562 49822
rect 27246 49810 27298 49822
rect 20514 49758 20526 49810
rect 20578 49758 20590 49810
rect 20738 49758 20750 49810
rect 20802 49758 20814 49810
rect 23538 49758 23550 49810
rect 23602 49758 23614 49810
rect 18510 49746 18562 49758
rect 27246 49746 27298 49758
rect 27918 49810 27970 49822
rect 27918 49746 27970 49758
rect 29710 49810 29762 49822
rect 29710 49746 29762 49758
rect 30270 49810 30322 49822
rect 30270 49746 30322 49758
rect 30942 49810 30994 49822
rect 30942 49746 30994 49758
rect 31614 49810 31666 49822
rect 31614 49746 31666 49758
rect 32398 49810 32450 49822
rect 34526 49810 34578 49822
rect 45726 49810 45778 49822
rect 33954 49758 33966 49810
rect 34018 49758 34030 49810
rect 42018 49758 42030 49810
rect 42082 49758 42094 49810
rect 32398 49746 32450 49758
rect 34526 49746 34578 49758
rect 45726 49746 45778 49758
rect 46062 49810 46114 49822
rect 46062 49746 46114 49758
rect 48190 49810 48242 49822
rect 48190 49746 48242 49758
rect 49534 49810 49586 49822
rect 52334 49810 52386 49822
rect 52210 49758 52222 49810
rect 52274 49758 52286 49810
rect 49534 49746 49586 49758
rect 52334 49746 52386 49758
rect 55470 49810 55522 49822
rect 55470 49746 55522 49758
rect 55694 49810 55746 49822
rect 55694 49746 55746 49758
rect 57486 49810 57538 49822
rect 57486 49746 57538 49758
rect 58158 49810 58210 49822
rect 58158 49746 58210 49758
rect 2046 49698 2098 49710
rect 2046 49634 2098 49646
rect 2942 49698 2994 49710
rect 8990 49698 9042 49710
rect 6066 49646 6078 49698
rect 6130 49646 6142 49698
rect 7298 49646 7310 49698
rect 7362 49646 7374 49698
rect 2942 49634 2994 49646
rect 8990 49634 9042 49646
rect 13246 49698 13298 49710
rect 13246 49634 13298 49646
rect 14814 49698 14866 49710
rect 16494 49698 16546 49710
rect 15810 49646 15822 49698
rect 15874 49646 15886 49698
rect 14814 49634 14866 49646
rect 16494 49634 16546 49646
rect 16942 49698 16994 49710
rect 26126 49698 26178 49710
rect 22530 49646 22542 49698
rect 22594 49646 22606 49698
rect 23762 49646 23774 49698
rect 23826 49646 23838 49698
rect 24770 49646 24782 49698
rect 24834 49646 24846 49698
rect 16942 49634 16994 49646
rect 26126 49634 26178 49646
rect 27022 49698 27074 49710
rect 27022 49634 27074 49646
rect 28366 49698 28418 49710
rect 28366 49634 28418 49646
rect 28814 49698 28866 49710
rect 28814 49634 28866 49646
rect 34638 49698 34690 49710
rect 34638 49634 34690 49646
rect 35534 49698 35586 49710
rect 35534 49634 35586 49646
rect 35758 49698 35810 49710
rect 35758 49634 35810 49646
rect 36542 49698 36594 49710
rect 36542 49634 36594 49646
rect 37102 49698 37154 49710
rect 37102 49634 37154 49646
rect 37550 49698 37602 49710
rect 42590 49698 42642 49710
rect 41906 49646 41918 49698
rect 41970 49646 41982 49698
rect 37550 49634 37602 49646
rect 42590 49634 42642 49646
rect 43822 49698 43874 49710
rect 43822 49634 43874 49646
rect 49758 49698 49810 49710
rect 49758 49634 49810 49646
rect 50878 49698 50930 49710
rect 50878 49634 50930 49646
rect 51438 49698 51490 49710
rect 51438 49634 51490 49646
rect 52446 49698 52498 49710
rect 52446 49634 52498 49646
rect 53790 49698 53842 49710
rect 53790 49634 53842 49646
rect 55918 49698 55970 49710
rect 55918 49634 55970 49646
rect 56702 49698 56754 49710
rect 56702 49634 56754 49646
rect 5070 49586 5122 49598
rect 2034 49534 2046 49586
rect 2098 49583 2110 49586
rect 3154 49583 3166 49586
rect 2098 49537 3166 49583
rect 2098 49534 2110 49537
rect 3154 49534 3166 49537
rect 3218 49534 3230 49586
rect 5070 49522 5122 49534
rect 10894 49586 10946 49598
rect 10894 49522 10946 49534
rect 11006 49586 11058 49598
rect 11006 49522 11058 49534
rect 14590 49586 14642 49598
rect 14590 49522 14642 49534
rect 15486 49586 15538 49598
rect 32734 49586 32786 49598
rect 25554 49534 25566 49586
rect 25618 49583 25630 49586
rect 26114 49583 26126 49586
rect 25618 49537 26126 49583
rect 25618 49534 25630 49537
rect 26114 49534 26126 49537
rect 26178 49534 26190 49586
rect 15486 49522 15538 49534
rect 32734 49522 32786 49534
rect 43598 49586 43650 49598
rect 43598 49522 43650 49534
rect 48414 49586 48466 49598
rect 48414 49522 48466 49534
rect 48750 49586 48802 49598
rect 51886 49586 51938 49598
rect 50082 49534 50094 49586
rect 50146 49534 50158 49586
rect 48750 49522 48802 49534
rect 51886 49522 51938 49534
rect 56366 49586 56418 49598
rect 56366 49522 56418 49534
rect 1344 49418 59024 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 59024 49418
rect 1344 49332 59024 49366
rect 5742 49250 5794 49262
rect 42142 49250 42194 49262
rect 1922 49198 1934 49250
rect 1986 49247 1998 49250
rect 2594 49247 2606 49250
rect 1986 49201 2606 49247
rect 1986 49198 1998 49201
rect 2594 49198 2606 49201
rect 2658 49247 2670 49250
rect 3042 49247 3054 49250
rect 2658 49201 3054 49247
rect 2658 49198 2670 49201
rect 3042 49198 3054 49201
rect 3106 49198 3118 49250
rect 13906 49198 13918 49250
rect 13970 49247 13982 49250
rect 14466 49247 14478 49250
rect 13970 49201 14478 49247
rect 13970 49198 13982 49201
rect 14466 49198 14478 49201
rect 14530 49198 14542 49250
rect 22866 49198 22878 49250
rect 22930 49198 22942 49250
rect 30706 49198 30718 49250
rect 30770 49198 30782 49250
rect 5742 49186 5794 49198
rect 42142 49186 42194 49198
rect 44606 49250 44658 49262
rect 52670 49250 52722 49262
rect 47170 49198 47182 49250
rect 47234 49198 47246 49250
rect 44606 49186 44658 49198
rect 52670 49186 52722 49198
rect 55470 49250 55522 49262
rect 55470 49186 55522 49198
rect 1934 49138 1986 49150
rect 1934 49074 1986 49086
rect 3838 49138 3890 49150
rect 3838 49074 3890 49086
rect 4958 49138 5010 49150
rect 4958 49074 5010 49086
rect 7310 49138 7362 49150
rect 7310 49074 7362 49086
rect 9214 49138 9266 49150
rect 12350 49138 12402 49150
rect 11442 49086 11454 49138
rect 11506 49086 11518 49138
rect 9214 49074 9266 49086
rect 12350 49074 12402 49086
rect 13918 49138 13970 49150
rect 13918 49074 13970 49086
rect 14366 49138 14418 49150
rect 14366 49074 14418 49086
rect 16942 49138 16994 49150
rect 16942 49074 16994 49086
rect 17390 49138 17442 49150
rect 26350 49138 26402 49150
rect 18386 49086 18398 49138
rect 18450 49086 18462 49138
rect 20850 49086 20862 49138
rect 20914 49086 20926 49138
rect 22642 49086 22654 49138
rect 22706 49086 22718 49138
rect 24882 49086 24894 49138
rect 24946 49086 24958 49138
rect 17390 49074 17442 49086
rect 26350 49074 26402 49086
rect 27918 49138 27970 49150
rect 27918 49074 27970 49086
rect 28366 49138 28418 49150
rect 28366 49074 28418 49086
rect 28814 49138 28866 49150
rect 36542 49138 36594 49150
rect 30482 49086 30494 49138
rect 30546 49086 30558 49138
rect 35746 49086 35758 49138
rect 35810 49086 35822 49138
rect 28814 49074 28866 49086
rect 36542 49074 36594 49086
rect 38334 49138 38386 49150
rect 49534 49138 49586 49150
rect 54126 49138 54178 49150
rect 46722 49086 46734 49138
rect 46786 49086 46798 49138
rect 51762 49086 51774 49138
rect 51826 49086 51838 49138
rect 56466 49086 56478 49138
rect 56530 49086 56542 49138
rect 57026 49086 57038 49138
rect 57090 49086 57102 49138
rect 38334 49074 38386 49086
rect 49534 49074 49586 49086
rect 54126 49074 54178 49086
rect 9886 49026 9938 49038
rect 9886 48962 9938 48974
rect 9998 49026 10050 49038
rect 9998 48962 10050 48974
rect 10334 49026 10386 49038
rect 10334 48962 10386 48974
rect 12126 49026 12178 49038
rect 12126 48962 12178 48974
rect 12798 49026 12850 49038
rect 12798 48962 12850 48974
rect 14926 49026 14978 49038
rect 14926 48962 14978 48974
rect 15262 49026 15314 49038
rect 15262 48962 15314 48974
rect 15598 49026 15650 49038
rect 15598 48962 15650 48974
rect 18062 49026 18114 49038
rect 21982 49026 22034 49038
rect 24222 49026 24274 49038
rect 25006 49026 25058 49038
rect 19618 48974 19630 49026
rect 19682 48974 19694 49026
rect 20066 48974 20078 49026
rect 20130 48974 20142 49026
rect 23090 48974 23102 49026
rect 23154 48974 23166 49026
rect 23762 48974 23774 49026
rect 23826 48974 23838 49026
rect 24770 48974 24782 49026
rect 24834 48974 24846 49026
rect 18062 48962 18114 48974
rect 21982 48962 22034 48974
rect 24222 48962 24274 48974
rect 25006 48962 25058 48974
rect 25230 49026 25282 49038
rect 32958 49026 33010 49038
rect 34862 49026 34914 49038
rect 44718 49026 44770 49038
rect 48974 49026 49026 49038
rect 30706 48974 30718 49026
rect 30770 48974 30782 49026
rect 32610 48974 32622 49026
rect 32674 48974 32686 49026
rect 34402 48974 34414 49026
rect 34466 48974 34478 49026
rect 36082 48974 36094 49026
rect 36146 48974 36158 49026
rect 46386 48974 46398 49026
rect 46450 48974 46462 49026
rect 25230 48962 25282 48974
rect 32958 48962 33010 48974
rect 34862 48962 34914 48974
rect 44718 48962 44770 48974
rect 48974 48962 49026 48974
rect 49422 49026 49474 49038
rect 49422 48962 49474 48974
rect 49646 49026 49698 49038
rect 52558 49026 52610 49038
rect 51650 48974 51662 49026
rect 51714 48974 51726 49026
rect 51986 48974 51998 49026
rect 52050 48974 52062 49026
rect 49646 48962 49698 48974
rect 52558 48962 52610 48974
rect 53678 49026 53730 49038
rect 57822 49026 57874 49038
rect 56690 48974 56702 49026
rect 56754 48974 56766 49026
rect 57586 48974 57598 49026
rect 57650 48974 57662 49026
rect 53678 48962 53730 48974
rect 57822 48962 57874 48974
rect 58270 49026 58322 49038
rect 58270 48962 58322 48974
rect 6974 48914 7026 48926
rect 6974 48850 7026 48862
rect 18174 48914 18226 48926
rect 18174 48850 18226 48862
rect 21646 48914 21698 48926
rect 21646 48850 21698 48862
rect 21758 48914 21810 48926
rect 21758 48850 21810 48862
rect 25454 48914 25506 48926
rect 25454 48850 25506 48862
rect 39566 48914 39618 48926
rect 39566 48850 39618 48862
rect 41806 48914 41858 48926
rect 41806 48850 41858 48862
rect 43262 48914 43314 48926
rect 43262 48850 43314 48862
rect 43374 48914 43426 48926
rect 43374 48850 43426 48862
rect 52334 48914 52386 48926
rect 52334 48850 52386 48862
rect 53342 48914 53394 48926
rect 53342 48850 53394 48862
rect 53566 48914 53618 48926
rect 53566 48850 53618 48862
rect 55358 48914 55410 48926
rect 55358 48850 55410 48862
rect 2382 48802 2434 48814
rect 2382 48738 2434 48750
rect 2830 48802 2882 48814
rect 2830 48738 2882 48750
rect 3278 48802 3330 48814
rect 3278 48738 3330 48750
rect 4622 48802 4674 48814
rect 4622 48738 4674 48750
rect 5854 48802 5906 48814
rect 5854 48738 5906 48750
rect 5966 48802 6018 48814
rect 5966 48738 6018 48750
rect 7198 48802 7250 48814
rect 7198 48738 7250 48750
rect 7422 48802 7474 48814
rect 7422 48738 7474 48750
rect 7870 48802 7922 48814
rect 7870 48738 7922 48750
rect 8430 48802 8482 48814
rect 8430 48738 8482 48750
rect 8878 48802 8930 48814
rect 8878 48738 8930 48750
rect 10110 48802 10162 48814
rect 10110 48738 10162 48750
rect 11006 48802 11058 48814
rect 11006 48738 11058 48750
rect 12574 48802 12626 48814
rect 12574 48738 12626 48750
rect 12686 48802 12738 48814
rect 12686 48738 12738 48750
rect 15038 48802 15090 48814
rect 15038 48738 15090 48750
rect 16046 48802 16098 48814
rect 16046 48738 16098 48750
rect 16494 48802 16546 48814
rect 16494 48738 16546 48750
rect 18398 48802 18450 48814
rect 18398 48738 18450 48750
rect 18510 48802 18562 48814
rect 18510 48738 18562 48750
rect 26014 48802 26066 48814
rect 26014 48738 26066 48750
rect 26798 48802 26850 48814
rect 26798 48738 26850 48750
rect 27582 48802 27634 48814
rect 27582 48738 27634 48750
rect 37550 48802 37602 48814
rect 37550 48738 37602 48750
rect 37886 48802 37938 48814
rect 37886 48738 37938 48750
rect 39230 48802 39282 48814
rect 39230 48738 39282 48750
rect 39454 48802 39506 48814
rect 39454 48738 39506 48750
rect 42030 48802 42082 48814
rect 42030 48738 42082 48750
rect 43598 48802 43650 48814
rect 43598 48738 43650 48750
rect 44606 48802 44658 48814
rect 44606 48738 44658 48750
rect 51102 48802 51154 48814
rect 51102 48738 51154 48750
rect 55470 48802 55522 48814
rect 55470 48738 55522 48750
rect 1344 48634 59024 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 59024 48634
rect 1344 48548 59024 48582
rect 2046 48466 2098 48478
rect 2046 48402 2098 48414
rect 2830 48466 2882 48478
rect 2830 48402 2882 48414
rect 3390 48466 3442 48478
rect 9774 48466 9826 48478
rect 8754 48414 8766 48466
rect 8818 48414 8830 48466
rect 3390 48402 3442 48414
rect 9774 48402 9826 48414
rect 11790 48466 11842 48478
rect 11790 48402 11842 48414
rect 12238 48466 12290 48478
rect 12238 48402 12290 48414
rect 14590 48466 14642 48478
rect 14590 48402 14642 48414
rect 15710 48466 15762 48478
rect 15710 48402 15762 48414
rect 16942 48466 16994 48478
rect 16942 48402 16994 48414
rect 19294 48466 19346 48478
rect 22654 48466 22706 48478
rect 21074 48414 21086 48466
rect 21138 48414 21150 48466
rect 19294 48402 19346 48414
rect 22654 48402 22706 48414
rect 23438 48466 23490 48478
rect 23438 48402 23490 48414
rect 25790 48466 25842 48478
rect 25790 48402 25842 48414
rect 49534 48466 49586 48478
rect 49534 48402 49586 48414
rect 52558 48466 52610 48478
rect 52558 48402 52610 48414
rect 53118 48466 53170 48478
rect 53118 48402 53170 48414
rect 15486 48354 15538 48366
rect 5394 48302 5406 48354
rect 5458 48302 5470 48354
rect 15486 48290 15538 48302
rect 16158 48354 16210 48366
rect 23326 48354 23378 48366
rect 20850 48302 20862 48354
rect 20914 48302 20926 48354
rect 21522 48302 21534 48354
rect 21586 48302 21598 48354
rect 16158 48290 16210 48302
rect 23326 48290 23378 48302
rect 26574 48354 26626 48366
rect 26574 48290 26626 48302
rect 33630 48354 33682 48366
rect 33630 48290 33682 48302
rect 40462 48354 40514 48366
rect 40462 48290 40514 48302
rect 43822 48354 43874 48366
rect 43822 48290 43874 48302
rect 46622 48354 46674 48366
rect 46622 48290 46674 48302
rect 52670 48354 52722 48366
rect 52670 48290 52722 48302
rect 57486 48354 57538 48366
rect 57486 48290 57538 48302
rect 7534 48242 7586 48254
rect 10110 48242 10162 48254
rect 5170 48190 5182 48242
rect 5234 48190 5246 48242
rect 6738 48190 6750 48242
rect 6802 48190 6814 48242
rect 8418 48190 8430 48242
rect 8482 48190 8494 48242
rect 9762 48190 9774 48242
rect 9826 48190 9838 48242
rect 7534 48178 7586 48190
rect 10110 48178 10162 48190
rect 10222 48242 10274 48254
rect 10222 48178 10274 48190
rect 10558 48242 10610 48254
rect 10558 48178 10610 48190
rect 11342 48242 11394 48254
rect 11342 48178 11394 48190
rect 12798 48242 12850 48254
rect 12798 48178 12850 48190
rect 12910 48242 12962 48254
rect 12910 48178 12962 48190
rect 13134 48242 13186 48254
rect 13134 48178 13186 48190
rect 13358 48242 13410 48254
rect 14366 48242 14418 48254
rect 15934 48242 15986 48254
rect 23550 48242 23602 48254
rect 14130 48190 14142 48242
rect 14194 48190 14206 48242
rect 14802 48190 14814 48242
rect 14866 48190 14878 48242
rect 17938 48190 17950 48242
rect 18002 48190 18014 48242
rect 20178 48190 20190 48242
rect 20242 48190 20254 48242
rect 20738 48190 20750 48242
rect 20802 48190 20814 48242
rect 21746 48190 21758 48242
rect 21810 48190 21822 48242
rect 13358 48178 13410 48190
rect 14366 48178 14418 48190
rect 15934 48178 15986 48190
rect 23550 48178 23602 48190
rect 23998 48242 24050 48254
rect 30830 48242 30882 48254
rect 36430 48242 36482 48254
rect 28242 48190 28254 48242
rect 28306 48190 28318 48242
rect 30034 48190 30046 48242
rect 30098 48190 30110 48242
rect 31154 48190 31166 48242
rect 31218 48190 31230 48242
rect 33842 48190 33854 48242
rect 33906 48190 33918 48242
rect 34066 48190 34078 48242
rect 34130 48190 34142 48242
rect 35970 48190 35982 48242
rect 36034 48190 36046 48242
rect 23998 48178 24050 48190
rect 30830 48178 30882 48190
rect 36430 48178 36482 48190
rect 37886 48242 37938 48254
rect 46510 48242 46562 48254
rect 38098 48190 38110 48242
rect 38162 48190 38174 48242
rect 39554 48190 39566 48242
rect 39618 48190 39630 48242
rect 43138 48190 43150 48242
rect 43202 48190 43214 48242
rect 46162 48190 46174 48242
rect 46226 48190 46238 48242
rect 37886 48178 37938 48190
rect 46510 48178 46562 48190
rect 51662 48242 51714 48254
rect 52446 48242 52498 48254
rect 51986 48190 51998 48242
rect 52050 48190 52062 48242
rect 51662 48178 51714 48190
rect 52446 48178 52498 48190
rect 54798 48242 54850 48254
rect 57598 48242 57650 48254
rect 55346 48190 55358 48242
rect 55410 48190 55422 48242
rect 57922 48190 57934 48242
rect 57986 48190 57998 48242
rect 54798 48178 54850 48190
rect 57598 48178 57650 48190
rect 2382 48130 2434 48142
rect 2382 48066 2434 48078
rect 3950 48130 4002 48142
rect 3950 48066 4002 48078
rect 14478 48130 14530 48142
rect 14478 48066 14530 48078
rect 16270 48130 16322 48142
rect 23774 48130 23826 48142
rect 17826 48078 17838 48130
rect 17890 48078 17902 48130
rect 16270 48066 16322 48078
rect 23774 48066 23826 48078
rect 24446 48130 24498 48142
rect 24446 48066 24498 48078
rect 24894 48130 24946 48142
rect 36990 48130 37042 48142
rect 28130 48078 28142 48130
rect 28194 48078 28206 48130
rect 29922 48078 29934 48130
rect 29986 48078 29998 48130
rect 35634 48078 35646 48130
rect 35698 48078 35710 48130
rect 24894 48066 24946 48078
rect 36990 48066 37042 48078
rect 38782 48130 38834 48142
rect 49646 48130 49698 48142
rect 39666 48078 39678 48130
rect 39730 48078 39742 48130
rect 43362 48078 43374 48130
rect 43426 48078 43438 48130
rect 38782 48066 38834 48078
rect 49646 48066 49698 48078
rect 50206 48130 50258 48142
rect 50206 48066 50258 48078
rect 50654 48130 50706 48142
rect 50654 48066 50706 48078
rect 51214 48130 51266 48142
rect 56702 48130 56754 48142
rect 55682 48078 55694 48130
rect 55746 48078 55758 48130
rect 51214 48066 51266 48078
rect 56702 48066 56754 48078
rect 50878 48018 50930 48030
rect 18386 47966 18398 48018
rect 18450 47966 18462 48018
rect 27906 47966 27918 48018
rect 27970 47966 27982 48018
rect 50878 47954 50930 47966
rect 52222 48018 52274 48030
rect 52222 47954 52274 47966
rect 1344 47850 59024 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 59024 47850
rect 1344 47764 59024 47798
rect 3838 47682 3890 47694
rect 3838 47618 3890 47630
rect 9326 47682 9378 47694
rect 9326 47618 9378 47630
rect 9774 47682 9826 47694
rect 36206 47682 36258 47694
rect 12002 47630 12014 47682
rect 12066 47679 12078 47682
rect 12898 47679 12910 47682
rect 12066 47633 12910 47679
rect 12066 47630 12078 47633
rect 12898 47630 12910 47633
rect 12962 47630 12974 47682
rect 26114 47630 26126 47682
rect 26178 47679 26190 47682
rect 26562 47679 26574 47682
rect 26178 47633 26574 47679
rect 26178 47630 26190 47633
rect 26562 47630 26574 47633
rect 26626 47679 26638 47682
rect 26786 47679 26798 47682
rect 26626 47633 26798 47679
rect 26626 47630 26638 47633
rect 26786 47630 26798 47633
rect 26850 47630 26862 47682
rect 34514 47630 34526 47682
rect 34578 47630 34590 47682
rect 52210 47630 52222 47682
rect 52274 47630 52286 47682
rect 9774 47618 9826 47630
rect 36206 47618 36258 47630
rect 2830 47570 2882 47582
rect 2830 47506 2882 47518
rect 3502 47570 3554 47582
rect 3502 47506 3554 47518
rect 7310 47570 7362 47582
rect 7310 47506 7362 47518
rect 7534 47570 7586 47582
rect 7534 47506 7586 47518
rect 8654 47570 8706 47582
rect 12014 47570 12066 47582
rect 11442 47518 11454 47570
rect 11506 47518 11518 47570
rect 8654 47506 8706 47518
rect 12014 47506 12066 47518
rect 13022 47570 13074 47582
rect 13022 47506 13074 47518
rect 15150 47570 15202 47582
rect 21982 47570 22034 47582
rect 17602 47518 17614 47570
rect 17666 47518 17678 47570
rect 18050 47518 18062 47570
rect 18114 47518 18126 47570
rect 20066 47518 20078 47570
rect 20130 47518 20142 47570
rect 15150 47506 15202 47518
rect 21982 47506 22034 47518
rect 22878 47570 22930 47582
rect 22878 47506 22930 47518
rect 26126 47570 26178 47582
rect 26126 47506 26178 47518
rect 26574 47570 26626 47582
rect 26574 47506 26626 47518
rect 27246 47570 27298 47582
rect 27246 47506 27298 47518
rect 28366 47570 28418 47582
rect 28366 47506 28418 47518
rect 28814 47570 28866 47582
rect 38558 47570 38610 47582
rect 31266 47518 31278 47570
rect 31330 47518 31342 47570
rect 32946 47518 32958 47570
rect 33010 47518 33022 47570
rect 28814 47506 28866 47518
rect 38558 47506 38610 47518
rect 40798 47570 40850 47582
rect 40798 47506 40850 47518
rect 42478 47570 42530 47582
rect 42478 47506 42530 47518
rect 45614 47570 45666 47582
rect 45614 47506 45666 47518
rect 46734 47570 46786 47582
rect 56366 47570 56418 47582
rect 55346 47518 55358 47570
rect 55410 47518 55422 47570
rect 46734 47506 46786 47518
rect 56366 47506 56418 47518
rect 2606 47458 2658 47470
rect 6078 47458 6130 47470
rect 7646 47458 7698 47470
rect 4162 47406 4174 47458
rect 4226 47406 4238 47458
rect 7074 47406 7086 47458
rect 7138 47406 7150 47458
rect 2606 47394 2658 47406
rect 6078 47394 6130 47406
rect 7646 47394 7698 47406
rect 9438 47458 9490 47470
rect 9438 47394 9490 47406
rect 9998 47458 10050 47470
rect 9998 47394 10050 47406
rect 10670 47458 10722 47470
rect 10670 47394 10722 47406
rect 15710 47458 15762 47470
rect 15710 47394 15762 47406
rect 15934 47458 15986 47470
rect 19854 47458 19906 47470
rect 23326 47458 23378 47470
rect 16258 47406 16270 47458
rect 16322 47406 16334 47458
rect 17266 47406 17278 47458
rect 17330 47406 17342 47458
rect 18162 47406 18174 47458
rect 18226 47406 18238 47458
rect 20626 47406 20638 47458
rect 20690 47406 20702 47458
rect 15934 47394 15986 47406
rect 19854 47394 19906 47406
rect 23326 47394 23378 47406
rect 27134 47458 27186 47470
rect 27134 47394 27186 47406
rect 27358 47458 27410 47470
rect 37438 47458 37490 47470
rect 31714 47406 31726 47458
rect 31778 47406 31790 47458
rect 33170 47406 33182 47458
rect 33234 47406 33246 47458
rect 34066 47406 34078 47458
rect 34130 47406 34142 47458
rect 34514 47406 34526 47458
rect 34578 47406 34590 47458
rect 36194 47406 36206 47458
rect 36258 47406 36270 47458
rect 27358 47394 27410 47406
rect 37438 47394 37490 47406
rect 38446 47458 38498 47470
rect 38446 47394 38498 47406
rect 39118 47458 39170 47470
rect 39118 47394 39170 47406
rect 41022 47458 41074 47470
rect 41022 47394 41074 47406
rect 41582 47458 41634 47470
rect 44606 47458 44658 47470
rect 41794 47406 41806 47458
rect 41858 47406 41870 47458
rect 44034 47406 44046 47458
rect 44098 47406 44110 47458
rect 41582 47394 41634 47406
rect 44606 47394 44658 47406
rect 45390 47458 45442 47470
rect 45390 47394 45442 47406
rect 46062 47458 46114 47470
rect 46062 47394 46114 47406
rect 51662 47458 51714 47470
rect 51662 47394 51714 47406
rect 51886 47458 51938 47470
rect 51886 47394 51938 47406
rect 54574 47458 54626 47470
rect 56814 47458 56866 47470
rect 55234 47406 55246 47458
rect 55298 47406 55310 47458
rect 54574 47394 54626 47406
rect 56814 47394 56866 47406
rect 3390 47346 3442 47358
rect 9214 47346 9266 47358
rect 3602 47294 3614 47346
rect 3666 47294 3678 47346
rect 3390 47282 3442 47294
rect 9214 47282 9266 47294
rect 10894 47346 10946 47358
rect 10894 47282 10946 47294
rect 11006 47346 11058 47358
rect 19294 47346 19346 47358
rect 11106 47294 11118 47346
rect 11170 47294 11182 47346
rect 18498 47294 18510 47346
rect 18562 47294 18574 47346
rect 11006 47282 11058 47294
rect 19294 47282 19346 47294
rect 20190 47346 20242 47358
rect 20190 47282 20242 47294
rect 24558 47346 24610 47358
rect 24558 47282 24610 47294
rect 27582 47346 27634 47358
rect 27582 47282 27634 47294
rect 36542 47346 36594 47358
rect 36542 47282 36594 47294
rect 39454 47346 39506 47358
rect 39454 47282 39506 47294
rect 40350 47346 40402 47358
rect 40350 47282 40402 47294
rect 40574 47346 40626 47358
rect 40574 47282 40626 47294
rect 44718 47346 44770 47358
rect 44718 47282 44770 47294
rect 45838 47346 45890 47358
rect 45838 47282 45890 47294
rect 46622 47346 46674 47358
rect 46622 47282 46674 47294
rect 46846 47346 46898 47358
rect 46846 47282 46898 47294
rect 48190 47346 48242 47358
rect 48190 47282 48242 47294
rect 56254 47346 56306 47358
rect 56254 47282 56306 47294
rect 56590 47346 56642 47358
rect 56590 47282 56642 47294
rect 1822 47234 1874 47246
rect 4958 47234 5010 47246
rect 2258 47182 2270 47234
rect 2322 47182 2334 47234
rect 1822 47170 1874 47182
rect 4958 47170 5010 47182
rect 12462 47234 12514 47246
rect 12462 47170 12514 47182
rect 13694 47234 13746 47246
rect 13694 47170 13746 47182
rect 14478 47234 14530 47246
rect 14478 47170 14530 47182
rect 15822 47234 15874 47246
rect 15822 47170 15874 47182
rect 20078 47234 20130 47246
rect 20078 47170 20130 47182
rect 21646 47234 21698 47246
rect 21646 47170 21698 47182
rect 22430 47234 22482 47246
rect 22430 47170 22482 47182
rect 23774 47234 23826 47246
rect 23774 47170 23826 47182
rect 24334 47234 24386 47246
rect 24334 47170 24386 47182
rect 24446 47234 24498 47246
rect 24446 47170 24498 47182
rect 24782 47234 24834 47246
rect 24782 47170 24834 47182
rect 25678 47234 25730 47246
rect 25678 47170 25730 47182
rect 29710 47234 29762 47246
rect 29710 47170 29762 47182
rect 37998 47234 38050 47246
rect 37998 47170 38050 47182
rect 38670 47234 38722 47246
rect 38670 47170 38722 47182
rect 48302 47234 48354 47246
rect 48302 47170 48354 47182
rect 48526 47234 48578 47246
rect 48526 47170 48578 47182
rect 48862 47234 48914 47246
rect 48862 47170 48914 47182
rect 51102 47234 51154 47246
rect 51102 47170 51154 47182
rect 1344 47066 59024 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 59024 47066
rect 1344 46980 59024 47014
rect 2382 46898 2434 46910
rect 2382 46834 2434 46846
rect 3166 46898 3218 46910
rect 3166 46834 3218 46846
rect 4846 46898 4898 46910
rect 4846 46834 4898 46846
rect 6078 46898 6130 46910
rect 6078 46834 6130 46846
rect 6862 46898 6914 46910
rect 6862 46834 6914 46846
rect 8766 46898 8818 46910
rect 8766 46834 8818 46846
rect 10670 46898 10722 46910
rect 10670 46834 10722 46846
rect 11454 46898 11506 46910
rect 11454 46834 11506 46846
rect 12910 46898 12962 46910
rect 12910 46834 12962 46846
rect 14142 46898 14194 46910
rect 22990 46898 23042 46910
rect 16930 46846 16942 46898
rect 16994 46846 17006 46898
rect 14142 46834 14194 46846
rect 22990 46834 23042 46846
rect 32622 46898 32674 46910
rect 36654 46898 36706 46910
rect 33618 46846 33630 46898
rect 33682 46846 33694 46898
rect 32622 46834 32674 46846
rect 36654 46834 36706 46846
rect 38110 46898 38162 46910
rect 38110 46834 38162 46846
rect 38446 46898 38498 46910
rect 38446 46834 38498 46846
rect 45614 46898 45666 46910
rect 45614 46834 45666 46846
rect 49646 46898 49698 46910
rect 49646 46834 49698 46846
rect 49982 46898 50034 46910
rect 49982 46834 50034 46846
rect 3390 46786 3442 46798
rect 3390 46722 3442 46734
rect 3502 46786 3554 46798
rect 3502 46722 3554 46734
rect 4734 46786 4786 46798
rect 4734 46722 4786 46734
rect 4958 46786 5010 46798
rect 4958 46722 5010 46734
rect 6638 46786 6690 46798
rect 6638 46722 6690 46734
rect 7646 46786 7698 46798
rect 7646 46722 7698 46734
rect 8990 46786 9042 46798
rect 8990 46722 9042 46734
rect 10334 46786 10386 46798
rect 10334 46722 10386 46734
rect 10558 46786 10610 46798
rect 10558 46722 10610 46734
rect 14254 46786 14306 46798
rect 23774 46786 23826 46798
rect 14354 46734 14366 46786
rect 14418 46734 14430 46786
rect 18498 46734 18510 46786
rect 18562 46734 18574 46786
rect 21186 46734 21198 46786
rect 21250 46734 21262 46786
rect 14254 46722 14306 46734
rect 23774 46722 23826 46734
rect 36206 46786 36258 46798
rect 36206 46722 36258 46734
rect 36878 46786 36930 46798
rect 36878 46722 36930 46734
rect 37886 46786 37938 46798
rect 37886 46722 37938 46734
rect 40014 46786 40066 46798
rect 40014 46722 40066 46734
rect 45502 46786 45554 46798
rect 45502 46722 45554 46734
rect 53230 46786 53282 46798
rect 53230 46722 53282 46734
rect 55694 46786 55746 46798
rect 55694 46722 55746 46734
rect 57486 46786 57538 46798
rect 57486 46722 57538 46734
rect 2830 46674 2882 46686
rect 2830 46610 2882 46622
rect 6974 46674 7026 46686
rect 6974 46610 7026 46622
rect 7198 46674 7250 46686
rect 7198 46610 7250 46622
rect 10782 46674 10834 46686
rect 10782 46610 10834 46622
rect 11790 46674 11842 46686
rect 11790 46610 11842 46622
rect 12350 46674 12402 46686
rect 12350 46610 12402 46622
rect 12798 46674 12850 46686
rect 12798 46610 12850 46622
rect 13022 46674 13074 46686
rect 13022 46610 13074 46622
rect 13918 46674 13970 46686
rect 13918 46610 13970 46622
rect 15262 46674 15314 46686
rect 15262 46610 15314 46622
rect 16606 46674 16658 46686
rect 23998 46674 24050 46686
rect 26238 46674 26290 46686
rect 30158 46674 30210 46686
rect 34190 46674 34242 46686
rect 36990 46674 37042 46686
rect 17826 46622 17838 46674
rect 17890 46622 17902 46674
rect 19842 46622 19854 46674
rect 19906 46622 19918 46674
rect 21298 46622 21310 46674
rect 21362 46622 21374 46674
rect 23538 46622 23550 46674
rect 23602 46622 23614 46674
rect 24210 46622 24222 46674
rect 24274 46622 24286 46674
rect 28242 46622 28254 46674
rect 28306 46622 28318 46674
rect 29922 46622 29934 46674
rect 29986 46622 29998 46674
rect 30594 46622 30606 46674
rect 30658 46622 30670 46674
rect 30818 46622 30830 46674
rect 30882 46622 30894 46674
rect 35746 46622 35758 46674
rect 35810 46622 35822 46674
rect 16606 46610 16658 46622
rect 23998 46610 24050 46622
rect 26238 46610 26290 46622
rect 30158 46610 30210 46622
rect 34190 46610 34242 46622
rect 36990 46610 37042 46622
rect 37774 46674 37826 46686
rect 48750 46674 48802 46686
rect 39554 46622 39566 46674
rect 39618 46622 39630 46674
rect 47842 46622 47854 46674
rect 47906 46622 47918 46674
rect 37774 46610 37826 46622
rect 48750 46610 48802 46622
rect 49534 46674 49586 46686
rect 49534 46610 49586 46622
rect 49758 46674 49810 46686
rect 49758 46610 49810 46622
rect 55246 46674 55298 46686
rect 55246 46610 55298 46622
rect 55470 46674 55522 46686
rect 55470 46610 55522 46622
rect 55918 46674 55970 46686
rect 58146 46622 58158 46674
rect 58210 46622 58222 46674
rect 55918 46610 55970 46622
rect 1934 46562 1986 46574
rect 1934 46498 1986 46510
rect 4174 46562 4226 46574
rect 4174 46498 4226 46510
rect 5630 46562 5682 46574
rect 5630 46498 5682 46510
rect 8094 46562 8146 46574
rect 8094 46498 8146 46510
rect 8878 46562 8930 46574
rect 8878 46498 8930 46510
rect 9774 46562 9826 46574
rect 15822 46562 15874 46574
rect 14690 46510 14702 46562
rect 14754 46510 14766 46562
rect 9774 46498 9826 46510
rect 15822 46498 15874 46510
rect 16382 46562 16434 46574
rect 16382 46498 16434 46510
rect 20414 46562 20466 46574
rect 20414 46498 20466 46510
rect 22542 46562 22594 46574
rect 22542 46498 22594 46510
rect 23886 46562 23938 46574
rect 23886 46498 23938 46510
rect 25006 46562 25058 46574
rect 42590 46562 42642 46574
rect 27794 46510 27806 46562
rect 27858 46510 27870 46562
rect 35858 46510 35870 46562
rect 35922 46510 35934 46562
rect 39218 46510 39230 46562
rect 39282 46510 39294 46562
rect 25006 46498 25058 46510
rect 42590 46498 42642 46510
rect 47070 46562 47122 46574
rect 54014 46562 54066 46574
rect 47954 46510 47966 46562
rect 48018 46510 48030 46562
rect 53106 46510 53118 46562
rect 53170 46510 53182 46562
rect 47070 46498 47122 46510
rect 54014 46498 54066 46510
rect 56478 46562 56530 46574
rect 57810 46510 57822 46562
rect 57874 46510 57886 46562
rect 56478 46498 56530 46510
rect 11454 46450 11506 46462
rect 11454 46386 11506 46398
rect 11566 46450 11618 46462
rect 26014 46450 26066 46462
rect 33966 46450 34018 46462
rect 25666 46398 25678 46450
rect 25730 46398 25742 46450
rect 29362 46398 29374 46450
rect 29426 46398 29438 46450
rect 11566 46386 11618 46398
rect 26014 46386 26066 46398
rect 33966 46386 34018 46398
rect 53454 46450 53506 46462
rect 53454 46386 53506 46398
rect 56030 46450 56082 46462
rect 56030 46386 56082 46398
rect 1344 46282 59024 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 59024 46282
rect 1344 46196 59024 46230
rect 3614 46114 3666 46126
rect 39342 46114 39394 46126
rect 30930 46062 30942 46114
rect 30994 46111 31006 46114
rect 31714 46111 31726 46114
rect 30994 46065 31726 46111
rect 30994 46062 31006 46065
rect 31714 46062 31726 46065
rect 31778 46062 31790 46114
rect 38546 46062 38558 46114
rect 38610 46062 38622 46114
rect 3614 46050 3666 46062
rect 39342 46050 39394 46062
rect 39678 46114 39730 46126
rect 39678 46050 39730 46062
rect 43150 46114 43202 46126
rect 43150 46050 43202 46062
rect 46734 46114 46786 46126
rect 46734 46050 46786 46062
rect 55582 46114 55634 46126
rect 57822 46114 57874 46126
rect 57474 46062 57486 46114
rect 57538 46062 57550 46114
rect 55582 46050 55634 46062
rect 57822 46050 57874 46062
rect 1934 46002 1986 46014
rect 1934 45938 1986 45950
rect 6750 46002 6802 46014
rect 6750 45938 6802 45950
rect 9774 46002 9826 46014
rect 9774 45938 9826 45950
rect 12126 46002 12178 46014
rect 12126 45938 12178 45950
rect 12686 46002 12738 46014
rect 22878 46002 22930 46014
rect 15250 45950 15262 46002
rect 15314 45950 15326 46002
rect 12686 45938 12738 45950
rect 22878 45938 22930 45950
rect 26910 46002 26962 46014
rect 31166 46002 31218 46014
rect 29586 45950 29598 46002
rect 29650 45950 29662 46002
rect 26910 45938 26962 45950
rect 31166 45938 31218 45950
rect 31614 46002 31666 46014
rect 31614 45938 31666 45950
rect 33406 46002 33458 46014
rect 33406 45938 33458 45950
rect 34190 46002 34242 46014
rect 34190 45938 34242 45950
rect 35646 46002 35698 46014
rect 41246 46002 41298 46014
rect 37986 45950 37998 46002
rect 38050 45950 38062 46002
rect 35646 45938 35698 45950
rect 41246 45938 41298 45950
rect 44718 46002 44770 46014
rect 44718 45938 44770 45950
rect 45614 46002 45666 46014
rect 54462 46002 54514 46014
rect 48738 45950 48750 46002
rect 48802 45950 48814 46002
rect 45614 45938 45666 45950
rect 54462 45938 54514 45950
rect 56142 46002 56194 46014
rect 56142 45938 56194 45950
rect 56590 46002 56642 46014
rect 56590 45938 56642 45950
rect 3278 45890 3330 45902
rect 2818 45838 2830 45890
rect 2882 45838 2894 45890
rect 3278 45826 3330 45838
rect 6526 45890 6578 45902
rect 6526 45826 6578 45838
rect 6638 45890 6690 45902
rect 6638 45826 6690 45838
rect 7534 45890 7586 45902
rect 7534 45826 7586 45838
rect 7982 45890 8034 45902
rect 7982 45826 8034 45838
rect 8766 45890 8818 45902
rect 8766 45826 8818 45838
rect 9102 45890 9154 45902
rect 18174 45890 18226 45902
rect 22654 45890 22706 45902
rect 10322 45838 10334 45890
rect 10386 45838 10398 45890
rect 14690 45838 14702 45890
rect 14754 45838 14766 45890
rect 15362 45838 15374 45890
rect 15426 45838 15438 45890
rect 17378 45838 17390 45890
rect 17442 45838 17454 45890
rect 18498 45838 18510 45890
rect 18562 45838 18574 45890
rect 20514 45838 20526 45890
rect 20578 45838 20590 45890
rect 9102 45826 9154 45838
rect 18174 45826 18226 45838
rect 22654 45826 22706 45838
rect 23326 45890 23378 45902
rect 25454 45890 25506 45902
rect 24322 45838 24334 45890
rect 24386 45838 24398 45890
rect 23326 45826 23378 45838
rect 25454 45826 25506 45838
rect 30718 45890 30770 45902
rect 30718 45826 30770 45838
rect 33518 45890 33570 45902
rect 33518 45826 33570 45838
rect 34302 45890 34354 45902
rect 34302 45826 34354 45838
rect 34750 45890 34802 45902
rect 34750 45826 34802 45838
rect 36206 45890 36258 45902
rect 42142 45890 42194 45902
rect 37762 45838 37774 45890
rect 37826 45838 37838 45890
rect 41682 45838 41694 45890
rect 41746 45838 41758 45890
rect 36206 45826 36258 45838
rect 42142 45826 42194 45838
rect 42814 45890 42866 45902
rect 42814 45826 42866 45838
rect 45726 45890 45778 45902
rect 45726 45826 45778 45838
rect 45950 45890 46002 45902
rect 51326 45890 51378 45902
rect 48962 45838 48974 45890
rect 49026 45838 49038 45890
rect 45950 45826 46002 45838
rect 51326 45826 51378 45838
rect 51550 45890 51602 45902
rect 55918 45890 55970 45902
rect 53778 45838 53790 45890
rect 53842 45838 53854 45890
rect 54226 45838 54238 45890
rect 54290 45838 54302 45890
rect 51550 45826 51602 45838
rect 55918 45826 55970 45838
rect 58046 45890 58098 45902
rect 58046 45826 58098 45838
rect 4398 45778 4450 45790
rect 2482 45726 2494 45778
rect 2546 45726 2558 45778
rect 4398 45714 4450 45726
rect 4510 45778 4562 45790
rect 4510 45714 4562 45726
rect 7086 45778 7138 45790
rect 7086 45714 7138 45726
rect 8206 45778 8258 45790
rect 8206 45714 8258 45726
rect 10894 45778 10946 45790
rect 10894 45714 10946 45726
rect 13918 45778 13970 45790
rect 13918 45714 13970 45726
rect 14030 45778 14082 45790
rect 24782 45778 24834 45790
rect 16034 45726 16046 45778
rect 16098 45726 16110 45778
rect 20178 45726 20190 45778
rect 20242 45726 20254 45778
rect 24210 45726 24222 45778
rect 24274 45726 24286 45778
rect 14030 45714 14082 45726
rect 24782 45714 24834 45726
rect 25566 45778 25618 45790
rect 25566 45714 25618 45726
rect 25790 45778 25842 45790
rect 25790 45714 25842 45726
rect 26798 45778 26850 45790
rect 26798 45714 26850 45726
rect 27134 45778 27186 45790
rect 27134 45714 27186 45726
rect 27358 45778 27410 45790
rect 27358 45714 27410 45726
rect 29710 45778 29762 45790
rect 29710 45714 29762 45726
rect 29934 45778 29986 45790
rect 29934 45714 29986 45726
rect 30606 45778 30658 45790
rect 30606 45714 30658 45726
rect 33070 45778 33122 45790
rect 33070 45714 33122 45726
rect 34078 45778 34130 45790
rect 34078 45714 34130 45726
rect 35758 45778 35810 45790
rect 35758 45714 35810 45726
rect 40238 45778 40290 45790
rect 40238 45714 40290 45726
rect 43038 45778 43090 45790
rect 43038 45714 43090 45726
rect 45502 45778 45554 45790
rect 45502 45714 45554 45726
rect 46622 45778 46674 45790
rect 46622 45714 46674 45726
rect 49646 45778 49698 45790
rect 49646 45714 49698 45726
rect 4734 45666 4786 45678
rect 4734 45602 4786 45614
rect 5854 45666 5906 45678
rect 5854 45602 5906 45614
rect 6862 45666 6914 45678
rect 6862 45602 6914 45614
rect 7758 45666 7810 45678
rect 7758 45602 7810 45614
rect 8878 45666 8930 45678
rect 8878 45602 8930 45614
rect 14254 45666 14306 45678
rect 21534 45666 21586 45678
rect 19842 45614 19854 45666
rect 19906 45614 19918 45666
rect 14254 45602 14306 45614
rect 21534 45602 21586 45614
rect 22094 45666 22146 45678
rect 22094 45602 22146 45614
rect 23102 45666 23154 45678
rect 23102 45602 23154 45614
rect 23214 45666 23266 45678
rect 23214 45602 23266 45614
rect 24558 45666 24610 45678
rect 24558 45602 24610 45614
rect 24670 45666 24722 45678
rect 24670 45602 24722 45614
rect 25342 45666 25394 45678
rect 25342 45602 25394 45614
rect 28030 45666 28082 45678
rect 28030 45602 28082 45614
rect 28366 45666 28418 45678
rect 28366 45602 28418 45614
rect 28926 45666 28978 45678
rect 28926 45602 28978 45614
rect 30382 45666 30434 45678
rect 30382 45602 30434 45614
rect 32174 45666 32226 45678
rect 32174 45602 32226 45614
rect 33294 45666 33346 45678
rect 33294 45602 33346 45614
rect 35534 45666 35586 45678
rect 35534 45602 35586 45614
rect 36654 45666 36706 45678
rect 36654 45602 36706 45614
rect 39566 45666 39618 45678
rect 39566 45602 39618 45614
rect 40574 45666 40626 45678
rect 40574 45602 40626 45614
rect 44158 45666 44210 45678
rect 44158 45602 44210 45614
rect 46734 45666 46786 45678
rect 54910 45666 54962 45678
rect 51874 45614 51886 45666
rect 51938 45614 51950 45666
rect 46734 45602 46786 45614
rect 54910 45602 54962 45614
rect 1344 45498 59024 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 59024 45498
rect 1344 45412 59024 45446
rect 3054 45330 3106 45342
rect 3054 45266 3106 45278
rect 4398 45330 4450 45342
rect 4398 45266 4450 45278
rect 5182 45330 5234 45342
rect 5182 45266 5234 45278
rect 5406 45330 5458 45342
rect 15598 45330 15650 45342
rect 7186 45278 7198 45330
rect 7250 45278 7262 45330
rect 10770 45278 10782 45330
rect 10834 45278 10846 45330
rect 5406 45266 5458 45278
rect 15598 45266 15650 45278
rect 16942 45330 16994 45342
rect 23998 45330 24050 45342
rect 18274 45278 18286 45330
rect 18338 45278 18350 45330
rect 16942 45266 16994 45278
rect 23998 45266 24050 45278
rect 24110 45330 24162 45342
rect 24110 45266 24162 45278
rect 25006 45330 25058 45342
rect 25006 45266 25058 45278
rect 29486 45330 29538 45342
rect 29486 45266 29538 45278
rect 30270 45330 30322 45342
rect 30270 45266 30322 45278
rect 30494 45330 30546 45342
rect 30494 45266 30546 45278
rect 30606 45330 30658 45342
rect 30606 45266 30658 45278
rect 31726 45330 31778 45342
rect 31726 45266 31778 45278
rect 34638 45330 34690 45342
rect 34638 45266 34690 45278
rect 34750 45330 34802 45342
rect 34750 45266 34802 45278
rect 37102 45330 37154 45342
rect 37102 45266 37154 45278
rect 38446 45330 38498 45342
rect 38446 45266 38498 45278
rect 38782 45330 38834 45342
rect 38782 45266 38834 45278
rect 41470 45330 41522 45342
rect 41470 45266 41522 45278
rect 42814 45330 42866 45342
rect 42814 45266 42866 45278
rect 44494 45330 44546 45342
rect 44494 45266 44546 45278
rect 45054 45330 45106 45342
rect 45054 45266 45106 45278
rect 45166 45330 45218 45342
rect 45166 45266 45218 45278
rect 53566 45330 53618 45342
rect 53566 45266 53618 45278
rect 57934 45330 57986 45342
rect 57934 45266 57986 45278
rect 2158 45218 2210 45230
rect 2158 45154 2210 45166
rect 4174 45218 4226 45230
rect 27246 45218 27298 45230
rect 29374 45218 29426 45230
rect 11330 45166 11342 45218
rect 11394 45166 11406 45218
rect 12786 45166 12798 45218
rect 12850 45166 12862 45218
rect 14802 45166 14814 45218
rect 14866 45166 14878 45218
rect 17826 45166 17838 45218
rect 17890 45166 17902 45218
rect 20962 45166 20974 45218
rect 21026 45166 21038 45218
rect 21634 45166 21646 45218
rect 21698 45166 21710 45218
rect 27570 45166 27582 45218
rect 27634 45166 27646 45218
rect 4174 45154 4226 45166
rect 27246 45154 27298 45166
rect 29374 45154 29426 45166
rect 30830 45218 30882 45230
rect 30830 45154 30882 45166
rect 31614 45218 31666 45230
rect 31614 45154 31666 45166
rect 36654 45218 36706 45230
rect 36654 45154 36706 45166
rect 38222 45218 38274 45230
rect 38222 45154 38274 45166
rect 39790 45218 39842 45230
rect 39790 45154 39842 45166
rect 43598 45218 43650 45230
rect 43598 45154 43650 45166
rect 44158 45218 44210 45230
rect 44158 45154 44210 45166
rect 44270 45218 44322 45230
rect 44270 45154 44322 45166
rect 47518 45218 47570 45230
rect 47518 45154 47570 45166
rect 52894 45218 52946 45230
rect 52894 45154 52946 45166
rect 54014 45218 54066 45230
rect 54014 45154 54066 45166
rect 56366 45218 56418 45230
rect 56366 45154 56418 45166
rect 57598 45218 57650 45230
rect 57598 45154 57650 45166
rect 5070 45106 5122 45118
rect 2482 45054 2494 45106
rect 2546 45054 2558 45106
rect 5070 45042 5122 45054
rect 6638 45106 6690 45118
rect 6638 45042 6690 45054
rect 6862 45106 6914 45118
rect 6862 45042 6914 45054
rect 7198 45106 7250 45118
rect 7198 45042 7250 45054
rect 7646 45106 7698 45118
rect 7646 45042 7698 45054
rect 8094 45106 8146 45118
rect 24222 45106 24274 45118
rect 10770 45054 10782 45106
rect 10834 45054 10846 45106
rect 11666 45054 11678 45106
rect 11730 45054 11742 45106
rect 12562 45054 12574 45106
rect 12626 45054 12638 45106
rect 14466 45054 14478 45106
rect 14530 45054 14542 45106
rect 18050 45054 18062 45106
rect 18114 45054 18126 45106
rect 20178 45054 20190 45106
rect 20242 45054 20254 45106
rect 20850 45054 20862 45106
rect 20914 45054 20926 45106
rect 21746 45054 21758 45106
rect 21810 45054 21822 45106
rect 23762 45054 23774 45106
rect 23826 45054 23838 45106
rect 8094 45042 8146 45054
rect 24222 45042 24274 45054
rect 24334 45106 24386 45118
rect 26910 45106 26962 45118
rect 25666 45054 25678 45106
rect 25730 45054 25742 45106
rect 24334 45042 24386 45054
rect 26910 45042 26962 45054
rect 27694 45106 27746 45118
rect 27694 45042 27746 45054
rect 27806 45106 27858 45118
rect 27806 45042 27858 45054
rect 28590 45106 28642 45118
rect 28590 45042 28642 45054
rect 28814 45106 28866 45118
rect 28814 45042 28866 45054
rect 29262 45106 29314 45118
rect 29262 45042 29314 45054
rect 30382 45106 30434 45118
rect 30382 45042 30434 45054
rect 31390 45106 31442 45118
rect 31390 45042 31442 45054
rect 32062 45106 32114 45118
rect 32062 45042 32114 45054
rect 34526 45106 34578 45118
rect 34526 45042 34578 45054
rect 34862 45106 34914 45118
rect 35758 45106 35810 45118
rect 38110 45106 38162 45118
rect 35074 45054 35086 45106
rect 35138 45054 35150 45106
rect 35970 45054 35982 45106
rect 36034 45054 36046 45106
rect 34862 45042 34914 45054
rect 35758 45042 35810 45054
rect 38110 45042 38162 45054
rect 39678 45106 39730 45118
rect 39678 45042 39730 45054
rect 40014 45106 40066 45118
rect 40014 45042 40066 45054
rect 42254 45106 42306 45118
rect 42254 45042 42306 45054
rect 42702 45106 42754 45118
rect 42702 45042 42754 45054
rect 42926 45106 42978 45118
rect 48750 45106 48802 45118
rect 53342 45106 53394 45118
rect 47058 45054 47070 45106
rect 47122 45054 47134 45106
rect 49858 45054 49870 45106
rect 49922 45054 49934 45106
rect 51986 45054 51998 45106
rect 52050 45054 52062 45106
rect 42926 45042 42978 45054
rect 48750 45042 48802 45054
rect 53342 45042 53394 45054
rect 53790 45106 53842 45118
rect 53790 45042 53842 45054
rect 57822 45106 57874 45118
rect 57822 45042 57874 45054
rect 58046 45106 58098 45118
rect 58046 45042 58098 45054
rect 58494 45106 58546 45118
rect 58494 45042 58546 45054
rect 3614 44994 3666 45006
rect 6078 44994 6130 45006
rect 2370 44942 2382 44994
rect 2434 44942 2446 44994
rect 4498 44942 4510 44994
rect 4562 44942 4574 44994
rect 3614 44930 3666 44942
rect 6078 44930 6130 44942
rect 8654 44994 8706 45006
rect 8654 44930 8706 44942
rect 9662 44994 9714 45006
rect 9662 44930 9714 44942
rect 10222 44994 10274 45006
rect 10222 44930 10274 44942
rect 16158 44994 16210 45006
rect 16158 44930 16210 44942
rect 16494 44994 16546 45006
rect 16494 44930 16546 44942
rect 18846 44994 18898 45006
rect 18846 44930 18898 44942
rect 19294 44994 19346 45006
rect 22766 44994 22818 45006
rect 21522 44942 21534 44994
rect 21586 44942 21598 44994
rect 19294 44930 19346 44942
rect 22766 44930 22818 44942
rect 23214 44994 23266 45006
rect 23214 44930 23266 44942
rect 29038 44994 29090 45006
rect 29038 44930 29090 44942
rect 32510 44994 32562 45006
rect 32510 44930 32562 44942
rect 32958 44994 33010 45006
rect 32958 44930 33010 44942
rect 33630 44994 33682 45006
rect 33630 44930 33682 44942
rect 37550 44994 37602 45006
rect 37550 44930 37602 44942
rect 40350 44994 40402 45006
rect 40350 44930 40402 44942
rect 45726 44994 45778 45006
rect 48526 44994 48578 45006
rect 50542 44994 50594 45006
rect 46610 44942 46622 44994
rect 46674 44942 46686 44994
rect 49634 44942 49646 44994
rect 49698 44942 49710 44994
rect 52098 44942 52110 44994
rect 52162 44942 52174 44994
rect 56242 44942 56254 44994
rect 56306 44942 56318 44994
rect 45726 44930 45778 44942
rect 48526 44930 48578 44942
rect 50542 44930 50594 44942
rect 7086 44882 7138 44894
rect 7086 44818 7138 44830
rect 25678 44882 25730 44894
rect 25678 44818 25730 44830
rect 26014 44882 26066 44894
rect 26014 44818 26066 44830
rect 27022 44882 27074 44894
rect 27022 44818 27074 44830
rect 45278 44882 45330 44894
rect 56590 44882 56642 44894
rect 48178 44830 48190 44882
rect 48242 44830 48254 44882
rect 45278 44818 45330 44830
rect 56590 44818 56642 44830
rect 1344 44714 59024 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 59024 44714
rect 1344 44628 59024 44662
rect 6190 44546 6242 44558
rect 6190 44482 6242 44494
rect 6862 44546 6914 44558
rect 6862 44482 6914 44494
rect 24558 44546 24610 44558
rect 24558 44482 24610 44494
rect 24670 44546 24722 44558
rect 24670 44482 24722 44494
rect 24894 44546 24946 44558
rect 24894 44482 24946 44494
rect 25006 44546 25058 44558
rect 25006 44482 25058 44494
rect 27694 44546 27746 44558
rect 27694 44482 27746 44494
rect 28142 44546 28194 44558
rect 30046 44546 30098 44558
rect 28578 44494 28590 44546
rect 28642 44543 28654 44546
rect 28802 44543 28814 44546
rect 28642 44497 28814 44543
rect 28642 44494 28654 44497
rect 28802 44494 28814 44497
rect 28866 44494 28878 44546
rect 36082 44494 36094 44546
rect 36146 44494 36158 44546
rect 56690 44494 56702 44546
rect 56754 44494 56766 44546
rect 28142 44482 28194 44494
rect 30046 44482 30098 44494
rect 3166 44434 3218 44446
rect 13806 44434 13858 44446
rect 25790 44434 25842 44446
rect 4386 44382 4398 44434
rect 4450 44382 4462 44434
rect 10658 44382 10670 44434
rect 10722 44382 10734 44434
rect 14914 44382 14926 44434
rect 14978 44382 14990 44434
rect 20850 44382 20862 44434
rect 20914 44382 20926 44434
rect 3166 44370 3218 44382
rect 13806 44370 13858 44382
rect 25790 44370 25842 44382
rect 27918 44434 27970 44446
rect 27918 44370 27970 44382
rect 30382 44434 30434 44446
rect 39902 44434 39954 44446
rect 35970 44382 35982 44434
rect 36034 44382 36046 44434
rect 37874 44382 37886 44434
rect 37938 44382 37950 44434
rect 30382 44370 30434 44382
rect 39902 44370 39954 44382
rect 40238 44434 40290 44446
rect 40238 44370 40290 44382
rect 44270 44434 44322 44446
rect 49086 44434 49138 44446
rect 45826 44382 45838 44434
rect 45890 44382 45902 44434
rect 48290 44382 48302 44434
rect 48354 44382 48366 44434
rect 44270 44370 44322 44382
rect 49086 44370 49138 44382
rect 49758 44434 49810 44446
rect 51998 44434 52050 44446
rect 57710 44434 57762 44446
rect 51090 44382 51102 44434
rect 51154 44382 51166 44434
rect 56578 44382 56590 44434
rect 56642 44382 56654 44434
rect 49758 44370 49810 44382
rect 51998 44370 52050 44382
rect 57710 44370 57762 44382
rect 5966 44322 6018 44334
rect 2706 44270 2718 44322
rect 2770 44270 2782 44322
rect 2930 44270 2942 44322
rect 2994 44270 3006 44322
rect 4274 44270 4286 44322
rect 4338 44270 4350 44322
rect 5966 44258 6018 44270
rect 6414 44322 6466 44334
rect 6414 44258 6466 44270
rect 8430 44322 8482 44334
rect 11790 44322 11842 44334
rect 14814 44322 14866 44334
rect 10322 44270 10334 44322
rect 10386 44270 10398 44322
rect 11218 44270 11230 44322
rect 11282 44270 11294 44322
rect 12002 44270 12014 44322
rect 12066 44270 12078 44322
rect 14354 44270 14366 44322
rect 14418 44270 14430 44322
rect 8430 44258 8482 44270
rect 11790 44258 11842 44270
rect 14814 44258 14866 44270
rect 15822 44322 15874 44334
rect 15822 44258 15874 44270
rect 16046 44322 16098 44334
rect 16046 44258 16098 44270
rect 17726 44322 17778 44334
rect 17726 44258 17778 44270
rect 18174 44322 18226 44334
rect 18174 44258 18226 44270
rect 18286 44322 18338 44334
rect 18286 44258 18338 44270
rect 19070 44322 19122 44334
rect 19070 44258 19122 44270
rect 21646 44322 21698 44334
rect 22094 44322 22146 44334
rect 26462 44322 26514 44334
rect 21858 44270 21870 44322
rect 21922 44270 21934 44322
rect 22194 44270 22206 44322
rect 22258 44270 22270 44322
rect 21646 44258 21698 44270
rect 22094 44258 22146 44270
rect 26462 44258 26514 44270
rect 27022 44322 27074 44334
rect 31502 44322 31554 44334
rect 33406 44322 33458 44334
rect 38782 44322 38834 44334
rect 27458 44270 27470 44322
rect 27522 44270 27534 44322
rect 31826 44270 31838 44322
rect 31890 44270 31902 44322
rect 34738 44270 34750 44322
rect 34802 44270 34814 44322
rect 35298 44270 35310 44322
rect 35362 44270 35374 44322
rect 38210 44270 38222 44322
rect 38274 44270 38286 44322
rect 27022 44258 27074 44270
rect 31502 44258 31554 44270
rect 33406 44258 33458 44270
rect 38782 44258 38834 44270
rect 41246 44322 41298 44334
rect 41246 44258 41298 44270
rect 41582 44322 41634 44334
rect 41582 44258 41634 44270
rect 42590 44322 42642 44334
rect 44158 44322 44210 44334
rect 42802 44270 42814 44322
rect 42866 44270 42878 44322
rect 42590 44258 42642 44270
rect 44158 44258 44210 44270
rect 44382 44322 44434 44334
rect 46622 44322 46674 44334
rect 49870 44322 49922 44334
rect 46162 44270 46174 44322
rect 46226 44270 46238 44322
rect 48402 44270 48414 44322
rect 48466 44270 48478 44322
rect 44382 44258 44434 44270
rect 46622 44258 46674 44270
rect 49870 44258 49922 44270
rect 50094 44322 50146 44334
rect 51314 44270 51326 44322
rect 51378 44270 51390 44322
rect 56802 44270 56814 44322
rect 56866 44270 56878 44322
rect 50094 44258 50146 44270
rect 4958 44210 5010 44222
rect 4050 44158 4062 44210
rect 4114 44158 4126 44210
rect 4958 44146 5010 44158
rect 5742 44210 5794 44222
rect 14926 44210 14978 44222
rect 8978 44158 8990 44210
rect 9042 44158 9054 44210
rect 9202 44158 9214 44210
rect 9266 44158 9278 44210
rect 10434 44158 10446 44210
rect 10498 44158 10510 44210
rect 5742 44146 5794 44158
rect 14926 44146 14978 44158
rect 19182 44210 19234 44222
rect 19182 44146 19234 44158
rect 19518 44210 19570 44222
rect 19518 44146 19570 44158
rect 20302 44210 20354 44222
rect 20302 44146 20354 44158
rect 20414 44210 20466 44222
rect 26350 44210 26402 44222
rect 20514 44158 20526 44210
rect 20578 44158 20590 44210
rect 20414 44146 20466 44158
rect 26350 44146 26402 44158
rect 29486 44210 29538 44222
rect 29486 44146 29538 44158
rect 30158 44210 30210 44222
rect 30158 44146 30210 44158
rect 39678 44210 39730 44222
rect 39678 44146 39730 44158
rect 41358 44210 41410 44222
rect 41358 44146 41410 44158
rect 43486 44210 43538 44222
rect 43486 44146 43538 44158
rect 44718 44210 44770 44222
rect 44718 44146 44770 44158
rect 49646 44210 49698 44222
rect 49646 44146 49698 44158
rect 7422 44098 7474 44110
rect 7422 44034 7474 44046
rect 7870 44098 7922 44110
rect 11902 44098 11954 44110
rect 8530 44046 8542 44098
rect 8594 44046 8606 44098
rect 7870 44034 7922 44046
rect 11902 44034 11954 44046
rect 14590 44098 14642 44110
rect 16830 44098 16882 44110
rect 16370 44046 16382 44098
rect 16434 44046 16446 44098
rect 14590 44034 14642 44046
rect 16830 44034 16882 44046
rect 17278 44098 17330 44110
rect 17278 44034 17330 44046
rect 18398 44098 18450 44110
rect 18398 44034 18450 44046
rect 19406 44098 19458 44110
rect 19406 44034 19458 44046
rect 20078 44098 20130 44110
rect 22990 44098 23042 44110
rect 22082 44046 22094 44098
rect 22146 44046 22158 44098
rect 20078 44034 20130 44046
rect 22990 44034 23042 44046
rect 23550 44098 23602 44110
rect 23550 44034 23602 44046
rect 23886 44098 23938 44110
rect 23886 44034 23938 44046
rect 26574 44098 26626 44110
rect 26574 44034 26626 44046
rect 27582 44098 27634 44110
rect 27582 44034 27634 44046
rect 28814 44098 28866 44110
rect 28814 44034 28866 44046
rect 30830 44098 30882 44110
rect 30830 44034 30882 44046
rect 42030 44098 42082 44110
rect 42030 44034 42082 44046
rect 1344 43930 59024 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 59024 43930
rect 1344 43844 59024 43878
rect 1934 43762 1986 43774
rect 1934 43698 1986 43710
rect 5294 43762 5346 43774
rect 5294 43698 5346 43710
rect 8206 43762 8258 43774
rect 8206 43698 8258 43710
rect 9886 43762 9938 43774
rect 9886 43698 9938 43710
rect 12574 43762 12626 43774
rect 12574 43698 12626 43710
rect 14702 43762 14754 43774
rect 14702 43698 14754 43710
rect 16830 43762 16882 43774
rect 16830 43698 16882 43710
rect 17950 43762 18002 43774
rect 17950 43698 18002 43710
rect 26014 43762 26066 43774
rect 26014 43698 26066 43710
rect 26462 43762 26514 43774
rect 26462 43698 26514 43710
rect 28030 43762 28082 43774
rect 28030 43698 28082 43710
rect 28142 43762 28194 43774
rect 28142 43698 28194 43710
rect 28254 43762 28306 43774
rect 28254 43698 28306 43710
rect 30270 43762 30322 43774
rect 30270 43698 30322 43710
rect 35422 43762 35474 43774
rect 35422 43698 35474 43710
rect 38222 43762 38274 43774
rect 38222 43698 38274 43710
rect 44494 43762 44546 43774
rect 44494 43698 44546 43710
rect 45502 43762 45554 43774
rect 45502 43698 45554 43710
rect 56590 43762 56642 43774
rect 56590 43698 56642 43710
rect 5070 43650 5122 43662
rect 5070 43586 5122 43598
rect 5406 43650 5458 43662
rect 5406 43586 5458 43598
rect 9774 43650 9826 43662
rect 11454 43650 11506 43662
rect 10434 43598 10446 43650
rect 10498 43598 10510 43650
rect 9774 43586 9826 43598
rect 11454 43586 11506 43598
rect 12238 43650 12290 43662
rect 13470 43650 13522 43662
rect 16606 43650 16658 43662
rect 12338 43598 12350 43650
rect 12402 43598 12414 43650
rect 16258 43598 16270 43650
rect 16322 43598 16334 43650
rect 12238 43586 12290 43598
rect 13470 43586 13522 43598
rect 16606 43586 16658 43598
rect 18062 43650 18114 43662
rect 23998 43650 24050 43662
rect 20850 43598 20862 43650
rect 20914 43598 20926 43650
rect 18062 43586 18114 43598
rect 23998 43586 24050 43598
rect 24558 43650 24610 43662
rect 24558 43586 24610 43598
rect 28478 43650 28530 43662
rect 28478 43586 28530 43598
rect 31054 43650 31106 43662
rect 39678 43650 39730 43662
rect 43934 43650 43986 43662
rect 34514 43598 34526 43650
rect 34578 43598 34590 43650
rect 40338 43598 40350 43650
rect 40402 43598 40414 43650
rect 31054 43586 31106 43598
rect 39678 43586 39730 43598
rect 43934 43586 43986 43598
rect 56366 43650 56418 43662
rect 56366 43586 56418 43598
rect 57486 43650 57538 43662
rect 57486 43586 57538 43598
rect 5518 43538 5570 43550
rect 3154 43486 3166 43538
rect 3218 43486 3230 43538
rect 3714 43486 3726 43538
rect 3778 43486 3790 43538
rect 5518 43474 5570 43486
rect 6750 43538 6802 43550
rect 6750 43474 6802 43486
rect 7646 43538 7698 43550
rect 12910 43538 12962 43550
rect 10658 43486 10670 43538
rect 10722 43486 10734 43538
rect 12002 43486 12014 43538
rect 12066 43486 12078 43538
rect 7646 43474 7698 43486
rect 12910 43474 12962 43486
rect 14366 43538 14418 43550
rect 14366 43474 14418 43486
rect 14702 43538 14754 43550
rect 14702 43474 14754 43486
rect 15038 43538 15090 43550
rect 18734 43538 18786 43550
rect 16370 43486 16382 43538
rect 16434 43486 16446 43538
rect 17714 43486 17726 43538
rect 17778 43486 17790 43538
rect 15038 43474 15090 43486
rect 18734 43474 18786 43486
rect 18958 43538 19010 43550
rect 27918 43538 27970 43550
rect 35086 43538 35138 43550
rect 20402 43486 20414 43538
rect 20466 43486 20478 43538
rect 21634 43486 21646 43538
rect 21698 43486 21710 43538
rect 32834 43486 32846 43538
rect 32898 43486 32910 43538
rect 34290 43486 34302 43538
rect 34354 43486 34366 43538
rect 18958 43474 19010 43486
rect 27918 43474 27970 43486
rect 35086 43474 35138 43486
rect 35982 43538 36034 43550
rect 35982 43474 36034 43486
rect 37326 43538 37378 43550
rect 41582 43538 41634 43550
rect 54126 43538 54178 43550
rect 56254 43538 56306 43550
rect 40562 43486 40574 43538
rect 40626 43486 40638 43538
rect 42242 43486 42254 43538
rect 42306 43486 42318 43538
rect 55010 43486 55022 43538
rect 55074 43486 55086 43538
rect 56018 43486 56030 43538
rect 56082 43486 56094 43538
rect 37326 43474 37378 43486
rect 41582 43474 41634 43486
rect 54126 43474 54178 43486
rect 56254 43474 56306 43486
rect 56478 43538 56530 43550
rect 57922 43486 57934 43538
rect 57986 43486 57998 43538
rect 56478 43474 56530 43486
rect 2494 43426 2546 43438
rect 2494 43362 2546 43374
rect 4174 43426 4226 43438
rect 4174 43362 4226 43374
rect 6302 43426 6354 43438
rect 6302 43362 6354 43374
rect 7198 43426 7250 43438
rect 7198 43362 7250 43374
rect 8542 43426 8594 43438
rect 8542 43362 8594 43374
rect 8990 43426 9042 43438
rect 8990 43362 9042 43374
rect 9998 43426 10050 43438
rect 9998 43362 10050 43374
rect 13022 43426 13074 43438
rect 13022 43362 13074 43374
rect 13918 43426 13970 43438
rect 13918 43362 13970 43374
rect 15486 43426 15538 43438
rect 19182 43426 19234 43438
rect 16482 43374 16494 43426
rect 16546 43374 16558 43426
rect 18834 43374 18846 43426
rect 18898 43374 18910 43426
rect 15486 43362 15538 43374
rect 19182 43362 19234 43374
rect 19406 43426 19458 43438
rect 19406 43362 19458 43374
rect 21086 43426 21138 43438
rect 21086 43362 21138 43374
rect 21198 43426 21250 43438
rect 21198 43362 21250 43374
rect 22766 43426 22818 43438
rect 22766 43362 22818 43374
rect 23102 43426 23154 43438
rect 23102 43362 23154 43374
rect 23662 43426 23714 43438
rect 23662 43362 23714 43374
rect 25006 43426 25058 43438
rect 25006 43362 25058 43374
rect 26798 43426 26850 43438
rect 26798 43362 26850 43374
rect 27246 43426 27298 43438
rect 27246 43362 27298 43374
rect 29262 43426 29314 43438
rect 29262 43362 29314 43374
rect 29710 43426 29762 43438
rect 29710 43362 29762 43374
rect 33518 43426 33570 43438
rect 33518 43362 33570 43374
rect 36542 43426 36594 43438
rect 36542 43362 36594 43374
rect 36878 43426 36930 43438
rect 36878 43362 36930 43374
rect 37886 43426 37938 43438
rect 37886 43362 37938 43374
rect 38670 43426 38722 43438
rect 38670 43362 38722 43374
rect 39118 43426 39170 43438
rect 44942 43426 44994 43438
rect 40786 43374 40798 43426
rect 40850 43374 40862 43426
rect 42354 43374 42366 43426
rect 42418 43374 42430 43426
rect 44034 43374 44046 43426
rect 44098 43374 44110 43426
rect 39118 43362 39170 43374
rect 44942 43362 44994 43374
rect 46062 43426 46114 43438
rect 46062 43362 46114 43374
rect 46622 43426 46674 43438
rect 46622 43362 46674 43374
rect 46958 43426 47010 43438
rect 46958 43362 47010 43374
rect 47406 43426 47458 43438
rect 47406 43362 47458 43374
rect 47854 43426 47906 43438
rect 47854 43362 47906 43374
rect 48414 43426 48466 43438
rect 48414 43362 48466 43374
rect 48862 43426 48914 43438
rect 54898 43374 54910 43426
rect 54962 43374 54974 43426
rect 58370 43374 58382 43426
rect 58434 43374 58446 43426
rect 48862 43362 48914 43374
rect 10222 43314 10274 43326
rect 4050 43262 4062 43314
rect 4114 43262 4126 43314
rect 7186 43262 7198 43314
rect 7250 43311 7262 43314
rect 8866 43311 8878 43314
rect 7250 43265 8878 43311
rect 7250 43262 7262 43265
rect 8866 43262 8878 43265
rect 8930 43262 8942 43314
rect 10222 43250 10274 43262
rect 19630 43314 19682 43326
rect 31278 43314 31330 43326
rect 23650 43262 23662 43314
rect 23714 43311 23726 43314
rect 25106 43311 25118 43314
rect 23714 43265 25118 43311
rect 23714 43262 23726 43265
rect 25106 43262 25118 43265
rect 25170 43262 25182 43314
rect 19630 43250 19682 43262
rect 31278 43250 31330 43262
rect 31614 43314 31666 43326
rect 31614 43250 31666 43262
rect 32510 43314 32562 43326
rect 32510 43250 32562 43262
rect 32846 43314 32898 43326
rect 43710 43314 43762 43326
rect 38770 43262 38782 43314
rect 38834 43311 38846 43314
rect 39106 43311 39118 43314
rect 38834 43265 39118 43311
rect 38834 43262 38846 43265
rect 39106 43262 39118 43265
rect 39170 43262 39182 43314
rect 42802 43262 42814 43314
rect 42866 43262 42878 43314
rect 44258 43262 44270 43314
rect 44322 43311 44334 43314
rect 45042 43311 45054 43314
rect 44322 43265 45054 43311
rect 44322 43262 44334 43265
rect 45042 43262 45054 43265
rect 45106 43262 45118 43314
rect 32846 43250 32898 43262
rect 43710 43250 43762 43262
rect 1344 43146 59024 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 59024 43146
rect 1344 43060 59024 43094
rect 12126 42978 12178 42990
rect 6626 42926 6638 42978
rect 6690 42926 6702 42978
rect 12126 42914 12178 42926
rect 22094 42978 22146 42990
rect 29934 42978 29986 42990
rect 45838 42978 45890 42990
rect 27682 42926 27694 42978
rect 27746 42975 27758 42978
rect 28242 42975 28254 42978
rect 27746 42929 28254 42975
rect 27746 42926 27758 42929
rect 28242 42926 28254 42929
rect 28306 42926 28318 42978
rect 36194 42926 36206 42978
rect 36258 42926 36270 42978
rect 45490 42926 45502 42978
rect 45554 42926 45566 42978
rect 22094 42914 22146 42926
rect 29934 42914 29986 42926
rect 45838 42914 45890 42926
rect 48974 42978 49026 42990
rect 48974 42914 49026 42926
rect 2158 42866 2210 42878
rect 2158 42802 2210 42814
rect 2606 42866 2658 42878
rect 2606 42802 2658 42814
rect 2942 42866 2994 42878
rect 10334 42866 10386 42878
rect 15150 42866 15202 42878
rect 18398 42866 18450 42878
rect 26686 42866 26738 42878
rect 3602 42814 3614 42866
rect 3666 42814 3678 42866
rect 14242 42814 14254 42866
rect 14306 42814 14318 42866
rect 15922 42814 15934 42866
rect 15986 42814 15998 42866
rect 17826 42814 17838 42866
rect 17890 42814 17902 42866
rect 18722 42814 18734 42866
rect 18786 42814 18798 42866
rect 25106 42814 25118 42866
rect 25170 42814 25182 42866
rect 25890 42814 25902 42866
rect 25954 42814 25966 42866
rect 2942 42802 2994 42814
rect 10334 42802 10386 42814
rect 15150 42802 15202 42814
rect 18398 42802 18450 42814
rect 26686 42802 26738 42814
rect 27918 42866 27970 42878
rect 40462 42866 40514 42878
rect 35746 42814 35758 42866
rect 35810 42814 35822 42866
rect 27918 42802 27970 42814
rect 40462 42802 40514 42814
rect 47742 42866 47794 42878
rect 47742 42802 47794 42814
rect 53902 42866 53954 42878
rect 53902 42802 53954 42814
rect 55022 42866 55074 42878
rect 55022 42802 55074 42814
rect 56702 42866 56754 42878
rect 56702 42802 56754 42814
rect 4062 42754 4114 42766
rect 4062 42690 4114 42702
rect 6078 42754 6130 42766
rect 6078 42690 6130 42702
rect 6414 42754 6466 42766
rect 8094 42754 8146 42766
rect 8766 42754 8818 42766
rect 6850 42702 6862 42754
rect 6914 42702 6926 42754
rect 8530 42702 8542 42754
rect 8594 42702 8606 42754
rect 6414 42690 6466 42702
rect 8094 42690 8146 42702
rect 8766 42690 8818 42702
rect 8990 42754 9042 42766
rect 11790 42754 11842 42766
rect 9202 42702 9214 42754
rect 9266 42702 9278 42754
rect 8990 42690 9042 42702
rect 11790 42690 11842 42702
rect 13918 42754 13970 42766
rect 15710 42754 15762 42766
rect 14354 42702 14366 42754
rect 14418 42702 14430 42754
rect 13918 42690 13970 42702
rect 15710 42690 15762 42702
rect 17054 42754 17106 42766
rect 21982 42754 22034 42766
rect 26798 42754 26850 42766
rect 17714 42702 17726 42754
rect 17778 42702 17790 42754
rect 22194 42702 22206 42754
rect 22258 42702 22270 42754
rect 23650 42702 23662 42754
rect 23714 42702 23726 42754
rect 23986 42702 23998 42754
rect 24050 42702 24062 42754
rect 26114 42702 26126 42754
rect 26178 42702 26190 42754
rect 17054 42690 17106 42702
rect 21982 42690 22034 42702
rect 26798 42690 26850 42702
rect 28814 42754 28866 42766
rect 33070 42754 33122 42766
rect 38110 42754 38162 42766
rect 31938 42702 31950 42754
rect 32002 42702 32014 42754
rect 33282 42702 33294 42754
rect 33346 42702 33358 42754
rect 34402 42702 34414 42754
rect 34466 42702 34478 42754
rect 35298 42702 35310 42754
rect 35362 42702 35374 42754
rect 28814 42690 28866 42702
rect 33070 42690 33122 42702
rect 38110 42690 38162 42702
rect 38894 42754 38946 42766
rect 46062 42754 46114 42766
rect 39106 42702 39118 42754
rect 39170 42702 39182 42754
rect 38894 42690 38946 42702
rect 46062 42690 46114 42702
rect 48750 42754 48802 42766
rect 48750 42690 48802 42702
rect 53342 42754 53394 42766
rect 53342 42690 53394 42702
rect 54014 42754 54066 42766
rect 54014 42690 54066 42702
rect 55582 42754 55634 42766
rect 55582 42690 55634 42702
rect 55918 42754 55970 42766
rect 55918 42690 55970 42702
rect 7758 42642 7810 42654
rect 7758 42578 7810 42590
rect 7870 42642 7922 42654
rect 7870 42578 7922 42590
rect 9886 42642 9938 42654
rect 13694 42642 13746 42654
rect 11106 42590 11118 42642
rect 11170 42590 11182 42642
rect 11554 42590 11566 42642
rect 11618 42590 11630 42642
rect 9886 42578 9938 42590
rect 13694 42578 13746 42590
rect 14142 42642 14194 42654
rect 14142 42578 14194 42590
rect 16046 42642 16098 42654
rect 17278 42642 17330 42654
rect 16146 42590 16158 42642
rect 16210 42590 16222 42642
rect 16046 42578 16098 42590
rect 17278 42578 17330 42590
rect 17390 42642 17442 42654
rect 17390 42578 17442 42590
rect 19966 42642 20018 42654
rect 19966 42578 20018 42590
rect 21646 42642 21698 42654
rect 21646 42578 21698 42590
rect 23102 42642 23154 42654
rect 23102 42578 23154 42590
rect 25902 42642 25954 42654
rect 25902 42578 25954 42590
rect 30046 42642 30098 42654
rect 30046 42578 30098 42590
rect 37774 42642 37826 42654
rect 37774 42578 37826 42590
rect 39790 42642 39842 42654
rect 39790 42578 39842 42590
rect 40350 42642 40402 42654
rect 40350 42578 40402 42590
rect 54910 42642 54962 42654
rect 54910 42578 54962 42590
rect 56254 42642 56306 42654
rect 56254 42578 56306 42590
rect 3502 42530 3554 42542
rect 3502 42466 3554 42478
rect 3726 42530 3778 42542
rect 3726 42466 3778 42478
rect 4622 42530 4674 42542
rect 4622 42466 4674 42478
rect 5070 42530 5122 42542
rect 8878 42530 8930 42542
rect 6514 42478 6526 42530
rect 6578 42478 6590 42530
rect 5070 42466 5122 42478
rect 8878 42466 8930 42478
rect 13022 42530 13074 42542
rect 13022 42466 13074 42478
rect 15934 42530 15986 42542
rect 15934 42466 15986 42478
rect 18622 42530 18674 42542
rect 18622 42466 18674 42478
rect 19518 42530 19570 42542
rect 19518 42466 19570 42478
rect 20414 42530 20466 42542
rect 20414 42466 20466 42478
rect 20862 42530 20914 42542
rect 20862 42466 20914 42478
rect 22430 42530 22482 42542
rect 22430 42466 22482 42478
rect 26350 42530 26402 42542
rect 26350 42466 26402 42478
rect 27470 42530 27522 42542
rect 27470 42466 27522 42478
rect 28366 42530 28418 42542
rect 28366 42466 28418 42478
rect 29934 42530 29986 42542
rect 29934 42466 29986 42478
rect 30830 42530 30882 42542
rect 30830 42466 30882 42478
rect 37886 42530 37938 42542
rect 37886 42466 37938 42478
rect 40574 42530 40626 42542
rect 40574 42466 40626 42478
rect 40798 42530 40850 42542
rect 40798 42466 40850 42478
rect 41358 42530 41410 42542
rect 41358 42466 41410 42478
rect 41806 42530 41858 42542
rect 41806 42466 41858 42478
rect 42702 42530 42754 42542
rect 42702 42466 42754 42478
rect 43374 42530 43426 42542
rect 43374 42466 43426 42478
rect 44718 42530 44770 42542
rect 44718 42466 44770 42478
rect 46510 42530 46562 42542
rect 46510 42466 46562 42478
rect 47406 42530 47458 42542
rect 47406 42466 47458 42478
rect 47630 42530 47682 42542
rect 47630 42466 47682 42478
rect 47854 42530 47906 42542
rect 47854 42466 47906 42478
rect 48302 42530 48354 42542
rect 48302 42466 48354 42478
rect 49086 42530 49138 42542
rect 49086 42466 49138 42478
rect 49310 42530 49362 42542
rect 49310 42466 49362 42478
rect 49758 42530 49810 42542
rect 49758 42466 49810 42478
rect 52222 42530 52274 42542
rect 52222 42466 52274 42478
rect 53790 42530 53842 42542
rect 53790 42466 53842 42478
rect 55134 42530 55186 42542
rect 55134 42466 55186 42478
rect 56142 42530 56194 42542
rect 56142 42466 56194 42478
rect 57150 42530 57202 42542
rect 57150 42466 57202 42478
rect 57598 42530 57650 42542
rect 57598 42466 57650 42478
rect 1344 42362 59024 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 59024 42362
rect 1344 42276 59024 42310
rect 3726 42194 3778 42206
rect 3726 42130 3778 42142
rect 10110 42194 10162 42206
rect 10110 42130 10162 42142
rect 10670 42194 10722 42206
rect 10670 42130 10722 42142
rect 13358 42194 13410 42206
rect 13358 42130 13410 42142
rect 13470 42194 13522 42206
rect 13470 42130 13522 42142
rect 13582 42194 13634 42206
rect 13582 42130 13634 42142
rect 14926 42194 14978 42206
rect 14926 42130 14978 42142
rect 17950 42194 18002 42206
rect 17950 42130 18002 42142
rect 19518 42194 19570 42206
rect 19518 42130 19570 42142
rect 19630 42194 19682 42206
rect 37438 42194 37490 42206
rect 32834 42142 32846 42194
rect 32898 42142 32910 42194
rect 19630 42130 19682 42142
rect 37438 42130 37490 42142
rect 37550 42194 37602 42206
rect 37550 42130 37602 42142
rect 37662 42194 37714 42206
rect 37662 42130 37714 42142
rect 38446 42194 38498 42206
rect 38446 42130 38498 42142
rect 44718 42194 44770 42206
rect 44718 42130 44770 42142
rect 53342 42194 53394 42206
rect 53342 42130 53394 42142
rect 2494 42082 2546 42094
rect 2494 42018 2546 42030
rect 2718 42082 2770 42094
rect 2718 42018 2770 42030
rect 3054 42082 3106 42094
rect 3054 42018 3106 42030
rect 3614 42082 3666 42094
rect 8766 42082 8818 42094
rect 6626 42030 6638 42082
rect 6690 42030 6702 42082
rect 3614 42018 3666 42030
rect 8766 42018 8818 42030
rect 21758 42082 21810 42094
rect 30830 42082 30882 42094
rect 26562 42030 26574 42082
rect 26626 42030 26638 42082
rect 29586 42030 29598 42082
rect 29650 42030 29662 42082
rect 21758 42018 21810 42030
rect 30830 42018 30882 42030
rect 31166 42082 31218 42094
rect 31166 42018 31218 42030
rect 36542 42082 36594 42094
rect 36542 42018 36594 42030
rect 37102 42082 37154 42094
rect 37102 42018 37154 42030
rect 37326 42082 37378 42094
rect 37326 42018 37378 42030
rect 38334 42082 38386 42094
rect 38334 42018 38386 42030
rect 42366 42082 42418 42094
rect 42366 42018 42418 42030
rect 48750 42082 48802 42094
rect 48750 42018 48802 42030
rect 53902 42082 53954 42094
rect 53902 42018 53954 42030
rect 57486 42082 57538 42094
rect 57486 42018 57538 42030
rect 3950 41970 4002 41982
rect 3950 41906 4002 41918
rect 4174 41970 4226 41982
rect 8542 41970 8594 41982
rect 6514 41918 6526 41970
rect 6578 41918 6590 41970
rect 7410 41918 7422 41970
rect 7474 41918 7486 41970
rect 4174 41906 4226 41918
rect 8542 41906 8594 41918
rect 9662 41970 9714 41982
rect 9662 41906 9714 41918
rect 11230 41970 11282 41982
rect 11230 41906 11282 41918
rect 12014 41970 12066 41982
rect 12014 41906 12066 41918
rect 12910 41970 12962 41982
rect 12910 41906 12962 41918
rect 14142 41970 14194 41982
rect 14142 41906 14194 41918
rect 14590 41970 14642 41982
rect 14590 41906 14642 41918
rect 14814 41970 14866 41982
rect 14814 41906 14866 41918
rect 15038 41970 15090 41982
rect 15038 41906 15090 41918
rect 15598 41970 15650 41982
rect 15598 41906 15650 41918
rect 16494 41970 16546 41982
rect 19742 41970 19794 41982
rect 19282 41918 19294 41970
rect 19346 41918 19358 41970
rect 16494 41906 16546 41918
rect 19742 41906 19794 41918
rect 19854 41970 19906 41982
rect 19854 41906 19906 41918
rect 20862 41970 20914 41982
rect 20862 41906 20914 41918
rect 21086 41970 21138 41982
rect 21086 41906 21138 41918
rect 21870 41970 21922 41982
rect 21870 41906 21922 41918
rect 21982 41970 22034 41982
rect 22878 41970 22930 41982
rect 30718 41970 30770 41982
rect 22418 41918 22430 41970
rect 22482 41918 22494 41970
rect 23650 41918 23662 41970
rect 23714 41918 23726 41970
rect 24210 41918 24222 41970
rect 24274 41918 24286 41970
rect 26674 41918 26686 41970
rect 26738 41918 26750 41970
rect 28354 41918 28366 41970
rect 28418 41918 28430 41970
rect 29026 41918 29038 41970
rect 29090 41918 29102 41970
rect 21982 41906 22034 41918
rect 22878 41906 22930 41918
rect 30718 41906 30770 41918
rect 33854 41970 33906 41982
rect 38670 41970 38722 41982
rect 44606 41970 44658 41982
rect 34066 41918 34078 41970
rect 34130 41918 34142 41970
rect 35858 41918 35870 41970
rect 35922 41918 35934 41970
rect 40114 41918 40126 41970
rect 40178 41918 40190 41970
rect 43362 41918 43374 41970
rect 43426 41918 43438 41970
rect 33854 41906 33906 41918
rect 38670 41906 38722 41918
rect 44606 41906 44658 41918
rect 44942 41970 44994 41982
rect 44942 41906 44994 41918
rect 45726 41970 45778 41982
rect 45726 41906 45778 41918
rect 46398 41970 46450 41982
rect 48638 41970 48690 41982
rect 52670 41970 52722 41982
rect 57598 41970 57650 41982
rect 48290 41918 48302 41970
rect 48354 41918 48366 41970
rect 50082 41918 50094 41970
rect 50146 41918 50158 41970
rect 51090 41918 51102 41970
rect 51154 41918 51166 41970
rect 56354 41918 56366 41970
rect 56418 41918 56430 41970
rect 57922 41918 57934 41970
rect 57986 41918 57998 41970
rect 46398 41906 46450 41918
rect 48638 41906 48690 41918
rect 52670 41906 52722 41918
rect 57598 41906 57650 41918
rect 2046 41858 2098 41870
rect 1698 41806 1710 41858
rect 1762 41806 1774 41858
rect 1713 41743 1759 41806
rect 2046 41794 2098 41806
rect 2942 41858 2994 41870
rect 2942 41794 2994 41806
rect 4958 41858 5010 41870
rect 4958 41794 5010 41806
rect 5518 41858 5570 41870
rect 5518 41794 5570 41806
rect 5966 41858 6018 41870
rect 7198 41858 7250 41870
rect 12574 41858 12626 41870
rect 6962 41806 6974 41858
rect 7026 41806 7038 41858
rect 8866 41806 8878 41858
rect 8930 41806 8942 41858
rect 5966 41794 6018 41806
rect 7198 41794 7250 41806
rect 12574 41794 12626 41806
rect 14366 41858 14418 41870
rect 14366 41794 14418 41806
rect 16046 41858 16098 41870
rect 16046 41794 16098 41806
rect 16942 41858 16994 41870
rect 16942 41794 16994 41806
rect 17838 41858 17890 41870
rect 17838 41794 17890 41806
rect 18846 41858 18898 41870
rect 25902 41858 25954 41870
rect 31054 41858 31106 41870
rect 24098 41806 24110 41858
rect 24162 41806 24174 41858
rect 27682 41806 27694 41858
rect 27746 41806 27758 41858
rect 28914 41806 28926 41858
rect 28978 41806 28990 41858
rect 18846 41794 18898 41806
rect 25902 41794 25954 41806
rect 31054 41794 31106 41806
rect 31726 41858 31778 41870
rect 31726 41794 31778 41806
rect 32286 41858 32338 41870
rect 39342 41858 39394 41870
rect 41470 41858 41522 41870
rect 35634 41806 35646 41858
rect 35698 41806 35710 41858
rect 39778 41806 39790 41858
rect 39842 41806 39854 41858
rect 32286 41794 32338 41806
rect 39342 41794 39394 41806
rect 41470 41794 41522 41806
rect 43150 41858 43202 41870
rect 43150 41794 43202 41806
rect 43822 41858 43874 41870
rect 43822 41794 43874 41806
rect 45278 41858 45330 41870
rect 49970 41806 49982 41858
rect 50034 41806 50046 41858
rect 56242 41806 56254 41858
rect 56306 41806 56318 41858
rect 45278 41794 45330 41806
rect 17726 41746 17778 41758
rect 2370 41743 2382 41746
rect 1713 41697 2382 41743
rect 2370 41694 2382 41697
rect 2434 41694 2446 41746
rect 17726 41682 17778 41694
rect 20526 41746 20578 41758
rect 32510 41746 32562 41758
rect 42142 41746 42194 41758
rect 24546 41694 24558 41746
rect 24610 41694 24622 41746
rect 34514 41694 34526 41746
rect 34578 41694 34590 41746
rect 20526 41682 20578 41694
rect 32510 41682 32562 41694
rect 42142 41682 42194 41694
rect 42478 41746 42530 41758
rect 42478 41682 42530 41694
rect 43038 41746 43090 41758
rect 43038 41682 43090 41694
rect 46622 41746 46674 41758
rect 46622 41682 46674 41694
rect 46846 41746 46898 41758
rect 46846 41682 46898 41694
rect 47294 41746 47346 41758
rect 52446 41746 52498 41758
rect 51762 41694 51774 41746
rect 51826 41694 51838 41746
rect 47294 41682 47346 41694
rect 52446 41682 52498 41694
rect 53006 41746 53058 41758
rect 53006 41682 53058 41694
rect 53230 41746 53282 41758
rect 53230 41682 53282 41694
rect 54014 41746 54066 41758
rect 54014 41682 54066 41694
rect 54238 41746 54290 41758
rect 54238 41682 54290 41694
rect 54462 41746 54514 41758
rect 54462 41682 54514 41694
rect 54574 41746 54626 41758
rect 55906 41694 55918 41746
rect 55970 41694 55982 41746
rect 54574 41682 54626 41694
rect 1344 41578 59024 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 59024 41578
rect 1344 41492 59024 41526
rect 3054 41410 3106 41422
rect 2258 41358 2270 41410
rect 2322 41407 2334 41410
rect 2818 41407 2830 41410
rect 2322 41361 2830 41407
rect 2322 41358 2334 41361
rect 2818 41358 2830 41361
rect 2882 41358 2894 41410
rect 3054 41346 3106 41358
rect 3614 41410 3666 41422
rect 8878 41410 8930 41422
rect 24446 41410 24498 41422
rect 6962 41358 6974 41410
rect 7026 41358 7038 41410
rect 10546 41358 10558 41410
rect 10610 41407 10622 41410
rect 11106 41407 11118 41410
rect 10610 41361 11118 41407
rect 10610 41358 10622 41361
rect 11106 41358 11118 41361
rect 11170 41358 11182 41410
rect 12002 41358 12014 41410
rect 12066 41407 12078 41410
rect 12786 41407 12798 41410
rect 12066 41361 12798 41407
rect 12066 41358 12078 41361
rect 12786 41358 12798 41361
rect 12850 41358 12862 41410
rect 14802 41358 14814 41410
rect 14866 41358 14878 41410
rect 17378 41358 17390 41410
rect 17442 41407 17454 41410
rect 17602 41407 17614 41410
rect 17442 41361 17614 41407
rect 17442 41358 17454 41361
rect 17602 41358 17614 41361
rect 17666 41358 17678 41410
rect 3614 41346 3666 41358
rect 8878 41346 8930 41358
rect 24446 41346 24498 41358
rect 24670 41410 24722 41422
rect 24670 41346 24722 41358
rect 27918 41410 27970 41422
rect 27918 41346 27970 41358
rect 28030 41410 28082 41422
rect 28030 41346 28082 41358
rect 28254 41410 28306 41422
rect 28254 41346 28306 41358
rect 34190 41410 34242 41422
rect 34190 41346 34242 41358
rect 34526 41410 34578 41422
rect 34526 41346 34578 41358
rect 44494 41410 44546 41422
rect 44494 41346 44546 41358
rect 48638 41410 48690 41422
rect 48638 41346 48690 41358
rect 50206 41410 50258 41422
rect 50206 41346 50258 41358
rect 53790 41410 53842 41422
rect 54686 41410 54738 41422
rect 54338 41358 54350 41410
rect 54402 41358 54414 41410
rect 53790 41346 53842 41358
rect 54686 41346 54738 41358
rect 3838 41298 3890 41310
rect 11566 41298 11618 41310
rect 7074 41246 7086 41298
rect 7138 41246 7150 41298
rect 9874 41246 9886 41298
rect 9938 41246 9950 41298
rect 3838 41234 3890 41246
rect 11566 41234 11618 41246
rect 12462 41298 12514 41310
rect 12462 41234 12514 41246
rect 15486 41298 15538 41310
rect 15486 41234 15538 41246
rect 17390 41298 17442 41310
rect 17390 41234 17442 41246
rect 17726 41298 17778 41310
rect 17726 41234 17778 41246
rect 18622 41298 18674 41310
rect 18622 41234 18674 41246
rect 19630 41298 19682 41310
rect 19630 41234 19682 41246
rect 20190 41298 20242 41310
rect 20190 41234 20242 41246
rect 20862 41298 20914 41310
rect 20862 41234 20914 41246
rect 23214 41298 23266 41310
rect 23214 41234 23266 41246
rect 23774 41298 23826 41310
rect 36542 41298 36594 41310
rect 28802 41246 28814 41298
rect 28866 41246 28878 41298
rect 30930 41246 30942 41298
rect 30994 41246 31006 41298
rect 23774 41234 23826 41246
rect 36542 41234 36594 41246
rect 39566 41298 39618 41310
rect 53678 41298 53730 41310
rect 46946 41246 46958 41298
rect 47010 41246 47022 41298
rect 39566 41234 39618 41246
rect 53678 41234 53730 41246
rect 54910 41298 54962 41310
rect 54910 41234 54962 41246
rect 55358 41298 55410 41310
rect 55358 41234 55410 41246
rect 56590 41298 56642 41310
rect 56590 41234 56642 41246
rect 57262 41298 57314 41310
rect 57262 41234 57314 41246
rect 3278 41186 3330 41198
rect 3278 41122 3330 41134
rect 4510 41186 4562 41198
rect 4510 41122 4562 41134
rect 5630 41186 5682 41198
rect 5630 41122 5682 41134
rect 8990 41186 9042 41198
rect 10670 41186 10722 41198
rect 9538 41134 9550 41186
rect 9602 41134 9614 41186
rect 8990 41122 9042 41134
rect 10670 41122 10722 41134
rect 14142 41186 14194 41198
rect 14142 41122 14194 41134
rect 19294 41186 19346 41198
rect 19294 41122 19346 41134
rect 19406 41186 19458 41198
rect 19406 41122 19458 41134
rect 24334 41186 24386 41198
rect 24334 41122 24386 41134
rect 27246 41186 27298 41198
rect 35982 41186 36034 41198
rect 29922 41134 29934 41186
rect 29986 41134 29998 41186
rect 32274 41134 32286 41186
rect 32338 41134 32350 41186
rect 33618 41134 33630 41186
rect 33682 41134 33694 41186
rect 27246 41122 27298 41134
rect 35982 41122 36034 41134
rect 36206 41186 36258 41198
rect 36206 41122 36258 41134
rect 36430 41186 36482 41198
rect 36430 41122 36482 41134
rect 37662 41186 37714 41198
rect 39454 41186 39506 41198
rect 37874 41134 37886 41186
rect 37938 41134 37950 41186
rect 37662 41122 37714 41134
rect 39454 41122 39506 41134
rect 39678 41186 39730 41198
rect 40462 41186 40514 41198
rect 40002 41134 40014 41186
rect 40066 41134 40078 41186
rect 39678 41122 39730 41134
rect 40462 41122 40514 41134
rect 43934 41186 43986 41198
rect 57150 41186 57202 41198
rect 46162 41134 46174 41186
rect 46226 41134 46238 41186
rect 48066 41134 48078 41186
rect 48130 41134 48142 41186
rect 49186 41134 49198 41186
rect 49250 41134 49262 41186
rect 49410 41134 49422 41186
rect 49474 41134 49486 41186
rect 53890 41134 53902 41186
rect 53954 41183 53966 41186
rect 54114 41183 54126 41186
rect 53954 41137 54126 41183
rect 53954 41134 53966 41137
rect 54114 41134 54126 41137
rect 54178 41134 54190 41186
rect 43934 41122 43986 41134
rect 57150 41122 57202 41134
rect 57374 41186 57426 41198
rect 57374 41122 57426 41134
rect 2606 41074 2658 41086
rect 2606 41010 2658 41022
rect 6078 41074 6130 41086
rect 9214 41074 9266 41086
rect 7410 41022 7422 41074
rect 7474 41022 7486 41074
rect 6078 41010 6130 41022
rect 9214 41010 9266 41022
rect 9774 41074 9826 41086
rect 9774 41010 9826 41022
rect 12910 41074 12962 41086
rect 12910 41010 12962 41022
rect 14254 41074 14306 41086
rect 14254 41010 14306 41022
rect 14366 41074 14418 41086
rect 14366 41010 14418 41022
rect 16942 41074 16994 41086
rect 16942 41010 16994 41022
rect 19742 41074 19794 41086
rect 38558 41074 38610 41086
rect 25218 41022 25230 41074
rect 25282 41022 25294 41074
rect 26450 41022 26462 41074
rect 26514 41022 26526 41074
rect 26786 41022 26798 41074
rect 26850 41022 26862 41074
rect 30146 41022 30158 41074
rect 30210 41022 30222 41074
rect 33506 41022 33518 41074
rect 33570 41022 33582 41074
rect 19742 41010 19794 41022
rect 38558 41010 38610 41022
rect 40798 41074 40850 41086
rect 40798 41010 40850 41022
rect 43598 41074 43650 41086
rect 43598 41010 43650 41022
rect 44382 41074 44434 41086
rect 50094 41074 50146 41086
rect 47394 41022 47406 41074
rect 47458 41022 47470 41074
rect 44382 41010 44434 41022
rect 50094 41010 50146 41022
rect 2046 40962 2098 40974
rect 2046 40898 2098 40910
rect 3950 40962 4002 40974
rect 3950 40898 4002 40910
rect 5070 40962 5122 40974
rect 5070 40898 5122 40910
rect 8318 40962 8370 40974
rect 8318 40898 8370 40910
rect 11230 40962 11282 40974
rect 11230 40898 11282 40910
rect 12014 40962 12066 40974
rect 12014 40898 12066 40910
rect 15934 40962 15986 40974
rect 15934 40898 15986 40910
rect 16382 40962 16434 40974
rect 16382 40898 16434 40910
rect 18174 40962 18226 40974
rect 18174 40898 18226 40910
rect 21534 40962 21586 40974
rect 21534 40898 21586 40910
rect 22318 40962 22370 40974
rect 22318 40898 22370 40910
rect 22766 40962 22818 40974
rect 32846 40962 32898 40974
rect 27122 40910 27134 40962
rect 27186 40910 27198 40962
rect 22766 40898 22818 40910
rect 32846 40898 32898 40910
rect 35198 40962 35250 40974
rect 35198 40898 35250 40910
rect 36654 40962 36706 40974
rect 36654 40898 36706 40910
rect 40686 40962 40738 40974
rect 40686 40898 40738 40910
rect 41246 40962 41298 40974
rect 41246 40898 41298 40910
rect 41806 40962 41858 40974
rect 41806 40898 41858 40910
rect 42142 40962 42194 40974
rect 42142 40898 42194 40910
rect 42702 40962 42754 40974
rect 42702 40898 42754 40910
rect 43150 40962 43202 40974
rect 43150 40898 43202 40910
rect 43710 40962 43762 40974
rect 43710 40898 43762 40910
rect 44494 40962 44546 40974
rect 44494 40898 44546 40910
rect 45502 40962 45554 40974
rect 45502 40898 45554 40910
rect 50206 40962 50258 40974
rect 50206 40898 50258 40910
rect 50766 40962 50818 40974
rect 50766 40898 50818 40910
rect 51214 40962 51266 40974
rect 51214 40898 51266 40910
rect 51886 40962 51938 40974
rect 51886 40898 51938 40910
rect 52670 40962 52722 40974
rect 52670 40898 52722 40910
rect 53566 40962 53618 40974
rect 53566 40898 53618 40910
rect 55806 40962 55858 40974
rect 55806 40898 55858 40910
rect 57598 40962 57650 40974
rect 57598 40898 57650 40910
rect 1344 40794 59024 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 59024 40794
rect 1344 40708 59024 40742
rect 2942 40626 2994 40638
rect 2942 40562 2994 40574
rect 4286 40626 4338 40638
rect 4286 40562 4338 40574
rect 4734 40626 4786 40638
rect 4734 40562 4786 40574
rect 5518 40626 5570 40638
rect 5518 40562 5570 40574
rect 6414 40626 6466 40638
rect 6414 40562 6466 40574
rect 6974 40626 7026 40638
rect 6974 40562 7026 40574
rect 8878 40626 8930 40638
rect 8878 40562 8930 40574
rect 11678 40626 11730 40638
rect 11678 40562 11730 40574
rect 13694 40626 13746 40638
rect 13694 40562 13746 40574
rect 13918 40626 13970 40638
rect 13918 40562 13970 40574
rect 14478 40626 14530 40638
rect 14478 40562 14530 40574
rect 15038 40626 15090 40638
rect 15038 40562 15090 40574
rect 17726 40626 17778 40638
rect 17726 40562 17778 40574
rect 18734 40626 18786 40638
rect 18734 40562 18786 40574
rect 19182 40626 19234 40638
rect 19182 40562 19234 40574
rect 19630 40626 19682 40638
rect 19630 40562 19682 40574
rect 21310 40626 21362 40638
rect 21310 40562 21362 40574
rect 21422 40626 21474 40638
rect 21422 40562 21474 40574
rect 22206 40626 22258 40638
rect 22206 40562 22258 40574
rect 25566 40626 25618 40638
rect 25566 40562 25618 40574
rect 27806 40626 27858 40638
rect 27806 40562 27858 40574
rect 28030 40626 28082 40638
rect 28030 40562 28082 40574
rect 29038 40626 29090 40638
rect 29038 40562 29090 40574
rect 30830 40626 30882 40638
rect 30830 40562 30882 40574
rect 32286 40626 32338 40638
rect 32286 40562 32338 40574
rect 35982 40626 36034 40638
rect 35982 40562 36034 40574
rect 37774 40626 37826 40638
rect 50990 40626 51042 40638
rect 42578 40574 42590 40626
rect 42642 40574 42654 40626
rect 37774 40562 37826 40574
rect 50990 40562 51042 40574
rect 54126 40626 54178 40638
rect 54126 40562 54178 40574
rect 54462 40626 54514 40638
rect 54462 40562 54514 40574
rect 57486 40626 57538 40638
rect 57486 40562 57538 40574
rect 1822 40514 1874 40526
rect 1822 40450 1874 40462
rect 5742 40514 5794 40526
rect 5742 40450 5794 40462
rect 11230 40514 11282 40526
rect 13022 40514 13074 40526
rect 11442 40462 11454 40514
rect 11506 40462 11518 40514
rect 11230 40450 11282 40462
rect 13022 40450 13074 40462
rect 15262 40514 15314 40526
rect 15262 40450 15314 40462
rect 16382 40514 16434 40526
rect 16382 40450 16434 40462
rect 16494 40514 16546 40526
rect 16494 40450 16546 40462
rect 16942 40514 16994 40526
rect 16942 40450 16994 40462
rect 22654 40514 22706 40526
rect 27694 40514 27746 40526
rect 24882 40462 24894 40514
rect 24946 40462 24958 40514
rect 22654 40450 22706 40462
rect 27694 40450 27746 40462
rect 29598 40514 29650 40526
rect 29598 40450 29650 40462
rect 31502 40514 31554 40526
rect 31502 40450 31554 40462
rect 38446 40514 38498 40526
rect 46846 40514 46898 40526
rect 43026 40462 43038 40514
rect 43090 40462 43102 40514
rect 38446 40450 38498 40462
rect 46846 40450 46898 40462
rect 48302 40514 48354 40526
rect 48302 40450 48354 40462
rect 48526 40514 48578 40526
rect 48526 40450 48578 40462
rect 50766 40514 50818 40526
rect 50766 40450 50818 40462
rect 57710 40514 57762 40526
rect 57710 40450 57762 40462
rect 58270 40514 58322 40526
rect 58270 40450 58322 40462
rect 5070 40402 5122 40414
rect 2258 40350 2270 40402
rect 2322 40350 2334 40402
rect 5070 40338 5122 40350
rect 5854 40402 5906 40414
rect 5854 40338 5906 40350
rect 7758 40402 7810 40414
rect 7758 40338 7810 40350
rect 8318 40402 8370 40414
rect 8318 40338 8370 40350
rect 8766 40402 8818 40414
rect 8766 40338 8818 40350
rect 8990 40402 9042 40414
rect 12014 40402 12066 40414
rect 10546 40350 10558 40402
rect 10610 40350 10622 40402
rect 8990 40338 9042 40350
rect 12014 40338 12066 40350
rect 12126 40402 12178 40414
rect 12126 40338 12178 40350
rect 13582 40402 13634 40414
rect 13582 40338 13634 40350
rect 14366 40402 14418 40414
rect 14366 40338 14418 40350
rect 14702 40402 14754 40414
rect 14702 40338 14754 40350
rect 15374 40402 15426 40414
rect 15374 40338 15426 40350
rect 16606 40402 16658 40414
rect 16606 40338 16658 40350
rect 18062 40402 18114 40414
rect 18062 40338 18114 40350
rect 18510 40402 18562 40414
rect 18510 40338 18562 40350
rect 20750 40402 20802 40414
rect 20750 40338 20802 40350
rect 21198 40402 21250 40414
rect 26574 40402 26626 40414
rect 23314 40350 23326 40402
rect 23378 40350 23390 40402
rect 23650 40350 23662 40402
rect 23714 40350 23726 40402
rect 21198 40338 21250 40350
rect 26574 40338 26626 40350
rect 26798 40402 26850 40414
rect 29822 40402 29874 40414
rect 27122 40350 27134 40402
rect 27186 40350 27198 40402
rect 26798 40338 26850 40350
rect 29822 40338 29874 40350
rect 32846 40402 32898 40414
rect 32846 40338 32898 40350
rect 33518 40402 33570 40414
rect 34526 40402 34578 40414
rect 34290 40350 34302 40402
rect 34354 40350 34366 40402
rect 33518 40338 33570 40350
rect 34526 40338 34578 40350
rect 34638 40402 34690 40414
rect 34638 40338 34690 40350
rect 36430 40402 36482 40414
rect 36430 40338 36482 40350
rect 37326 40402 37378 40414
rect 37326 40338 37378 40350
rect 38894 40402 38946 40414
rect 48190 40402 48242 40414
rect 39218 40350 39230 40402
rect 39282 40350 39294 40402
rect 40002 40350 40014 40402
rect 40066 40350 40078 40402
rect 42130 40350 42142 40402
rect 42194 40350 42206 40402
rect 44258 40350 44270 40402
rect 44322 40350 44334 40402
rect 45602 40350 45614 40402
rect 45666 40350 45678 40402
rect 38894 40338 38946 40350
rect 48190 40338 48242 40350
rect 49534 40402 49586 40414
rect 49534 40338 49586 40350
rect 49982 40402 50034 40414
rect 49982 40338 50034 40350
rect 50654 40402 50706 40414
rect 50654 40338 50706 40350
rect 53566 40402 53618 40414
rect 53566 40338 53618 40350
rect 57822 40402 57874 40414
rect 57822 40338 57874 40350
rect 3502 40290 3554 40302
rect 3502 40226 3554 40238
rect 9774 40290 9826 40302
rect 12574 40290 12626 40302
rect 11106 40238 11118 40290
rect 11170 40238 11182 40290
rect 9774 40226 9826 40238
rect 12574 40226 12626 40238
rect 15934 40290 15986 40302
rect 18622 40290 18674 40302
rect 18162 40287 18174 40290
rect 15934 40226 15986 40238
rect 17841 40241 18174 40287
rect 7086 40178 7138 40190
rect 7086 40114 7138 40126
rect 7310 40178 7362 40190
rect 7310 40114 7362 40126
rect 7870 40178 7922 40190
rect 7870 40114 7922 40126
rect 10222 40178 10274 40190
rect 10222 40114 10274 40126
rect 10558 40178 10610 40190
rect 17490 40126 17502 40178
rect 17554 40175 17566 40178
rect 17841 40175 17887 40241
rect 18162 40238 18174 40241
rect 18226 40238 18238 40290
rect 18622 40226 18674 40238
rect 20078 40290 20130 40302
rect 20078 40226 20130 40238
rect 26126 40290 26178 40302
rect 26126 40226 26178 40238
rect 28702 40290 28754 40302
rect 31726 40290 31778 40302
rect 31378 40238 31390 40290
rect 31442 40238 31454 40290
rect 28702 40226 28754 40238
rect 31726 40226 31778 40238
rect 35646 40290 35698 40302
rect 35646 40226 35698 40238
rect 36878 40290 36930 40302
rect 43822 40290 43874 40302
rect 39890 40238 39902 40290
rect 39954 40238 39966 40290
rect 44594 40238 44606 40290
rect 44658 40238 44670 40290
rect 45714 40238 45726 40290
rect 45778 40238 45790 40290
rect 36878 40226 36930 40238
rect 43822 40226 43874 40238
rect 47070 40178 47122 40190
rect 17554 40129 17887 40175
rect 17554 40126 17566 40129
rect 19506 40126 19518 40178
rect 19570 40175 19582 40178
rect 19954 40175 19966 40178
rect 19570 40129 19966 40175
rect 19570 40126 19582 40129
rect 19954 40126 19966 40129
rect 20018 40126 20030 40178
rect 28690 40126 28702 40178
rect 28754 40175 28766 40178
rect 29138 40175 29150 40178
rect 28754 40129 29150 40175
rect 28754 40126 28766 40129
rect 29138 40126 29150 40129
rect 29202 40126 29214 40178
rect 30146 40126 30158 40178
rect 30210 40126 30222 40178
rect 35074 40126 35086 40178
rect 35138 40126 35150 40178
rect 36194 40126 36206 40178
rect 36258 40175 36270 40178
rect 36866 40175 36878 40178
rect 36258 40129 36878 40175
rect 36258 40126 36270 40129
rect 36866 40126 36878 40129
rect 36930 40126 36942 40178
rect 40226 40126 40238 40178
rect 40290 40126 40302 40178
rect 46050 40126 46062 40178
rect 46114 40126 46126 40178
rect 10558 40114 10610 40126
rect 47070 40114 47122 40126
rect 47406 40178 47458 40190
rect 47406 40114 47458 40126
rect 1344 40010 59024 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 59024 40010
rect 1344 39924 59024 39958
rect 2718 39842 2770 39854
rect 9774 39842 9826 39854
rect 3490 39790 3502 39842
rect 3554 39839 3566 39842
rect 4722 39839 4734 39842
rect 3554 39793 4734 39839
rect 3554 39790 3566 39793
rect 4722 39790 4734 39793
rect 4786 39790 4798 39842
rect 2718 39778 2770 39790
rect 9774 39778 9826 39790
rect 11566 39842 11618 39854
rect 42814 39842 42866 39854
rect 34738 39790 34750 39842
rect 34802 39790 34814 39842
rect 11566 39778 11618 39790
rect 42814 39778 42866 39790
rect 2494 39730 2546 39742
rect 2494 39666 2546 39678
rect 3614 39730 3666 39742
rect 3614 39666 3666 39678
rect 4062 39730 4114 39742
rect 4062 39666 4114 39678
rect 4958 39730 5010 39742
rect 4958 39666 5010 39678
rect 5630 39730 5682 39742
rect 5630 39666 5682 39678
rect 7758 39730 7810 39742
rect 7758 39666 7810 39678
rect 8766 39730 8818 39742
rect 8766 39666 8818 39678
rect 9214 39730 9266 39742
rect 12910 39730 12962 39742
rect 16158 39730 16210 39742
rect 10770 39678 10782 39730
rect 10834 39678 10846 39730
rect 15026 39678 15038 39730
rect 15090 39678 15102 39730
rect 9214 39666 9266 39678
rect 12910 39666 12962 39678
rect 16158 39666 16210 39678
rect 18622 39730 18674 39742
rect 18622 39666 18674 39678
rect 19966 39730 20018 39742
rect 19966 39666 20018 39678
rect 22878 39730 22930 39742
rect 25678 39730 25730 39742
rect 38558 39730 38610 39742
rect 25106 39678 25118 39730
rect 25170 39678 25182 39730
rect 27234 39678 27246 39730
rect 27298 39678 27310 39730
rect 28466 39678 28478 39730
rect 28530 39678 28542 39730
rect 34402 39678 34414 39730
rect 34466 39678 34478 39730
rect 22878 39666 22930 39678
rect 25678 39666 25730 39678
rect 38558 39666 38610 39678
rect 40462 39730 40514 39742
rect 42030 39730 42082 39742
rect 41122 39678 41134 39730
rect 41186 39678 41198 39730
rect 40462 39666 40514 39678
rect 42030 39666 42082 39678
rect 42590 39730 42642 39742
rect 42590 39666 42642 39678
rect 43150 39730 43202 39742
rect 45502 39730 45554 39742
rect 43810 39678 43822 39730
rect 43874 39678 43886 39730
rect 43150 39666 43202 39678
rect 45502 39666 45554 39678
rect 50878 39730 50930 39742
rect 50878 39666 50930 39678
rect 7646 39618 7698 39630
rect 7646 39554 7698 39566
rect 7870 39618 7922 39630
rect 7870 39554 7922 39566
rect 9886 39618 9938 39630
rect 10670 39618 10722 39630
rect 10434 39566 10446 39618
rect 10498 39566 10510 39618
rect 9886 39554 9938 39566
rect 10670 39554 10722 39566
rect 11790 39618 11842 39630
rect 15374 39618 15426 39630
rect 12002 39566 12014 39618
rect 12066 39566 12078 39618
rect 14578 39566 14590 39618
rect 14642 39566 14654 39618
rect 14914 39566 14926 39618
rect 14978 39566 14990 39618
rect 11790 39554 11842 39566
rect 15374 39554 15426 39566
rect 16718 39618 16770 39630
rect 16718 39554 16770 39566
rect 16830 39618 16882 39630
rect 16830 39554 16882 39566
rect 17614 39618 17666 39630
rect 19406 39618 19458 39630
rect 18274 39566 18286 39618
rect 18338 39566 18350 39618
rect 17614 39554 17666 39566
rect 19406 39554 19458 39566
rect 20974 39618 21026 39630
rect 20974 39554 21026 39566
rect 21758 39618 21810 39630
rect 21758 39554 21810 39566
rect 22318 39618 22370 39630
rect 29822 39618 29874 39630
rect 31726 39618 31778 39630
rect 36094 39618 36146 39630
rect 23538 39566 23550 39618
rect 23602 39566 23614 39618
rect 23874 39566 23886 39618
rect 23938 39566 23950 39618
rect 27010 39566 27022 39618
rect 27074 39566 27086 39618
rect 30482 39566 30494 39618
rect 30546 39566 30558 39618
rect 32162 39566 32174 39618
rect 32226 39566 32238 39618
rect 35074 39566 35086 39618
rect 35138 39566 35150 39618
rect 22318 39554 22370 39566
rect 29822 39554 29874 39566
rect 31726 39554 31778 39566
rect 36094 39554 36146 39566
rect 36430 39618 36482 39630
rect 45726 39618 45778 39630
rect 50318 39618 50370 39630
rect 41570 39566 41582 39618
rect 41634 39566 41646 39618
rect 44258 39566 44270 39618
rect 44322 39566 44334 39618
rect 47282 39566 47294 39618
rect 47346 39566 47358 39618
rect 36430 39554 36482 39566
rect 45726 39554 45778 39566
rect 50318 39554 50370 39566
rect 51438 39618 51490 39630
rect 57150 39618 57202 39630
rect 53890 39566 53902 39618
rect 53954 39566 53966 39618
rect 51438 39554 51490 39566
rect 57150 39554 57202 39566
rect 57374 39618 57426 39630
rect 57810 39566 57822 39618
rect 57874 39566 57886 39618
rect 57374 39554 57426 39566
rect 4622 39506 4674 39518
rect 4622 39442 4674 39454
rect 6190 39506 6242 39518
rect 6190 39442 6242 39454
rect 6302 39506 6354 39518
rect 6302 39442 6354 39454
rect 7422 39506 7474 39518
rect 7422 39442 7474 39454
rect 10110 39506 10162 39518
rect 10110 39442 10162 39454
rect 11454 39506 11506 39518
rect 11454 39442 11506 39454
rect 12462 39506 12514 39518
rect 12462 39442 12514 39454
rect 17166 39506 17218 39518
rect 18734 39506 18786 39518
rect 17378 39454 17390 39506
rect 17442 39454 17454 39506
rect 17166 39442 17218 39454
rect 18734 39442 18786 39454
rect 19854 39506 19906 39518
rect 19854 39442 19906 39454
rect 21870 39506 21922 39518
rect 21870 39442 21922 39454
rect 35870 39506 35922 39518
rect 35870 39442 35922 39454
rect 44718 39506 44770 39518
rect 49982 39506 50034 39518
rect 47058 39454 47070 39506
rect 47122 39454 47134 39506
rect 44718 39442 44770 39454
rect 49982 39442 50034 39454
rect 53566 39506 53618 39518
rect 53566 39442 53618 39454
rect 54686 39506 54738 39518
rect 54686 39442 54738 39454
rect 2046 39394 2098 39406
rect 6526 39394 6578 39406
rect 3042 39342 3054 39394
rect 3106 39342 3118 39394
rect 2046 39330 2098 39342
rect 6526 39330 6578 39342
rect 8318 39394 8370 39406
rect 8318 39330 8370 39342
rect 13582 39394 13634 39406
rect 13582 39330 13634 39342
rect 14030 39394 14082 39406
rect 14030 39330 14082 39342
rect 15150 39394 15202 39406
rect 15150 39330 15202 39342
rect 17502 39394 17554 39406
rect 17502 39330 17554 39342
rect 18510 39394 18562 39406
rect 18510 39330 18562 39342
rect 18846 39394 18898 39406
rect 18846 39330 18898 39342
rect 20078 39394 20130 39406
rect 20078 39330 20130 39342
rect 22094 39394 22146 39406
rect 22094 39330 22146 39342
rect 26126 39394 26178 39406
rect 26126 39330 26178 39342
rect 35982 39394 36034 39406
rect 46510 39394 46562 39406
rect 50094 39394 50146 39406
rect 46050 39342 46062 39394
rect 46114 39342 46126 39394
rect 48626 39342 48638 39394
rect 48690 39342 48702 39394
rect 35982 39330 36034 39342
rect 46510 39330 46562 39342
rect 50094 39330 50146 39342
rect 50766 39394 50818 39406
rect 50766 39330 50818 39342
rect 50990 39394 51042 39406
rect 50990 39330 51042 39342
rect 53678 39394 53730 39406
rect 53678 39330 53730 39342
rect 54350 39394 54402 39406
rect 54350 39330 54402 39342
rect 54574 39394 54626 39406
rect 54574 39330 54626 39342
rect 56590 39394 56642 39406
rect 56590 39330 56642 39342
rect 1344 39226 59024 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 59024 39226
rect 1344 39140 59024 39174
rect 2382 39058 2434 39070
rect 2382 38994 2434 39006
rect 3726 39058 3778 39070
rect 3726 38994 3778 39006
rect 3838 39058 3890 39070
rect 3838 38994 3890 39006
rect 8990 39058 9042 39070
rect 8990 38994 9042 39006
rect 12462 39058 12514 39070
rect 12462 38994 12514 39006
rect 13246 39058 13298 39070
rect 13246 38994 13298 39006
rect 13694 39058 13746 39070
rect 13694 38994 13746 39006
rect 14590 39058 14642 39070
rect 14590 38994 14642 39006
rect 15486 39058 15538 39070
rect 15486 38994 15538 39006
rect 15710 39058 15762 39070
rect 15710 38994 15762 39006
rect 16046 39058 16098 39070
rect 16046 38994 16098 39006
rect 16718 39058 16770 39070
rect 16718 38994 16770 39006
rect 16830 39058 16882 39070
rect 16830 38994 16882 39006
rect 22654 39058 22706 39070
rect 22654 38994 22706 39006
rect 23102 39058 23154 39070
rect 23102 38994 23154 39006
rect 28590 39058 28642 39070
rect 28590 38994 28642 39006
rect 34078 39058 34130 39070
rect 34078 38994 34130 39006
rect 36318 39058 36370 39070
rect 36318 38994 36370 39006
rect 36654 39058 36706 39070
rect 36654 38994 36706 39006
rect 37102 39058 37154 39070
rect 37102 38994 37154 39006
rect 37550 39058 37602 39070
rect 37550 38994 37602 39006
rect 42030 39058 42082 39070
rect 42030 38994 42082 39006
rect 42590 39058 42642 39070
rect 42590 38994 42642 39006
rect 42926 39058 42978 39070
rect 42926 38994 42978 39006
rect 45502 39058 45554 39070
rect 45502 38994 45554 39006
rect 46734 39058 46786 39070
rect 46734 38994 46786 39006
rect 47182 39058 47234 39070
rect 47182 38994 47234 39006
rect 56478 39058 56530 39070
rect 56478 38994 56530 39006
rect 3614 38946 3666 38958
rect 3614 38882 3666 38894
rect 4622 38946 4674 38958
rect 4622 38882 4674 38894
rect 4846 38946 4898 38958
rect 4846 38882 4898 38894
rect 5182 38946 5234 38958
rect 5182 38882 5234 38894
rect 7310 38946 7362 38958
rect 7310 38882 7362 38894
rect 8206 38946 8258 38958
rect 8206 38882 8258 38894
rect 10894 38946 10946 38958
rect 10894 38882 10946 38894
rect 14478 38946 14530 38958
rect 14478 38882 14530 38894
rect 14814 38946 14866 38958
rect 14814 38882 14866 38894
rect 15374 38946 15426 38958
rect 15374 38882 15426 38894
rect 17726 38946 17778 38958
rect 17726 38882 17778 38894
rect 17950 38946 18002 38958
rect 17950 38882 18002 38894
rect 18286 38946 18338 38958
rect 18286 38882 18338 38894
rect 19518 38946 19570 38958
rect 23998 38946 24050 38958
rect 33630 38946 33682 38958
rect 20626 38894 20638 38946
rect 20690 38894 20702 38946
rect 27794 38894 27806 38946
rect 27858 38894 27870 38946
rect 29138 38894 29150 38946
rect 29202 38894 29214 38946
rect 19518 38882 19570 38894
rect 23998 38882 24050 38894
rect 33630 38882 33682 38894
rect 33854 38946 33906 38958
rect 33854 38882 33906 38894
rect 40798 38946 40850 38958
rect 40798 38882 40850 38894
rect 52222 38946 52274 38958
rect 52222 38882 52274 38894
rect 58494 38946 58546 38958
rect 58494 38882 58546 38894
rect 2606 38834 2658 38846
rect 2034 38782 2046 38834
rect 2098 38782 2110 38834
rect 2606 38770 2658 38782
rect 3166 38834 3218 38846
rect 3166 38770 3218 38782
rect 6078 38834 6130 38846
rect 6078 38770 6130 38782
rect 6414 38834 6466 38846
rect 6414 38770 6466 38782
rect 6750 38834 6802 38846
rect 6750 38770 6802 38782
rect 7646 38834 7698 38846
rect 7646 38770 7698 38782
rect 7758 38834 7810 38846
rect 7758 38770 7810 38782
rect 10334 38834 10386 38846
rect 10334 38770 10386 38782
rect 10670 38834 10722 38846
rect 10670 38770 10722 38782
rect 11790 38834 11842 38846
rect 11790 38770 11842 38782
rect 12014 38834 12066 38846
rect 12686 38834 12738 38846
rect 12338 38782 12350 38834
rect 12402 38782 12414 38834
rect 12014 38770 12066 38782
rect 12686 38770 12738 38782
rect 14254 38834 14306 38846
rect 19406 38834 19458 38846
rect 23550 38834 23602 38846
rect 30718 38834 30770 38846
rect 34190 38834 34242 38846
rect 35982 38834 36034 38846
rect 44942 38834 44994 38846
rect 50430 38834 50482 38846
rect 19170 38782 19182 38834
rect 19234 38782 19246 38834
rect 20514 38782 20526 38834
rect 20578 38782 20590 38834
rect 21522 38782 21534 38834
rect 21586 38782 21598 38834
rect 25778 38782 25790 38834
rect 25842 38782 25854 38834
rect 26002 38782 26014 38834
rect 26066 38782 26078 38834
rect 29698 38782 29710 38834
rect 29762 38782 29774 38834
rect 30034 38782 30046 38834
rect 30098 38782 30110 38834
rect 31714 38782 31726 38834
rect 31778 38782 31790 38834
rect 35522 38782 35534 38834
rect 35586 38782 35598 38834
rect 40114 38782 40126 38834
rect 40178 38782 40190 38834
rect 48066 38782 48078 38834
rect 48130 38782 48142 38834
rect 49858 38782 49870 38834
rect 49922 38782 49934 38834
rect 14254 38770 14306 38782
rect 19406 38770 19458 38782
rect 23550 38770 23602 38782
rect 30718 38770 30770 38782
rect 34190 38770 34242 38782
rect 35982 38770 36034 38782
rect 44942 38770 44994 38782
rect 50430 38770 50482 38782
rect 50542 38834 50594 38846
rect 51314 38782 51326 38834
rect 51378 38782 51390 38834
rect 53778 38782 53790 38834
rect 53842 38782 53854 38834
rect 54786 38782 54798 38834
rect 54850 38782 54862 38834
rect 56690 38782 56702 38834
rect 56754 38782 56766 38834
rect 57922 38782 57934 38834
rect 57986 38782 57998 38834
rect 50542 38770 50594 38782
rect 2494 38722 2546 38734
rect 2494 38658 2546 38670
rect 3390 38722 3442 38734
rect 3390 38658 3442 38670
rect 5070 38722 5122 38734
rect 5070 38658 5122 38670
rect 5630 38722 5682 38734
rect 5630 38658 5682 38670
rect 6302 38722 6354 38734
rect 6302 38658 6354 38670
rect 7982 38722 8034 38734
rect 7982 38658 8034 38670
rect 8094 38722 8146 38734
rect 8094 38658 8146 38670
rect 9774 38722 9826 38734
rect 9774 38658 9826 38670
rect 10782 38722 10834 38734
rect 16606 38722 16658 38734
rect 12562 38670 12574 38722
rect 12626 38670 12638 38722
rect 10782 38658 10834 38670
rect 16606 38658 16658 38670
rect 18174 38722 18226 38734
rect 18174 38658 18226 38670
rect 21198 38722 21250 38734
rect 21198 38658 21250 38670
rect 21310 38722 21362 38734
rect 21310 38658 21362 38670
rect 24558 38722 24610 38734
rect 24558 38658 24610 38670
rect 25006 38722 25058 38734
rect 31502 38722 31554 38734
rect 29810 38670 29822 38722
rect 29874 38670 29886 38722
rect 25006 38658 25058 38670
rect 31502 38658 31554 38670
rect 32622 38722 32674 38734
rect 38334 38722 38386 38734
rect 35186 38670 35198 38722
rect 35250 38670 35262 38722
rect 32622 38658 32674 38670
rect 38334 38658 38386 38670
rect 39342 38722 39394 38734
rect 46286 38722 46338 38734
rect 48750 38722 48802 38734
rect 56366 38722 56418 38734
rect 40338 38670 40350 38722
rect 40402 38670 40414 38722
rect 47954 38670 47966 38722
rect 48018 38670 48030 38722
rect 51426 38670 51438 38722
rect 51490 38670 51502 38722
rect 53890 38670 53902 38722
rect 53954 38670 53966 38722
rect 55570 38670 55582 38722
rect 55634 38670 55646 38722
rect 57586 38670 57598 38722
rect 57650 38670 57662 38722
rect 39342 38658 39394 38670
rect 46286 38658 46338 38670
rect 48750 38658 48802 38670
rect 56366 38658 56418 38670
rect 38446 38610 38498 38622
rect 19954 38558 19966 38610
rect 20018 38558 20030 38610
rect 31378 38558 31390 38610
rect 31442 38558 31454 38610
rect 38446 38546 38498 38558
rect 1344 38442 59024 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 59024 38442
rect 1344 38356 59024 38390
rect 8990 38274 9042 38286
rect 16270 38274 16322 38286
rect 35422 38274 35474 38286
rect 10098 38222 10110 38274
rect 10162 38271 10174 38274
rect 11218 38271 11230 38274
rect 10162 38225 11230 38271
rect 10162 38222 10174 38225
rect 11218 38222 11230 38225
rect 11282 38222 11294 38274
rect 18498 38222 18510 38274
rect 18562 38271 18574 38274
rect 19282 38271 19294 38274
rect 18562 38225 19294 38271
rect 18562 38222 18574 38225
rect 19282 38222 19294 38225
rect 19346 38222 19358 38274
rect 39218 38222 39230 38274
rect 39282 38222 39294 38274
rect 50306 38222 50318 38274
rect 50370 38222 50382 38274
rect 8990 38210 9042 38222
rect 16270 38210 16322 38222
rect 35422 38210 35474 38222
rect 2382 38162 2434 38174
rect 2382 38098 2434 38110
rect 5070 38162 5122 38174
rect 8654 38162 8706 38174
rect 7410 38110 7422 38162
rect 7474 38110 7486 38162
rect 5070 38098 5122 38110
rect 8654 38098 8706 38110
rect 10334 38162 10386 38174
rect 10334 38098 10386 38110
rect 11566 38162 11618 38174
rect 17614 38162 17666 38174
rect 15026 38110 15038 38162
rect 15090 38110 15102 38162
rect 11566 38098 11618 38110
rect 17614 38098 17666 38110
rect 18174 38162 18226 38174
rect 18174 38098 18226 38110
rect 18510 38162 18562 38174
rect 27246 38162 27298 38174
rect 36318 38162 36370 38174
rect 22642 38110 22654 38162
rect 22706 38110 22718 38162
rect 26338 38110 26350 38162
rect 26402 38110 26414 38162
rect 30594 38110 30606 38162
rect 30658 38110 30670 38162
rect 31826 38110 31838 38162
rect 31890 38110 31902 38162
rect 18510 38098 18562 38110
rect 27246 38098 27298 38110
rect 36318 38098 36370 38110
rect 2942 38050 2994 38062
rect 2942 37986 2994 37998
rect 3502 38050 3554 38062
rect 3502 37986 3554 37998
rect 4062 38050 4114 38062
rect 8542 38050 8594 38062
rect 21646 38050 21698 38062
rect 28142 38050 28194 38062
rect 34190 38050 34242 38062
rect 5730 37998 5742 38050
rect 5794 37998 5806 38050
rect 6738 37998 6750 38050
rect 6802 37998 6814 38050
rect 7634 37998 7646 38050
rect 7698 37998 7710 38050
rect 9090 37998 9102 38050
rect 9154 37998 9166 38050
rect 13906 37998 13918 38050
rect 13970 37998 13982 38050
rect 14802 37998 14814 38050
rect 14866 37998 14878 38050
rect 15922 37998 15934 38050
rect 15986 37998 15998 38050
rect 19394 37998 19406 38050
rect 19458 37998 19470 38050
rect 20514 37998 20526 38050
rect 20578 37998 20590 38050
rect 20738 37998 20750 38050
rect 20802 37998 20814 38050
rect 21858 37998 21870 38050
rect 21922 37998 21934 38050
rect 22754 37998 22766 38050
rect 22818 37998 22830 38050
rect 24098 37998 24110 38050
rect 24162 37998 24174 38050
rect 24434 37998 24446 38050
rect 24498 37998 24510 38050
rect 26562 37998 26574 38050
rect 26626 37998 26638 38050
rect 30706 37998 30718 38050
rect 30770 37998 30782 38050
rect 4062 37986 4114 37998
rect 8542 37986 8594 37998
rect 21646 37986 21698 37998
rect 28142 37986 28194 37998
rect 34190 37986 34242 37998
rect 35198 38050 35250 38062
rect 35198 37986 35250 37998
rect 38110 38050 38162 38062
rect 39006 38050 39058 38062
rect 38322 37998 38334 38050
rect 38386 37998 38398 38050
rect 38110 37986 38162 37998
rect 39006 37986 39058 37998
rect 3054 37938 3106 37950
rect 3054 37874 3106 37886
rect 3950 37938 4002 37950
rect 3950 37874 4002 37886
rect 4286 37938 4338 37950
rect 4286 37874 4338 37886
rect 4510 37938 4562 37950
rect 9774 37938 9826 37950
rect 6850 37886 6862 37938
rect 6914 37886 6926 37938
rect 7522 37886 7534 37938
rect 7586 37886 7598 37938
rect 8754 37886 8766 37938
rect 8818 37886 8830 37938
rect 4510 37874 4562 37886
rect 9774 37874 9826 37886
rect 14366 37938 14418 37950
rect 27806 37938 27858 37950
rect 15026 37886 15038 37938
rect 15090 37886 15102 37938
rect 20626 37886 20638 37938
rect 20690 37886 20702 37938
rect 22978 37886 22990 37938
rect 23042 37886 23054 37938
rect 25554 37886 25566 37938
rect 25618 37886 25630 37938
rect 14366 37874 14418 37886
rect 27806 37874 27858 37886
rect 33294 37938 33346 37950
rect 33294 37874 33346 37886
rect 33406 37938 33458 37950
rect 33406 37874 33458 37886
rect 33630 37938 33682 37950
rect 33630 37874 33682 37886
rect 34526 37938 34578 37950
rect 34526 37874 34578 37886
rect 1934 37826 1986 37838
rect 1934 37762 1986 37774
rect 3278 37826 3330 37838
rect 3278 37762 3330 37774
rect 10670 37826 10722 37838
rect 10670 37762 10722 37774
rect 11118 37826 11170 37838
rect 11118 37762 11170 37774
rect 12014 37826 12066 37838
rect 12014 37762 12066 37774
rect 12574 37826 12626 37838
rect 12574 37762 12626 37774
rect 12910 37826 12962 37838
rect 12910 37762 12962 37774
rect 16158 37826 16210 37838
rect 16158 37762 16210 37774
rect 16718 37826 16770 37838
rect 16718 37762 16770 37774
rect 17166 37826 17218 37838
rect 17166 37762 17218 37774
rect 19070 37826 19122 37838
rect 19070 37762 19122 37774
rect 27918 37826 27970 37838
rect 27918 37762 27970 37774
rect 28814 37826 28866 37838
rect 28814 37762 28866 37774
rect 29598 37826 29650 37838
rect 29598 37762 29650 37774
rect 30046 37826 30098 37838
rect 30046 37762 30098 37774
rect 32622 37826 32674 37838
rect 32622 37762 32674 37774
rect 34078 37826 34130 37838
rect 34078 37762 34130 37774
rect 34302 37826 34354 37838
rect 36654 37826 36706 37838
rect 35746 37774 35758 37826
rect 35810 37774 35822 37826
rect 34302 37762 34354 37774
rect 36654 37762 36706 37774
rect 37438 37826 37490 37838
rect 39233 37826 39279 38222
rect 40126 38162 40178 38174
rect 40126 38098 40178 38110
rect 46734 38162 46786 38174
rect 53902 38162 53954 38174
rect 56366 38162 56418 38174
rect 50754 38110 50766 38162
rect 50818 38110 50830 38162
rect 55234 38110 55246 38162
rect 55298 38110 55310 38162
rect 57810 38110 57822 38162
rect 57874 38110 57886 38162
rect 46734 38098 46786 38110
rect 53902 38098 53954 38110
rect 56366 38098 56418 38110
rect 39566 38050 39618 38062
rect 39566 37986 39618 37998
rect 40238 38050 40290 38062
rect 40238 37986 40290 37998
rect 43598 38050 43650 38062
rect 43598 37986 43650 37998
rect 44158 38050 44210 38062
rect 51550 38050 51602 38062
rect 50418 37998 50430 38050
rect 50482 37998 50494 38050
rect 44158 37986 44210 37998
rect 51550 37986 51602 37998
rect 51886 38050 51938 38062
rect 51886 37986 51938 37998
rect 53566 38050 53618 38062
rect 53566 37986 53618 37998
rect 54126 38050 54178 38062
rect 54126 37986 54178 37998
rect 56142 38050 56194 38062
rect 56142 37986 56194 37998
rect 56478 38050 56530 38062
rect 58382 38050 58434 38062
rect 57698 37998 57710 38050
rect 57762 37998 57774 38050
rect 56478 37986 56530 37998
rect 58382 37986 58434 37998
rect 51774 37938 51826 37950
rect 51774 37874 51826 37886
rect 53678 37938 53730 37950
rect 53678 37874 53730 37886
rect 54910 37938 54962 37950
rect 54910 37874 54962 37886
rect 40014 37826 40066 37838
rect 39218 37774 39230 37826
rect 39282 37774 39294 37826
rect 37438 37762 37490 37774
rect 40014 37762 40066 37774
rect 40798 37826 40850 37838
rect 40798 37762 40850 37774
rect 41246 37826 41298 37838
rect 41246 37762 41298 37774
rect 42142 37826 42194 37838
rect 42142 37762 42194 37774
rect 44046 37826 44098 37838
rect 44046 37762 44098 37774
rect 44270 37826 44322 37838
rect 44270 37762 44322 37774
rect 45726 37826 45778 37838
rect 45726 37762 45778 37774
rect 46622 37826 46674 37838
rect 46622 37762 46674 37774
rect 46846 37826 46898 37838
rect 46846 37762 46898 37774
rect 47070 37826 47122 37838
rect 47070 37762 47122 37774
rect 1344 37658 59024 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 59024 37658
rect 1344 37572 59024 37606
rect 1934 37490 1986 37502
rect 1934 37426 1986 37438
rect 10558 37490 10610 37502
rect 10558 37426 10610 37438
rect 12126 37490 12178 37502
rect 12126 37426 12178 37438
rect 17838 37490 17890 37502
rect 17838 37426 17890 37438
rect 17950 37490 18002 37502
rect 17950 37426 18002 37438
rect 19966 37490 20018 37502
rect 19966 37426 20018 37438
rect 21870 37490 21922 37502
rect 21870 37426 21922 37438
rect 22094 37490 22146 37502
rect 22094 37426 22146 37438
rect 23102 37490 23154 37502
rect 23102 37426 23154 37438
rect 23550 37490 23602 37502
rect 23550 37426 23602 37438
rect 23998 37490 24050 37502
rect 23998 37426 24050 37438
rect 24446 37490 24498 37502
rect 24446 37426 24498 37438
rect 24894 37490 24946 37502
rect 24894 37426 24946 37438
rect 25902 37490 25954 37502
rect 35310 37490 35362 37502
rect 29698 37438 29710 37490
rect 29762 37438 29774 37490
rect 32050 37438 32062 37490
rect 32114 37438 32126 37490
rect 25902 37426 25954 37438
rect 35310 37426 35362 37438
rect 38782 37490 38834 37502
rect 38782 37426 38834 37438
rect 39006 37490 39058 37502
rect 39006 37426 39058 37438
rect 41470 37490 41522 37502
rect 41470 37426 41522 37438
rect 54350 37490 54402 37502
rect 54350 37426 54402 37438
rect 54910 37490 54962 37502
rect 54910 37426 54962 37438
rect 57486 37490 57538 37502
rect 57486 37426 57538 37438
rect 3838 37378 3890 37390
rect 3838 37314 3890 37326
rect 4398 37378 4450 37390
rect 11118 37378 11170 37390
rect 8418 37326 8430 37378
rect 8482 37326 8494 37378
rect 9986 37326 9998 37378
rect 10050 37326 10062 37378
rect 4398 37314 4450 37326
rect 11118 37314 11170 37326
rect 11230 37378 11282 37390
rect 11230 37314 11282 37326
rect 13134 37378 13186 37390
rect 18062 37378 18114 37390
rect 14914 37326 14926 37378
rect 14978 37326 14990 37378
rect 13134 37314 13186 37326
rect 18062 37314 18114 37326
rect 18174 37378 18226 37390
rect 20974 37378 21026 37390
rect 18386 37326 18398 37378
rect 18450 37326 18462 37378
rect 18174 37314 18226 37326
rect 20974 37314 21026 37326
rect 21310 37378 21362 37390
rect 29150 37378 29202 37390
rect 27346 37326 27358 37378
rect 27410 37326 27422 37378
rect 21310 37314 21362 37326
rect 29150 37314 29202 37326
rect 29262 37378 29314 37390
rect 38110 37378 38162 37390
rect 34402 37326 34414 37378
rect 34466 37326 34478 37378
rect 36194 37326 36206 37378
rect 36258 37326 36270 37378
rect 29262 37314 29314 37326
rect 38110 37314 38162 37326
rect 38670 37378 38722 37390
rect 38670 37314 38722 37326
rect 45054 37378 45106 37390
rect 45054 37314 45106 37326
rect 57710 37378 57762 37390
rect 57710 37314 57762 37326
rect 57822 37378 57874 37390
rect 57822 37314 57874 37326
rect 3278 37266 3330 37278
rect 3278 37202 3330 37214
rect 3726 37266 3778 37278
rect 9774 37266 9826 37278
rect 12686 37266 12738 37278
rect 4722 37214 4734 37266
rect 4786 37214 4798 37266
rect 7074 37214 7086 37266
rect 7138 37214 7150 37266
rect 7410 37214 7422 37266
rect 7474 37214 7486 37266
rect 8194 37214 8206 37266
rect 8258 37214 8270 37266
rect 10546 37214 10558 37266
rect 10610 37214 10622 37266
rect 3726 37202 3778 37214
rect 9774 37202 9826 37214
rect 12686 37202 12738 37214
rect 12798 37266 12850 37278
rect 13582 37266 13634 37278
rect 16494 37266 16546 37278
rect 13346 37214 13358 37266
rect 13410 37214 13422 37266
rect 14802 37214 14814 37266
rect 14866 37214 14878 37266
rect 15810 37214 15822 37266
rect 15874 37214 15886 37266
rect 12798 37202 12850 37214
rect 13582 37202 13634 37214
rect 16494 37202 16546 37214
rect 20750 37266 20802 37278
rect 20750 37202 20802 37214
rect 21086 37266 21138 37278
rect 21086 37202 21138 37214
rect 21982 37266 22034 37278
rect 26350 37266 26402 37278
rect 29038 37266 29090 37278
rect 46846 37266 46898 37278
rect 22418 37214 22430 37266
rect 22482 37214 22494 37266
rect 27458 37214 27470 37266
rect 27522 37214 27534 37266
rect 27794 37214 27806 37266
rect 27858 37214 27870 37266
rect 31490 37214 31502 37266
rect 31554 37214 31566 37266
rect 31714 37214 31726 37266
rect 31778 37214 31790 37266
rect 34290 37214 34302 37266
rect 34354 37214 34366 37266
rect 37426 37214 37438 37266
rect 37490 37214 37502 37266
rect 39778 37214 39790 37266
rect 39842 37214 39854 37266
rect 42578 37214 42590 37266
rect 42642 37214 42654 37266
rect 44370 37214 44382 37266
rect 44434 37214 44446 37266
rect 46386 37214 46398 37266
rect 46450 37214 46462 37266
rect 47506 37214 47518 37266
rect 47570 37214 47582 37266
rect 21982 37202 22034 37214
rect 26350 37202 26402 37214
rect 29038 37202 29090 37214
rect 46846 37202 46898 37214
rect 2382 37154 2434 37166
rect 2382 37090 2434 37102
rect 3054 37154 3106 37166
rect 5182 37154 5234 37166
rect 3490 37102 3502 37154
rect 3554 37102 3566 37154
rect 3054 37090 3106 37102
rect 5182 37090 5234 37102
rect 5630 37154 5682 37166
rect 5630 37090 5682 37102
rect 6078 37154 6130 37166
rect 6078 37090 6130 37102
rect 6526 37154 6578 37166
rect 6526 37090 6578 37102
rect 7982 37154 8034 37166
rect 14590 37154 14642 37166
rect 13682 37102 13694 37154
rect 13746 37102 13758 37154
rect 7982 37090 8034 37102
rect 14590 37090 14642 37102
rect 19406 37154 19458 37166
rect 30158 37154 30210 37166
rect 27570 37102 27582 37154
rect 27634 37102 27646 37154
rect 19406 37090 19458 37102
rect 30158 37090 30210 37102
rect 30718 37154 30770 37166
rect 32846 37154 32898 37166
rect 32162 37102 32174 37154
rect 32226 37102 32238 37154
rect 30718 37090 30770 37102
rect 32846 37090 32898 37102
rect 33518 37154 33570 37166
rect 40574 37154 40626 37166
rect 43374 37154 43426 37166
rect 56366 37154 56418 37166
rect 34850 37102 34862 37154
rect 34914 37102 34926 37154
rect 35970 37102 35982 37154
rect 36034 37102 36046 37154
rect 39890 37102 39902 37154
rect 39954 37102 39966 37154
rect 42690 37102 42702 37154
rect 42754 37102 42766 37154
rect 44146 37102 44158 37154
rect 44210 37102 44222 37154
rect 48290 37102 48302 37154
rect 48354 37102 48366 37154
rect 33518 37090 33570 37102
rect 40574 37090 40626 37102
rect 43374 37090 43426 37102
rect 56366 37090 56418 37102
rect 56702 37154 56754 37166
rect 56702 37090 56754 37102
rect 4734 37042 4786 37054
rect 10222 37042 10274 37054
rect 5282 36990 5294 37042
rect 5346 37039 5358 37042
rect 6402 37039 6414 37042
rect 5346 36993 6414 37039
rect 5346 36990 5358 36993
rect 6402 36990 6414 36993
rect 6466 36990 6478 37042
rect 4734 36978 4786 36990
rect 10222 36978 10274 36990
rect 11230 37042 11282 37054
rect 11230 36978 11282 36990
rect 16382 37042 16434 37054
rect 16382 36978 16434 36990
rect 16718 37042 16770 37054
rect 16718 36978 16770 36990
rect 16830 37042 16882 37054
rect 20526 37042 20578 37054
rect 19394 36990 19406 37042
rect 19458 37039 19470 37042
rect 19954 37039 19966 37042
rect 19458 36993 19966 37039
rect 19458 36990 19470 36993
rect 19954 36990 19966 36993
rect 20018 36990 20030 37042
rect 24098 36990 24110 37042
rect 24162 37039 24174 37042
rect 24882 37039 24894 37042
rect 24162 36993 24894 37039
rect 24162 36990 24174 36993
rect 24882 36990 24894 36993
rect 24946 36990 24958 37042
rect 55906 36990 55918 37042
rect 55970 37039 55982 37042
rect 56354 37039 56366 37042
rect 55970 36993 56366 37039
rect 55970 36990 55982 36993
rect 56354 36990 56366 36993
rect 56418 36990 56430 37042
rect 16830 36978 16882 36990
rect 20526 36978 20578 36990
rect 1344 36874 59024 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 59024 36874
rect 1344 36788 59024 36822
rect 9998 36706 10050 36718
rect 1810 36654 1822 36706
rect 1874 36703 1886 36706
rect 2370 36703 2382 36706
rect 1874 36657 2382 36703
rect 1874 36654 1886 36657
rect 2370 36654 2382 36657
rect 2434 36654 2446 36706
rect 9998 36642 10050 36654
rect 16718 36706 16770 36718
rect 16718 36642 16770 36654
rect 17390 36706 17442 36718
rect 17390 36642 17442 36654
rect 19406 36706 19458 36718
rect 42926 36706 42978 36718
rect 20178 36654 20190 36706
rect 20242 36703 20254 36706
rect 20514 36703 20526 36706
rect 20242 36657 20526 36703
rect 20242 36654 20254 36657
rect 20514 36654 20526 36657
rect 20578 36654 20590 36706
rect 23650 36654 23662 36706
rect 23714 36703 23726 36706
rect 24322 36703 24334 36706
rect 23714 36657 24334 36703
rect 23714 36654 23726 36657
rect 24322 36654 24334 36657
rect 24386 36654 24398 36706
rect 28354 36654 28366 36706
rect 28418 36654 28430 36706
rect 31042 36654 31054 36706
rect 31106 36703 31118 36706
rect 31106 36657 31215 36703
rect 31106 36654 31118 36657
rect 19406 36642 19458 36654
rect 1822 36594 1874 36606
rect 1822 36530 1874 36542
rect 6190 36594 6242 36606
rect 6190 36530 6242 36542
rect 7870 36594 7922 36606
rect 12126 36594 12178 36606
rect 10882 36542 10894 36594
rect 10946 36542 10958 36594
rect 7870 36530 7922 36542
rect 12126 36530 12178 36542
rect 17838 36594 17890 36606
rect 17838 36530 17890 36542
rect 23662 36594 23714 36606
rect 23662 36530 23714 36542
rect 30046 36594 30098 36606
rect 31169 36591 31215 36657
rect 42926 36642 42978 36654
rect 43262 36706 43314 36718
rect 43262 36642 43314 36654
rect 43934 36706 43986 36718
rect 43934 36642 43986 36654
rect 46286 36706 46338 36718
rect 46286 36642 46338 36654
rect 31950 36594 32002 36606
rect 31490 36591 31502 36594
rect 31169 36545 31502 36591
rect 31490 36542 31502 36545
rect 31554 36542 31566 36594
rect 30046 36530 30098 36542
rect 31950 36530 32002 36542
rect 32958 36594 33010 36606
rect 32958 36530 33010 36542
rect 33966 36594 34018 36606
rect 33966 36530 34018 36542
rect 34526 36594 34578 36606
rect 34526 36530 34578 36542
rect 35870 36594 35922 36606
rect 35870 36530 35922 36542
rect 36430 36594 36482 36606
rect 36430 36530 36482 36542
rect 38782 36594 38834 36606
rect 43822 36594 43874 36606
rect 47854 36594 47906 36606
rect 41682 36542 41694 36594
rect 41746 36542 41758 36594
rect 46498 36542 46510 36594
rect 46562 36542 46574 36594
rect 38782 36530 38834 36542
rect 43822 36530 43874 36542
rect 47854 36530 47906 36542
rect 50654 36594 50706 36606
rect 50654 36530 50706 36542
rect 53902 36594 53954 36606
rect 53902 36530 53954 36542
rect 55022 36594 55074 36606
rect 57822 36594 57874 36606
rect 57474 36542 57486 36594
rect 57538 36542 57550 36594
rect 55022 36530 55074 36542
rect 57822 36530 57874 36542
rect 5966 36482 6018 36494
rect 2818 36430 2830 36482
rect 2882 36430 2894 36482
rect 4050 36430 4062 36482
rect 4114 36430 4126 36482
rect 4498 36430 4510 36482
rect 4562 36430 4574 36482
rect 5966 36418 6018 36430
rect 6526 36482 6578 36494
rect 6526 36418 6578 36430
rect 7534 36482 7586 36494
rect 7534 36418 7586 36430
rect 7982 36482 8034 36494
rect 7982 36418 8034 36430
rect 8766 36482 8818 36494
rect 8766 36418 8818 36430
rect 9326 36482 9378 36494
rect 9326 36418 9378 36430
rect 9438 36482 9490 36494
rect 9438 36418 9490 36430
rect 10110 36482 10162 36494
rect 10110 36418 10162 36430
rect 11566 36482 11618 36494
rect 17614 36482 17666 36494
rect 13906 36430 13918 36482
rect 13970 36430 13982 36482
rect 14578 36430 14590 36482
rect 14642 36430 14654 36482
rect 15474 36430 15486 36482
rect 15538 36430 15550 36482
rect 11566 36418 11618 36430
rect 17614 36418 17666 36430
rect 18174 36482 18226 36494
rect 18174 36418 18226 36430
rect 18286 36482 18338 36494
rect 19182 36482 19234 36494
rect 18946 36430 18958 36482
rect 19010 36430 19022 36482
rect 18286 36418 18338 36430
rect 19182 36418 19234 36430
rect 21534 36482 21586 36494
rect 21534 36418 21586 36430
rect 21870 36482 21922 36494
rect 21870 36418 21922 36430
rect 22766 36482 22818 36494
rect 22766 36418 22818 36430
rect 25342 36482 25394 36494
rect 25342 36418 25394 36430
rect 25902 36482 25954 36494
rect 25902 36418 25954 36430
rect 26126 36482 26178 36494
rect 29486 36482 29538 36494
rect 26562 36430 26574 36482
rect 26626 36430 26638 36482
rect 28466 36430 28478 36482
rect 28530 36430 28542 36482
rect 26126 36418 26178 36430
rect 29486 36418 29538 36430
rect 29934 36482 29986 36494
rect 29934 36418 29986 36430
rect 31838 36482 31890 36494
rect 31838 36418 31890 36430
rect 33406 36482 33458 36494
rect 33406 36418 33458 36430
rect 33854 36482 33906 36494
rect 33854 36418 33906 36430
rect 35310 36482 35362 36494
rect 35310 36418 35362 36430
rect 37886 36482 37938 36494
rect 37886 36418 37938 36430
rect 39678 36482 39730 36494
rect 39678 36418 39730 36430
rect 40014 36482 40066 36494
rect 40014 36418 40066 36430
rect 41134 36482 41186 36494
rect 41134 36418 41186 36430
rect 41358 36482 41410 36494
rect 41358 36418 41410 36430
rect 47070 36482 47122 36494
rect 47070 36418 47122 36430
rect 47406 36482 47458 36494
rect 47406 36418 47458 36430
rect 50878 36482 50930 36494
rect 50878 36418 50930 36430
rect 53342 36482 53394 36494
rect 57362 36430 57374 36482
rect 57426 36430 57438 36482
rect 53342 36418 53394 36430
rect 6414 36370 6466 36382
rect 3938 36318 3950 36370
rect 4002 36318 4014 36370
rect 4834 36318 4846 36370
rect 4898 36318 4910 36370
rect 6414 36306 6466 36318
rect 7646 36370 7698 36382
rect 10894 36370 10946 36382
rect 16718 36370 16770 36382
rect 10658 36318 10670 36370
rect 10722 36318 10734 36370
rect 13794 36318 13806 36370
rect 13858 36318 13870 36370
rect 14466 36318 14478 36370
rect 14530 36318 14542 36370
rect 7646 36306 7698 36318
rect 10894 36306 10946 36318
rect 16718 36306 16770 36318
rect 16830 36370 16882 36382
rect 16830 36306 16882 36318
rect 19966 36370 20018 36382
rect 19966 36306 20018 36318
rect 22206 36370 22258 36382
rect 22206 36306 22258 36318
rect 25006 36370 25058 36382
rect 25006 36306 25058 36318
rect 26014 36370 26066 36382
rect 30158 36370 30210 36382
rect 28802 36318 28814 36370
rect 28866 36318 28878 36370
rect 26014 36306 26066 36318
rect 30158 36306 30210 36318
rect 31614 36370 31666 36382
rect 31614 36306 31666 36318
rect 32062 36370 32114 36382
rect 32062 36306 32114 36318
rect 34078 36370 34130 36382
rect 34078 36306 34130 36318
rect 39790 36370 39842 36382
rect 39790 36306 39842 36318
rect 42702 36370 42754 36382
rect 42702 36306 42754 36318
rect 50206 36370 50258 36382
rect 50206 36306 50258 36318
rect 50430 36370 50482 36382
rect 50430 36306 50482 36318
rect 54574 36370 54626 36382
rect 54574 36306 54626 36318
rect 54798 36370 54850 36382
rect 54798 36306 54850 36318
rect 55134 36370 55186 36382
rect 55134 36306 55186 36318
rect 2270 36258 2322 36270
rect 9214 36258 9266 36270
rect 3826 36206 3838 36258
rect 3890 36206 3902 36258
rect 2270 36194 2322 36206
rect 9214 36194 9266 36206
rect 10446 36258 10498 36270
rect 10446 36194 10498 36206
rect 12910 36258 12962 36270
rect 18062 36258 18114 36270
rect 14802 36206 14814 36258
rect 14866 36206 14878 36258
rect 12910 36194 12962 36206
rect 18062 36194 18114 36206
rect 19070 36258 19122 36270
rect 19070 36194 19122 36206
rect 20414 36258 20466 36270
rect 20414 36194 20466 36206
rect 20862 36258 20914 36270
rect 20862 36194 20914 36206
rect 21758 36258 21810 36270
rect 21758 36194 21810 36206
rect 22878 36258 22930 36270
rect 22878 36194 22930 36206
rect 23102 36258 23154 36270
rect 23102 36194 23154 36206
rect 23998 36258 24050 36270
rect 23998 36194 24050 36206
rect 24446 36258 24498 36270
rect 24446 36194 24498 36206
rect 25118 36258 25170 36270
rect 25118 36194 25170 36206
rect 31054 36258 31106 36270
rect 31054 36194 31106 36206
rect 32622 36258 32674 36270
rect 32622 36194 32674 36206
rect 35758 36258 35810 36270
rect 35758 36194 35810 36206
rect 35982 36258 36034 36270
rect 35982 36194 36034 36206
rect 37438 36258 37490 36270
rect 37438 36194 37490 36206
rect 38334 36258 38386 36270
rect 38334 36194 38386 36206
rect 40462 36258 40514 36270
rect 40462 36194 40514 36206
rect 42254 36258 42306 36270
rect 42254 36194 42306 36206
rect 44382 36258 44434 36270
rect 44382 36194 44434 36206
rect 45502 36258 45554 36270
rect 45502 36194 45554 36206
rect 46510 36258 46562 36270
rect 46510 36194 46562 36206
rect 47294 36258 47346 36270
rect 47294 36194 47346 36206
rect 51214 36258 51266 36270
rect 51214 36194 51266 36206
rect 53790 36258 53842 36270
rect 53790 36194 53842 36206
rect 54014 36258 54066 36270
rect 54014 36194 54066 36206
rect 1344 36090 59024 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 59024 36090
rect 1344 36004 59024 36038
rect 7198 35922 7250 35934
rect 7198 35858 7250 35870
rect 8542 35922 8594 35934
rect 8542 35858 8594 35870
rect 8990 35922 9042 35934
rect 8990 35858 9042 35870
rect 10894 35922 10946 35934
rect 10894 35858 10946 35870
rect 11790 35922 11842 35934
rect 11790 35858 11842 35870
rect 13022 35922 13074 35934
rect 13022 35858 13074 35870
rect 13470 35922 13522 35934
rect 13470 35858 13522 35870
rect 14254 35922 14306 35934
rect 16942 35922 16994 35934
rect 15026 35870 15038 35922
rect 15090 35870 15102 35922
rect 14254 35858 14306 35870
rect 16942 35858 16994 35870
rect 18622 35922 18674 35934
rect 18622 35858 18674 35870
rect 19406 35922 19458 35934
rect 19406 35858 19458 35870
rect 20302 35922 20354 35934
rect 20302 35858 20354 35870
rect 22206 35922 22258 35934
rect 22206 35858 22258 35870
rect 26014 35922 26066 35934
rect 26014 35858 26066 35870
rect 26126 35922 26178 35934
rect 26126 35858 26178 35870
rect 26798 35922 26850 35934
rect 26798 35858 26850 35870
rect 33854 35922 33906 35934
rect 33854 35858 33906 35870
rect 34974 35922 35026 35934
rect 34974 35858 35026 35870
rect 38558 35922 38610 35934
rect 38558 35858 38610 35870
rect 39678 35922 39730 35934
rect 39678 35858 39730 35870
rect 44494 35922 44546 35934
rect 44494 35858 44546 35870
rect 45502 35922 45554 35934
rect 45502 35858 45554 35870
rect 46734 35922 46786 35934
rect 46734 35858 46786 35870
rect 49758 35922 49810 35934
rect 49758 35858 49810 35870
rect 51998 35922 52050 35934
rect 51998 35858 52050 35870
rect 57710 35922 57762 35934
rect 57710 35858 57762 35870
rect 5518 35810 5570 35822
rect 5518 35746 5570 35758
rect 13694 35810 13746 35822
rect 16046 35810 16098 35822
rect 15138 35758 15150 35810
rect 15202 35758 15214 35810
rect 13694 35746 13746 35758
rect 16046 35746 16098 35758
rect 16270 35810 16322 35822
rect 16270 35746 16322 35758
rect 17726 35810 17778 35822
rect 17726 35746 17778 35758
rect 20078 35810 20130 35822
rect 40686 35810 40738 35822
rect 30818 35758 30830 35810
rect 30882 35758 30894 35810
rect 20078 35746 20130 35758
rect 40686 35746 40738 35758
rect 43486 35810 43538 35822
rect 43486 35746 43538 35758
rect 44942 35810 44994 35822
rect 44942 35746 44994 35758
rect 45390 35810 45442 35822
rect 45390 35746 45442 35758
rect 53902 35810 53954 35822
rect 53902 35746 53954 35758
rect 56590 35810 56642 35822
rect 56590 35746 56642 35758
rect 57486 35810 57538 35822
rect 57486 35746 57538 35758
rect 4734 35698 4786 35710
rect 3378 35646 3390 35698
rect 3442 35646 3454 35698
rect 4162 35646 4174 35698
rect 4226 35646 4238 35698
rect 4734 35634 4786 35646
rect 5406 35698 5458 35710
rect 5406 35634 5458 35646
rect 5742 35698 5794 35710
rect 5742 35634 5794 35646
rect 6750 35698 6802 35710
rect 6750 35634 6802 35646
rect 10110 35698 10162 35710
rect 10110 35634 10162 35646
rect 10558 35698 10610 35710
rect 10558 35634 10610 35646
rect 10782 35698 10834 35710
rect 10782 35634 10834 35646
rect 11006 35698 11058 35710
rect 13806 35698 13858 35710
rect 16606 35698 16658 35710
rect 11890 35646 11902 35698
rect 11954 35646 11966 35698
rect 12338 35646 12350 35698
rect 12402 35646 12414 35698
rect 14914 35646 14926 35698
rect 14978 35646 14990 35698
rect 11006 35634 11058 35646
rect 13806 35634 13858 35646
rect 16606 35634 16658 35646
rect 16830 35698 16882 35710
rect 16830 35634 16882 35646
rect 17950 35698 18002 35710
rect 17950 35634 18002 35646
rect 18286 35698 18338 35710
rect 18286 35634 18338 35646
rect 20526 35698 20578 35710
rect 20526 35634 20578 35646
rect 21086 35698 21138 35710
rect 21086 35634 21138 35646
rect 21310 35698 21362 35710
rect 21310 35634 21362 35646
rect 21758 35698 21810 35710
rect 25790 35698 25842 35710
rect 23314 35646 23326 35698
rect 23378 35646 23390 35698
rect 23874 35646 23886 35698
rect 23938 35646 23950 35698
rect 21758 35634 21810 35646
rect 25790 35634 25842 35646
rect 25902 35698 25954 35710
rect 31614 35698 31666 35710
rect 26338 35646 26350 35698
rect 26402 35646 26414 35698
rect 27458 35646 27470 35698
rect 27522 35646 27534 35698
rect 27794 35646 27806 35698
rect 27858 35646 27870 35698
rect 29474 35646 29486 35698
rect 29538 35646 29550 35698
rect 30258 35646 30270 35698
rect 30322 35646 30334 35698
rect 25902 35634 25954 35646
rect 31614 35634 31666 35646
rect 31838 35698 31890 35710
rect 31838 35634 31890 35646
rect 32174 35698 32226 35710
rect 34862 35698 34914 35710
rect 34626 35646 34638 35698
rect 34690 35646 34702 35698
rect 32174 35634 32226 35646
rect 34862 35634 34914 35646
rect 35086 35698 35138 35710
rect 36878 35698 36930 35710
rect 35298 35646 35310 35698
rect 35362 35646 35374 35698
rect 35086 35634 35138 35646
rect 36878 35634 36930 35646
rect 37326 35698 37378 35710
rect 37326 35634 37378 35646
rect 37550 35698 37602 35710
rect 53006 35698 53058 35710
rect 55582 35698 55634 35710
rect 39890 35646 39902 35698
rect 39954 35646 39966 35698
rect 41794 35646 41806 35698
rect 41858 35646 41870 35698
rect 42018 35646 42030 35698
rect 42082 35646 42094 35698
rect 45714 35646 45726 35698
rect 45778 35646 45790 35698
rect 49522 35646 49534 35698
rect 49586 35646 49598 35698
rect 51090 35646 51102 35698
rect 51154 35646 51166 35698
rect 53218 35646 53230 35698
rect 53282 35646 53294 35698
rect 54786 35646 54798 35698
rect 54850 35646 54862 35698
rect 37550 35634 37602 35646
rect 53006 35634 53058 35646
rect 55582 35634 55634 35646
rect 57710 35698 57762 35710
rect 57710 35634 57762 35646
rect 57934 35698 57986 35710
rect 57934 35634 57986 35646
rect 2158 35586 2210 35598
rect 2158 35522 2210 35534
rect 2606 35586 2658 35598
rect 7646 35586 7698 35598
rect 3490 35534 3502 35586
rect 3554 35534 3566 35586
rect 6290 35534 6302 35586
rect 6354 35534 6366 35586
rect 2606 35522 2658 35534
rect 7646 35522 7698 35534
rect 8206 35586 8258 35598
rect 8206 35522 8258 35534
rect 20414 35586 20466 35598
rect 20414 35522 20466 35534
rect 21534 35586 21586 35598
rect 21534 35522 21586 35534
rect 22654 35586 22706 35598
rect 31950 35586 32002 35598
rect 24770 35534 24782 35586
rect 24834 35534 24846 35586
rect 28914 35534 28926 35586
rect 28978 35534 28990 35586
rect 30370 35534 30382 35586
rect 30434 35534 30446 35586
rect 22654 35522 22706 35534
rect 31950 35522 32002 35534
rect 32510 35586 32562 35598
rect 35758 35586 35810 35598
rect 33954 35534 33966 35586
rect 34018 35534 34030 35586
rect 32510 35522 32562 35534
rect 35758 35522 35810 35534
rect 36206 35586 36258 35598
rect 36206 35522 36258 35534
rect 37102 35586 37154 35598
rect 37102 35522 37154 35534
rect 37438 35586 37490 35598
rect 37438 35522 37490 35534
rect 38110 35586 38162 35598
rect 38110 35522 38162 35534
rect 39118 35586 39170 35598
rect 41582 35586 41634 35598
rect 40786 35534 40798 35586
rect 40850 35534 40862 35586
rect 39118 35522 39170 35534
rect 41582 35522 41634 35534
rect 43038 35586 43090 35598
rect 43038 35522 43090 35534
rect 44046 35586 44098 35598
rect 44046 35522 44098 35534
rect 46174 35586 46226 35598
rect 46174 35522 46226 35534
rect 47742 35586 47794 35598
rect 47742 35522 47794 35534
rect 48190 35586 48242 35598
rect 51550 35586 51602 35598
rect 50754 35534 50766 35586
rect 50818 35534 50830 35586
rect 54674 35534 54686 35586
rect 54738 35534 54750 35586
rect 56690 35534 56702 35586
rect 56754 35534 56766 35586
rect 48190 35522 48242 35534
rect 51550 35522 51602 35534
rect 10334 35474 10386 35486
rect 3714 35422 3726 35474
rect 3778 35422 3790 35474
rect 7858 35422 7870 35474
rect 7922 35471 7934 35474
rect 8194 35471 8206 35474
rect 7922 35425 8206 35471
rect 7922 35422 7934 35425
rect 8194 35422 8206 35425
rect 8258 35422 8270 35474
rect 10334 35410 10386 35422
rect 18510 35474 18562 35486
rect 18510 35410 18562 35422
rect 33630 35474 33682 35486
rect 33630 35410 33682 35422
rect 39566 35474 39618 35486
rect 39566 35410 39618 35422
rect 40462 35474 40514 35486
rect 40462 35410 40514 35422
rect 49870 35474 49922 35486
rect 49870 35410 49922 35422
rect 56366 35474 56418 35486
rect 56366 35410 56418 35422
rect 1344 35306 59024 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 59024 35306
rect 1344 35220 59024 35254
rect 16830 35138 16882 35150
rect 15138 35086 15150 35138
rect 15202 35135 15214 35138
rect 15698 35135 15710 35138
rect 15202 35089 15710 35135
rect 15202 35086 15214 35089
rect 15698 35086 15710 35089
rect 15762 35086 15774 35138
rect 16830 35074 16882 35086
rect 20974 35138 21026 35150
rect 28254 35138 28306 35150
rect 22642 35086 22654 35138
rect 22706 35135 22718 35138
rect 23874 35135 23886 35138
rect 22706 35089 23886 35135
rect 22706 35086 22718 35089
rect 23874 35086 23886 35089
rect 23938 35086 23950 35138
rect 20974 35074 21026 35086
rect 28254 35074 28306 35086
rect 41694 35138 41746 35150
rect 41694 35074 41746 35086
rect 1822 35026 1874 35038
rect 9662 35026 9714 35038
rect 2370 34974 2382 35026
rect 2434 34974 2446 35026
rect 4386 34974 4398 35026
rect 4450 34974 4462 35026
rect 7186 34974 7198 35026
rect 7250 34974 7262 35026
rect 1822 34962 1874 34974
rect 9662 34962 9714 34974
rect 12126 35026 12178 35038
rect 12126 34962 12178 34974
rect 14254 35026 14306 35038
rect 14254 34962 14306 34974
rect 15486 35026 15538 35038
rect 15486 34962 15538 34974
rect 16046 35026 16098 35038
rect 16046 34962 16098 34974
rect 17502 35026 17554 35038
rect 17502 34962 17554 34974
rect 18398 35026 18450 35038
rect 18398 34962 18450 34974
rect 20526 35026 20578 35038
rect 20526 34962 20578 34974
rect 21534 35026 21586 35038
rect 21534 34962 21586 34974
rect 22654 35026 22706 35038
rect 28030 35026 28082 35038
rect 37998 35026 38050 35038
rect 27010 34974 27022 35026
rect 27074 34974 27086 35026
rect 30370 34974 30382 35026
rect 30434 34974 30446 35026
rect 22654 34962 22706 34974
rect 28030 34962 28082 34974
rect 3390 34914 3442 34926
rect 3390 34850 3442 34862
rect 3502 34914 3554 34926
rect 3502 34850 3554 34862
rect 6862 34914 6914 34926
rect 6862 34850 6914 34862
rect 7310 34914 7362 34926
rect 11902 34914 11954 34926
rect 18958 34914 19010 34926
rect 10546 34862 10558 34914
rect 10610 34862 10622 34914
rect 10994 34862 11006 34914
rect 11058 34862 11070 34914
rect 13906 34862 13918 34914
rect 13970 34862 13982 34914
rect 16482 34862 16494 34914
rect 16546 34862 16558 34914
rect 7310 34850 7362 34862
rect 11902 34850 11954 34862
rect 18958 34850 19010 34862
rect 20078 34914 20130 34926
rect 20078 34850 20130 34862
rect 20302 34914 20354 34926
rect 27470 34914 27522 34926
rect 24210 34862 24222 34914
rect 24274 34862 24286 34914
rect 24546 34862 24558 34914
rect 24610 34862 24622 34914
rect 20302 34850 20354 34862
rect 27470 34850 27522 34862
rect 30046 34914 30098 34926
rect 30046 34850 30098 34862
rect 30270 34914 30322 34926
rect 30270 34850 30322 34862
rect 3838 34802 3890 34814
rect 4286 34802 4338 34814
rect 4050 34750 4062 34802
rect 4114 34750 4126 34802
rect 3838 34738 3890 34750
rect 4286 34738 4338 34750
rect 6190 34802 6242 34814
rect 6190 34738 6242 34750
rect 7982 34802 8034 34814
rect 7982 34738 8034 34750
rect 8318 34802 8370 34814
rect 14478 34802 14530 34814
rect 8418 34750 8430 34802
rect 8482 34750 8494 34802
rect 10322 34750 10334 34802
rect 10386 34750 10398 34802
rect 8318 34738 8370 34750
rect 14478 34738 14530 34750
rect 19182 34802 19234 34814
rect 29710 34802 29762 34814
rect 25666 34750 25678 34802
rect 25730 34750 25742 34802
rect 30385 34799 30431 34974
rect 37998 34962 38050 34974
rect 40798 35026 40850 35038
rect 47518 35026 47570 35038
rect 42018 34974 42030 35026
rect 42082 34974 42094 35026
rect 45602 34974 45614 35026
rect 45666 34974 45678 35026
rect 40798 34962 40850 34974
rect 47518 34962 47570 34974
rect 50542 35026 50594 35038
rect 54462 35026 54514 35038
rect 57374 35026 57426 35038
rect 51762 34974 51774 35026
rect 51826 34974 51838 35026
rect 56466 34974 56478 35026
rect 56530 34974 56542 35026
rect 50542 34962 50594 34974
rect 54462 34962 54514 34974
rect 57374 34962 57426 34974
rect 31054 34914 31106 34926
rect 30818 34862 30830 34914
rect 30882 34862 30894 34914
rect 31054 34850 31106 34862
rect 31166 34914 31218 34926
rect 31166 34850 31218 34862
rect 32174 34914 32226 34926
rect 32174 34850 32226 34862
rect 32398 34914 32450 34926
rect 32398 34850 32450 34862
rect 32846 34914 32898 34926
rect 32846 34850 32898 34862
rect 33182 34914 33234 34926
rect 33182 34850 33234 34862
rect 34526 34914 34578 34926
rect 35870 34914 35922 34926
rect 34962 34862 34974 34914
rect 35026 34862 35038 34914
rect 34526 34850 34578 34862
rect 35870 34850 35922 34862
rect 37550 34914 37602 34926
rect 37550 34850 37602 34862
rect 37886 34914 37938 34926
rect 37886 34850 37938 34862
rect 38222 34914 38274 34926
rect 38222 34850 38274 34862
rect 42590 34914 42642 34926
rect 42590 34850 42642 34862
rect 43262 34914 43314 34926
rect 43262 34850 43314 34862
rect 43598 34914 43650 34926
rect 43598 34850 43650 34862
rect 43934 34914 43986 34926
rect 46958 34914 47010 34926
rect 52558 34914 52610 34926
rect 45826 34862 45838 34914
rect 45890 34862 45902 34914
rect 49074 34862 49086 34914
rect 49138 34862 49150 34914
rect 49858 34862 49870 34914
rect 49922 34862 49934 34914
rect 51650 34862 51662 34914
rect 51714 34862 51726 34914
rect 43934 34850 43986 34862
rect 46958 34850 47010 34862
rect 52558 34850 52610 34862
rect 53566 34914 53618 34926
rect 53778 34862 53790 34914
rect 53842 34862 53854 34914
rect 56690 34862 56702 34914
rect 56754 34862 56766 34914
rect 53566 34850 53618 34862
rect 33518 34802 33570 34814
rect 36094 34802 36146 34814
rect 30706 34799 30718 34802
rect 30385 34753 30718 34799
rect 30706 34750 30718 34753
rect 30770 34750 30782 34802
rect 35074 34750 35086 34802
rect 35138 34750 35150 34802
rect 19182 34738 19234 34750
rect 29710 34738 29762 34750
rect 33518 34738 33570 34750
rect 36094 34738 36146 34750
rect 36206 34802 36258 34814
rect 36206 34738 36258 34750
rect 38782 34802 38834 34814
rect 38782 34738 38834 34750
rect 39006 34802 39058 34814
rect 39006 34738 39058 34750
rect 42702 34802 42754 34814
rect 42702 34738 42754 34750
rect 46510 34802 46562 34814
rect 48962 34750 48974 34802
rect 49026 34750 49038 34802
rect 46510 34738 46562 34750
rect 2830 34690 2882 34702
rect 2830 34626 2882 34638
rect 5070 34690 5122 34702
rect 5070 34626 5122 34638
rect 5966 34690 6018 34702
rect 5966 34626 6018 34638
rect 6078 34690 6130 34702
rect 6078 34626 6130 34638
rect 6974 34690 7026 34702
rect 6974 34626 7026 34638
rect 7198 34690 7250 34702
rect 7198 34626 7250 34638
rect 8094 34690 8146 34702
rect 8094 34626 8146 34638
rect 8206 34690 8258 34702
rect 12350 34690 12402 34702
rect 11106 34638 11118 34690
rect 11170 34638 11182 34690
rect 8206 34626 8258 34638
rect 12350 34626 12402 34638
rect 12462 34690 12514 34702
rect 12462 34626 12514 34638
rect 12574 34690 12626 34702
rect 12574 34626 12626 34638
rect 15150 34690 15202 34702
rect 15150 34626 15202 34638
rect 16718 34690 16770 34702
rect 16718 34626 16770 34638
rect 17950 34690 18002 34702
rect 17950 34626 18002 34638
rect 19070 34690 19122 34702
rect 19070 34626 19122 34638
rect 19406 34690 19458 34702
rect 19406 34626 19458 34638
rect 21982 34690 22034 34702
rect 21982 34626 22034 34638
rect 23102 34690 23154 34702
rect 23102 34626 23154 34638
rect 23550 34690 23602 34702
rect 23550 34626 23602 34638
rect 26350 34690 26402 34702
rect 29934 34690 29986 34702
rect 32286 34690 32338 34702
rect 28578 34638 28590 34690
rect 28642 34638 28654 34690
rect 31602 34638 31614 34690
rect 31666 34638 31678 34690
rect 26350 34626 26402 34638
rect 29934 34626 29986 34638
rect 32286 34626 32338 34638
rect 33406 34690 33458 34702
rect 33406 34626 33458 34638
rect 34190 34690 34242 34702
rect 34190 34626 34242 34638
rect 36766 34690 36818 34702
rect 36766 34626 36818 34638
rect 38894 34690 38946 34702
rect 38894 34626 38946 34638
rect 39566 34690 39618 34702
rect 39566 34626 39618 34638
rect 39902 34690 39954 34702
rect 39902 34626 39954 34638
rect 40462 34690 40514 34702
rect 40462 34626 40514 34638
rect 41918 34690 41970 34702
rect 41918 34626 41970 34638
rect 42814 34690 42866 34702
rect 42814 34626 42866 34638
rect 43822 34690 43874 34702
rect 43822 34626 43874 34638
rect 44382 34690 44434 34702
rect 44382 34626 44434 34638
rect 47406 34690 47458 34702
rect 47406 34626 47458 34638
rect 47630 34690 47682 34702
rect 47630 34626 47682 34638
rect 1344 34522 59024 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 59024 34522
rect 1344 34436 59024 34470
rect 4174 34354 4226 34366
rect 4174 34290 4226 34302
rect 4510 34354 4562 34366
rect 4510 34290 4562 34302
rect 5406 34354 5458 34366
rect 5406 34290 5458 34302
rect 8542 34354 8594 34366
rect 8542 34290 8594 34302
rect 11902 34354 11954 34366
rect 11902 34290 11954 34302
rect 12238 34354 12290 34366
rect 12238 34290 12290 34302
rect 19182 34354 19234 34366
rect 19182 34290 19234 34302
rect 23550 34354 23602 34366
rect 23550 34290 23602 34302
rect 23998 34354 24050 34366
rect 23998 34290 24050 34302
rect 24446 34354 24498 34366
rect 24446 34290 24498 34302
rect 26014 34354 26066 34366
rect 26014 34290 26066 34302
rect 29822 34354 29874 34366
rect 29822 34290 29874 34302
rect 30606 34354 30658 34366
rect 30606 34290 30658 34302
rect 36654 34354 36706 34366
rect 36654 34290 36706 34302
rect 44942 34354 44994 34366
rect 44942 34290 44994 34302
rect 51214 34354 51266 34366
rect 51214 34290 51266 34302
rect 52110 34354 52162 34366
rect 52110 34290 52162 34302
rect 52334 34354 52386 34366
rect 52334 34290 52386 34302
rect 52670 34354 52722 34366
rect 56366 34354 56418 34366
rect 54002 34302 54014 34354
rect 54066 34302 54078 34354
rect 52670 34290 52722 34302
rect 56366 34290 56418 34302
rect 2942 34242 2994 34254
rect 2942 34178 2994 34190
rect 5294 34242 5346 34254
rect 5294 34178 5346 34190
rect 5966 34242 6018 34254
rect 8206 34242 8258 34254
rect 14142 34242 14194 34254
rect 7298 34190 7310 34242
rect 7362 34190 7374 34242
rect 7522 34190 7534 34242
rect 7586 34190 7598 34242
rect 12786 34190 12798 34242
rect 12850 34190 12862 34242
rect 5966 34178 6018 34190
rect 8206 34178 8258 34190
rect 14142 34178 14194 34190
rect 15598 34242 15650 34254
rect 15598 34178 15650 34190
rect 17838 34242 17890 34254
rect 17838 34178 17890 34190
rect 17950 34242 18002 34254
rect 17950 34178 18002 34190
rect 26462 34242 26514 34254
rect 26462 34178 26514 34190
rect 35310 34242 35362 34254
rect 40798 34242 40850 34254
rect 46958 34242 47010 34254
rect 39218 34190 39230 34242
rect 39282 34190 39294 34242
rect 39890 34190 39902 34242
rect 39954 34190 39966 34242
rect 42578 34190 42590 34242
rect 42642 34190 42654 34242
rect 35310 34178 35362 34190
rect 40798 34178 40850 34190
rect 46958 34178 47010 34190
rect 49534 34242 49586 34254
rect 49534 34178 49586 34190
rect 51998 34242 52050 34254
rect 51998 34178 52050 34190
rect 57486 34242 57538 34254
rect 57486 34178 57538 34190
rect 3502 34130 3554 34142
rect 3502 34066 3554 34078
rect 4062 34130 4114 34142
rect 4062 34066 4114 34078
rect 4286 34130 4338 34142
rect 4286 34066 4338 34078
rect 6414 34130 6466 34142
rect 6414 34066 6466 34078
rect 8094 34130 8146 34142
rect 14366 34130 14418 34142
rect 15822 34130 15874 34142
rect 10098 34078 10110 34130
rect 10162 34078 10174 34130
rect 10770 34078 10782 34130
rect 10834 34078 10846 34130
rect 13010 34078 13022 34130
rect 13074 34078 13086 34130
rect 13682 34078 13694 34130
rect 13746 34078 13758 34130
rect 14802 34078 14814 34130
rect 14866 34078 14878 34130
rect 8094 34066 8146 34078
rect 14366 34066 14418 34078
rect 15822 34066 15874 34078
rect 16046 34130 16098 34142
rect 16046 34066 16098 34078
rect 16158 34130 16210 34142
rect 16158 34066 16210 34078
rect 17614 34130 17666 34142
rect 17614 34066 17666 34078
rect 21086 34130 21138 34142
rect 21086 34066 21138 34078
rect 21534 34130 21586 34142
rect 21534 34066 21586 34078
rect 21646 34130 21698 34142
rect 21646 34066 21698 34078
rect 28590 34130 28642 34142
rect 34414 34130 34466 34142
rect 35758 34130 35810 34142
rect 41470 34130 41522 34142
rect 53454 34130 53506 34142
rect 31714 34078 31726 34130
rect 31778 34078 31790 34130
rect 31938 34078 31950 34130
rect 32002 34078 32014 34130
rect 34626 34078 34638 34130
rect 34690 34078 34702 34130
rect 38098 34078 38110 34130
rect 38162 34078 38174 34130
rect 39442 34078 39454 34130
rect 39506 34078 39518 34130
rect 40002 34078 40014 34130
rect 40066 34078 40078 34130
rect 43922 34078 43934 34130
rect 43986 34078 43998 34130
rect 46050 34078 46062 34130
rect 46114 34078 46126 34130
rect 47842 34078 47854 34130
rect 47906 34078 47918 34130
rect 49746 34078 49758 34130
rect 49810 34078 49822 34130
rect 49970 34078 49982 34130
rect 50034 34078 50046 34130
rect 28590 34066 28642 34078
rect 34414 34066 34466 34078
rect 35758 34066 35810 34078
rect 41470 34066 41522 34078
rect 53454 34066 53506 34078
rect 53678 34130 53730 34142
rect 53678 34066 53730 34078
rect 55918 34130 55970 34142
rect 55918 34066 55970 34078
rect 56142 34130 56194 34142
rect 56142 34066 56194 34078
rect 56478 34130 56530 34142
rect 57922 34078 57934 34130
rect 57986 34078 57998 34130
rect 56478 34066 56530 34078
rect 1934 34018 1986 34030
rect 1934 33954 1986 33966
rect 2494 34018 2546 34030
rect 2494 33954 2546 33966
rect 8990 34018 9042 34030
rect 15934 34018 15986 34030
rect 10546 33966 10558 34018
rect 10610 33966 10622 34018
rect 8990 33954 9042 33966
rect 15934 33954 15986 33966
rect 16942 34018 16994 34030
rect 16942 33954 16994 33966
rect 18734 34018 18786 34030
rect 18734 33954 18786 33966
rect 19742 34018 19794 34030
rect 19742 33954 19794 33966
rect 20190 34018 20242 34030
rect 20190 33954 20242 33966
rect 20638 34018 20690 34030
rect 20638 33954 20690 33966
rect 21310 34018 21362 34030
rect 21310 33954 21362 33966
rect 22318 34018 22370 34030
rect 22318 33954 22370 33966
rect 22654 34018 22706 34030
rect 22654 33954 22706 33966
rect 23102 34018 23154 34030
rect 23102 33954 23154 33966
rect 24894 34018 24946 34030
rect 24894 33954 24946 33966
rect 25566 34018 25618 34030
rect 33518 34018 33570 34030
rect 28018 33966 28030 34018
rect 28082 33966 28094 34018
rect 29026 33966 29038 34018
rect 29090 33966 29102 34018
rect 32050 33966 32062 34018
rect 32114 33966 32126 34018
rect 25566 33954 25618 33966
rect 33518 33954 33570 33966
rect 36206 34018 36258 34030
rect 36206 33954 36258 33966
rect 37102 34018 37154 34030
rect 37102 33954 37154 33966
rect 37550 34018 37602 34030
rect 44494 34018 44546 34030
rect 48526 34018 48578 34030
rect 40226 33966 40238 34018
rect 40290 33966 40302 34018
rect 42354 33966 42366 34018
rect 42418 33966 42430 34018
rect 46498 33966 46510 34018
rect 46562 33966 46574 34018
rect 47618 33966 47630 34018
rect 47682 33966 47694 34018
rect 58258 33966 58270 34018
rect 58322 33966 58334 34018
rect 37550 33954 37602 33966
rect 44494 33954 44546 33966
rect 48526 33954 48578 33966
rect 5518 33906 5570 33918
rect 27134 33906 27186 33918
rect 5730 33854 5742 33906
rect 5794 33903 5806 33906
rect 6178 33903 6190 33906
rect 5794 33857 6190 33903
rect 5794 33854 5806 33857
rect 6178 33854 6190 33857
rect 6242 33854 6254 33906
rect 10098 33854 10110 33906
rect 10162 33854 10174 33906
rect 22306 33854 22318 33906
rect 22370 33903 22382 33906
rect 22530 33903 22542 33906
rect 22370 33857 22542 33903
rect 22370 33854 22382 33857
rect 22530 33854 22542 33857
rect 22594 33903 22606 33906
rect 23314 33903 23326 33906
rect 22594 33857 23326 33903
rect 22594 33854 22606 33857
rect 23314 33854 23326 33857
rect 23378 33854 23390 33906
rect 23650 33854 23662 33906
rect 23714 33903 23726 33906
rect 24546 33903 24558 33906
rect 23714 33857 24558 33903
rect 23714 33854 23726 33857
rect 24546 33854 24558 33857
rect 24610 33854 24622 33906
rect 5518 33842 5570 33854
rect 27134 33842 27186 33854
rect 27246 33906 27298 33918
rect 27246 33842 27298 33854
rect 27470 33906 27522 33918
rect 27470 33842 27522 33854
rect 30382 33906 30434 33918
rect 30382 33842 30434 33854
rect 30718 33906 30770 33918
rect 32498 33854 32510 33906
rect 32562 33854 32574 33906
rect 30718 33842 30770 33854
rect 1344 33738 59024 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 59024 33738
rect 1344 33652 59024 33686
rect 9886 33570 9938 33582
rect 9886 33506 9938 33518
rect 10782 33570 10834 33582
rect 39118 33570 39170 33582
rect 34738 33518 34750 33570
rect 34802 33567 34814 33570
rect 35186 33567 35198 33570
rect 34802 33521 35198 33567
rect 34802 33518 34814 33521
rect 35186 33518 35198 33521
rect 35250 33518 35262 33570
rect 42466 33518 42478 33570
rect 42530 33567 42542 33570
rect 43362 33567 43374 33570
rect 42530 33521 43374 33567
rect 42530 33518 42542 33521
rect 43362 33518 43374 33521
rect 43426 33518 43438 33570
rect 48962 33518 48974 33570
rect 49026 33567 49038 33570
rect 49522 33567 49534 33570
rect 49026 33521 49534 33567
rect 49026 33518 49038 33521
rect 49522 33518 49534 33521
rect 49586 33518 49598 33570
rect 10782 33506 10834 33518
rect 39118 33506 39170 33518
rect 12910 33458 12962 33470
rect 16046 33458 16098 33470
rect 2258 33406 2270 33458
rect 2322 33406 2334 33458
rect 6066 33406 6078 33458
rect 6130 33406 6142 33458
rect 6626 33406 6638 33458
rect 6690 33406 6702 33458
rect 8082 33406 8094 33458
rect 8146 33406 8158 33458
rect 14242 33406 14254 33458
rect 14306 33406 14318 33458
rect 14802 33406 14814 33458
rect 14866 33406 14878 33458
rect 12910 33394 12962 33406
rect 16046 33394 16098 33406
rect 19630 33458 19682 33470
rect 19630 33394 19682 33406
rect 20414 33458 20466 33470
rect 26798 33458 26850 33470
rect 29822 33458 29874 33470
rect 22418 33406 22430 33458
rect 22482 33406 22494 33458
rect 27682 33406 27694 33458
rect 27746 33406 27758 33458
rect 20414 33394 20466 33406
rect 26798 33394 26850 33406
rect 29822 33394 29874 33406
rect 32958 33458 33010 33470
rect 32958 33394 33010 33406
rect 34302 33458 34354 33470
rect 34302 33394 34354 33406
rect 35198 33458 35250 33470
rect 35198 33394 35250 33406
rect 42478 33458 42530 33470
rect 42478 33394 42530 33406
rect 43374 33458 43426 33470
rect 43374 33394 43426 33406
rect 45502 33458 45554 33470
rect 57934 33458 57986 33470
rect 56466 33406 56478 33458
rect 56530 33406 56542 33458
rect 45502 33394 45554 33406
rect 57934 33394 57986 33406
rect 9998 33346 10050 33358
rect 15822 33346 15874 33358
rect 3378 33294 3390 33346
rect 3442 33294 3454 33346
rect 5618 33294 5630 33346
rect 5682 33294 5694 33346
rect 6402 33294 6414 33346
rect 6466 33294 6478 33346
rect 14354 33294 14366 33346
rect 14418 33294 14430 33346
rect 15026 33294 15038 33346
rect 15090 33294 15102 33346
rect 9998 33282 10050 33294
rect 15822 33282 15874 33294
rect 16270 33346 16322 33358
rect 16270 33282 16322 33294
rect 17838 33346 17890 33358
rect 17838 33282 17890 33294
rect 17950 33346 18002 33358
rect 17950 33282 18002 33294
rect 18398 33346 18450 33358
rect 18398 33282 18450 33294
rect 18846 33346 18898 33358
rect 18846 33282 18898 33294
rect 18958 33346 19010 33358
rect 21646 33346 21698 33358
rect 19954 33294 19966 33346
rect 20018 33294 20030 33346
rect 18958 33282 19010 33294
rect 21646 33282 21698 33294
rect 22878 33346 22930 33358
rect 22878 33282 22930 33294
rect 23214 33346 23266 33358
rect 37438 33346 37490 33358
rect 41246 33346 41298 33358
rect 24210 33294 24222 33346
rect 24274 33294 24286 33346
rect 24546 33294 24558 33346
rect 24610 33294 24622 33346
rect 27570 33294 27582 33346
rect 27634 33294 27646 33346
rect 28466 33294 28478 33346
rect 28530 33294 28542 33346
rect 31154 33294 31166 33346
rect 31218 33294 31230 33346
rect 32050 33294 32062 33346
rect 32114 33294 32126 33346
rect 35970 33294 35982 33346
rect 36034 33294 36046 33346
rect 38434 33294 38446 33346
rect 38498 33294 38510 33346
rect 23214 33282 23266 33294
rect 37438 33282 37490 33294
rect 41246 33282 41298 33294
rect 46398 33346 46450 33358
rect 46398 33282 46450 33294
rect 46734 33346 46786 33358
rect 58046 33346 58098 33358
rect 56242 33294 56254 33346
rect 56306 33294 56318 33346
rect 57474 33294 57486 33346
rect 57538 33294 57550 33346
rect 46734 33282 46786 33294
rect 58046 33282 58098 33294
rect 17614 33234 17666 33246
rect 4274 33182 4286 33234
rect 4338 33182 4350 33234
rect 11778 33182 11790 33234
rect 11842 33182 11854 33234
rect 17378 33182 17390 33234
rect 17442 33182 17454 33234
rect 17614 33170 17666 33182
rect 18622 33234 18674 33246
rect 18622 33170 18674 33182
rect 21982 33234 22034 33246
rect 32510 33234 32562 33246
rect 22082 33182 22094 33234
rect 22146 33182 22158 33234
rect 25778 33182 25790 33234
rect 25842 33182 25854 33234
rect 27906 33182 27918 33234
rect 27970 33182 27982 33234
rect 30706 33182 30718 33234
rect 30770 33182 30782 33234
rect 21982 33170 22034 33182
rect 32510 33170 32562 33182
rect 34750 33234 34802 33246
rect 34750 33170 34802 33182
rect 36318 33234 36370 33246
rect 36318 33170 36370 33182
rect 40014 33234 40066 33246
rect 40014 33170 40066 33182
rect 40910 33234 40962 33246
rect 40910 33170 40962 33182
rect 56926 33234 56978 33246
rect 56926 33170 56978 33182
rect 2830 33122 2882 33134
rect 2830 33058 2882 33070
rect 8542 33122 8594 33134
rect 8542 33058 8594 33070
rect 9214 33122 9266 33134
rect 9214 33058 9266 33070
rect 9886 33122 9938 33134
rect 9886 33058 9938 33070
rect 12462 33122 12514 33134
rect 12462 33058 12514 33070
rect 16382 33122 16434 33134
rect 16382 33058 16434 33070
rect 16494 33122 16546 33134
rect 16494 33058 16546 33070
rect 17726 33122 17778 33134
rect 17726 33058 17778 33070
rect 19742 33122 19794 33134
rect 19742 33058 19794 33070
rect 20862 33122 20914 33134
rect 20862 33058 20914 33070
rect 21870 33122 21922 33134
rect 21870 33058 21922 33070
rect 23102 33122 23154 33134
rect 23102 33058 23154 33070
rect 26350 33122 26402 33134
rect 26350 33058 26402 33070
rect 33406 33122 33458 33134
rect 33406 33058 33458 33070
rect 33854 33122 33906 33134
rect 33854 33058 33906 33070
rect 36430 33122 36482 33134
rect 36430 33058 36482 33070
rect 36542 33122 36594 33134
rect 36542 33058 36594 33070
rect 40126 33122 40178 33134
rect 40126 33058 40178 33070
rect 40238 33122 40290 33134
rect 40238 33058 40290 33070
rect 41022 33122 41074 33134
rect 41022 33058 41074 33070
rect 41582 33122 41634 33134
rect 41582 33058 41634 33070
rect 42030 33122 42082 33134
rect 42030 33058 42082 33070
rect 43038 33122 43090 33134
rect 43038 33058 43090 33070
rect 43822 33122 43874 33134
rect 43822 33058 43874 33070
rect 44382 33122 44434 33134
rect 44382 33058 44434 33070
rect 46510 33122 46562 33134
rect 46510 33058 46562 33070
rect 47070 33122 47122 33134
rect 47070 33058 47122 33070
rect 48974 33122 49026 33134
rect 48974 33058 49026 33070
rect 49422 33122 49474 33134
rect 49422 33058 49474 33070
rect 54798 33122 54850 33134
rect 54798 33058 54850 33070
rect 57822 33122 57874 33134
rect 57822 33058 57874 33070
rect 1344 32954 59024 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 59024 32954
rect 1344 32868 59024 32902
rect 1934 32786 1986 32798
rect 1934 32722 1986 32734
rect 2382 32786 2434 32798
rect 2382 32722 2434 32734
rect 5518 32786 5570 32798
rect 5518 32722 5570 32734
rect 6414 32786 6466 32798
rect 6414 32722 6466 32734
rect 13806 32786 13858 32798
rect 13806 32722 13858 32734
rect 15822 32786 15874 32798
rect 15822 32722 15874 32734
rect 18398 32786 18450 32798
rect 18398 32722 18450 32734
rect 19406 32786 19458 32798
rect 19406 32722 19458 32734
rect 22990 32786 23042 32798
rect 22990 32722 23042 32734
rect 31502 32786 31554 32798
rect 31502 32722 31554 32734
rect 31726 32786 31778 32798
rect 31726 32722 31778 32734
rect 32398 32786 32450 32798
rect 32398 32722 32450 32734
rect 34526 32786 34578 32798
rect 34526 32722 34578 32734
rect 39118 32786 39170 32798
rect 39118 32722 39170 32734
rect 44046 32786 44098 32798
rect 44046 32722 44098 32734
rect 49870 32786 49922 32798
rect 49870 32722 49922 32734
rect 50878 32786 50930 32798
rect 50878 32722 50930 32734
rect 57486 32786 57538 32798
rect 57486 32722 57538 32734
rect 6078 32674 6130 32686
rect 4274 32622 4286 32674
rect 4338 32622 4350 32674
rect 6078 32610 6130 32622
rect 6190 32674 6242 32686
rect 6190 32610 6242 32622
rect 8542 32674 8594 32686
rect 13470 32674 13522 32686
rect 12114 32622 12126 32674
rect 12178 32622 12190 32674
rect 8542 32610 8594 32622
rect 13470 32610 13522 32622
rect 13582 32674 13634 32686
rect 13582 32610 13634 32622
rect 14366 32674 14418 32686
rect 14366 32610 14418 32622
rect 14590 32674 14642 32686
rect 14590 32610 14642 32622
rect 16382 32674 16434 32686
rect 22766 32674 22818 32686
rect 20290 32622 20302 32674
rect 20354 32622 20366 32674
rect 20738 32622 20750 32674
rect 20802 32622 20814 32674
rect 16382 32610 16434 32622
rect 22766 32610 22818 32622
rect 23326 32674 23378 32686
rect 31838 32674 31890 32686
rect 38334 32674 38386 32686
rect 25666 32622 25678 32674
rect 25730 32622 25742 32674
rect 30818 32622 30830 32674
rect 30882 32622 30894 32674
rect 35410 32622 35422 32674
rect 35474 32622 35486 32674
rect 23326 32610 23378 32622
rect 31838 32610 31890 32622
rect 38334 32610 38386 32622
rect 44830 32674 44882 32686
rect 44830 32610 44882 32622
rect 44942 32674 44994 32686
rect 44942 32610 44994 32622
rect 54462 32674 54514 32686
rect 54462 32610 54514 32622
rect 56030 32674 56082 32686
rect 56030 32610 56082 32622
rect 57710 32674 57762 32686
rect 57710 32610 57762 32622
rect 7646 32562 7698 32574
rect 4498 32510 4510 32562
rect 4562 32510 4574 32562
rect 5058 32510 5070 32562
rect 5122 32510 5134 32562
rect 7410 32510 7422 32562
rect 7474 32510 7486 32562
rect 7646 32498 7698 32510
rect 9102 32562 9154 32574
rect 14254 32562 14306 32574
rect 10210 32510 10222 32562
rect 10274 32510 10286 32562
rect 11218 32510 11230 32562
rect 11282 32510 11294 32562
rect 11666 32510 11678 32562
rect 11730 32510 11742 32562
rect 12562 32510 12574 32562
rect 12626 32510 12638 32562
rect 9102 32498 9154 32510
rect 14254 32498 14306 32510
rect 14702 32562 14754 32574
rect 14702 32498 14754 32510
rect 16718 32562 16770 32574
rect 18622 32562 18674 32574
rect 23214 32562 23266 32574
rect 16930 32510 16942 32562
rect 16994 32510 17006 32562
rect 20178 32510 20190 32562
rect 20242 32510 20254 32562
rect 21074 32510 21086 32562
rect 21138 32510 21150 32562
rect 21746 32510 21758 32562
rect 21810 32510 21822 32562
rect 16718 32498 16770 32510
rect 18622 32498 18674 32510
rect 23214 32498 23266 32510
rect 24334 32562 24386 32574
rect 28142 32562 28194 32574
rect 34414 32562 34466 32574
rect 26002 32510 26014 32562
rect 26066 32510 26078 32562
rect 26898 32510 26910 32562
rect 26962 32510 26974 32562
rect 28690 32510 28702 32562
rect 28754 32510 28766 32562
rect 29922 32510 29934 32562
rect 29986 32510 29998 32562
rect 30482 32510 30494 32562
rect 30546 32510 30558 32562
rect 24334 32498 24386 32510
rect 28142 32498 28194 32510
rect 34414 32498 34466 32510
rect 34750 32562 34802 32574
rect 36990 32562 37042 32574
rect 35298 32510 35310 32562
rect 35362 32510 35374 32562
rect 34750 32498 34802 32510
rect 36990 32498 37042 32510
rect 38222 32562 38274 32574
rect 38222 32498 38274 32510
rect 38558 32562 38610 32574
rect 38558 32498 38610 32510
rect 39230 32562 39282 32574
rect 39230 32498 39282 32510
rect 39902 32562 39954 32574
rect 41918 32562 41970 32574
rect 45166 32562 45218 32574
rect 40114 32510 40126 32562
rect 40178 32510 40190 32562
rect 42914 32510 42926 32562
rect 42978 32510 42990 32562
rect 39902 32498 39954 32510
rect 41918 32498 41970 32510
rect 45166 32498 45218 32510
rect 50430 32562 50482 32574
rect 50430 32498 50482 32510
rect 50766 32562 50818 32574
rect 50766 32498 50818 32510
rect 50990 32562 51042 32574
rect 57822 32562 57874 32574
rect 53778 32510 53790 32562
rect 53842 32510 53854 32562
rect 55346 32510 55358 32562
rect 55410 32510 55422 32562
rect 50990 32498 51042 32510
rect 57822 32498 57874 32510
rect 2942 32450 2994 32462
rect 2942 32386 2994 32398
rect 3390 32450 3442 32462
rect 8094 32450 8146 32462
rect 4050 32398 4062 32450
rect 4114 32398 4126 32450
rect 3390 32386 3442 32398
rect 8094 32386 8146 32398
rect 9998 32450 10050 32462
rect 15374 32450 15426 32462
rect 12338 32398 12350 32450
rect 12402 32398 12414 32450
rect 9998 32386 10050 32398
rect 15374 32386 15426 32398
rect 16494 32450 16546 32462
rect 16494 32386 16546 32398
rect 17950 32450 18002 32462
rect 17950 32386 18002 32398
rect 18174 32450 18226 32462
rect 24110 32450 24162 32462
rect 18498 32398 18510 32450
rect 18562 32398 18574 32450
rect 19954 32398 19966 32450
rect 20018 32398 20030 32450
rect 23314 32398 23326 32450
rect 23378 32398 23390 32450
rect 18174 32386 18226 32398
rect 24110 32386 24162 32398
rect 25902 32450 25954 32462
rect 25902 32386 25954 32398
rect 27918 32450 27970 32462
rect 27918 32386 27970 32398
rect 32734 32450 32786 32462
rect 32734 32386 32786 32398
rect 33630 32450 33682 32462
rect 33630 32386 33682 32398
rect 37438 32450 37490 32462
rect 37438 32386 37490 32398
rect 40798 32450 40850 32462
rect 43598 32450 43650 32462
rect 42690 32398 42702 32450
rect 42754 32398 42766 32450
rect 40798 32386 40850 32398
rect 43598 32386 43650 32398
rect 45502 32450 45554 32462
rect 45502 32386 45554 32398
rect 51550 32450 51602 32462
rect 54002 32398 54014 32450
rect 54066 32398 54078 32450
rect 55122 32398 55134 32450
rect 55186 32398 55198 32450
rect 51550 32386 51602 32398
rect 17726 32338 17778 32350
rect 6962 32286 6974 32338
rect 7026 32286 7038 32338
rect 10098 32286 10110 32338
rect 10162 32286 10174 32338
rect 17726 32274 17778 32286
rect 24558 32338 24610 32350
rect 24558 32274 24610 32286
rect 25006 32338 25058 32350
rect 36094 32338 36146 32350
rect 27570 32286 27582 32338
rect 27634 32286 27646 32338
rect 25006 32274 25058 32286
rect 36094 32274 36146 32286
rect 36430 32338 36482 32350
rect 36430 32274 36482 32286
rect 39118 32338 39170 32350
rect 39118 32274 39170 32286
rect 42030 32338 42082 32350
rect 42030 32274 42082 32286
rect 1344 32170 59024 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 59024 32170
rect 1344 32084 59024 32118
rect 2034 31950 2046 32002
rect 2098 31999 2110 32002
rect 2482 31999 2494 32002
rect 2098 31953 2494 31999
rect 2098 31950 2110 31953
rect 2482 31950 2494 31953
rect 2546 31950 2558 32002
rect 18498 31950 18510 32002
rect 18562 31999 18574 32002
rect 19282 31999 19294 32002
rect 18562 31953 19294 31999
rect 18562 31950 18574 31953
rect 19282 31950 19294 31953
rect 19346 31950 19358 32002
rect 28130 31950 28142 32002
rect 28194 31999 28206 32002
rect 28466 31999 28478 32002
rect 28194 31953 28478 31999
rect 28194 31950 28206 31953
rect 28466 31950 28478 31953
rect 28530 31950 28542 32002
rect 58146 31950 58158 32002
rect 58210 31950 58222 32002
rect 2382 31890 2434 31902
rect 5070 31890 5122 31902
rect 3378 31838 3390 31890
rect 3442 31838 3454 31890
rect 2382 31826 2434 31838
rect 5070 31826 5122 31838
rect 5854 31890 5906 31902
rect 5854 31826 5906 31838
rect 6302 31890 6354 31902
rect 6302 31826 6354 31838
rect 12910 31890 12962 31902
rect 12910 31826 12962 31838
rect 16830 31890 16882 31902
rect 16830 31826 16882 31838
rect 17726 31890 17778 31902
rect 17726 31826 17778 31838
rect 18286 31890 18338 31902
rect 18286 31826 18338 31838
rect 19070 31890 19122 31902
rect 19070 31826 19122 31838
rect 20190 31890 20242 31902
rect 20190 31826 20242 31838
rect 22878 31890 22930 31902
rect 24446 31890 24498 31902
rect 23538 31838 23550 31890
rect 23602 31838 23614 31890
rect 22878 31826 22930 31838
rect 24446 31826 24498 31838
rect 25006 31890 25058 31902
rect 27918 31890 27970 31902
rect 26562 31838 26574 31890
rect 26626 31838 26638 31890
rect 25006 31826 25058 31838
rect 27918 31826 27970 31838
rect 34190 31890 34242 31902
rect 47070 31890 47122 31902
rect 53902 31890 53954 31902
rect 40002 31838 40014 31890
rect 40066 31838 40078 31890
rect 44370 31838 44382 31890
rect 44434 31838 44446 31890
rect 48290 31838 48302 31890
rect 48354 31838 48366 31890
rect 34190 31826 34242 31838
rect 47070 31826 47122 31838
rect 53902 31826 53954 31838
rect 54462 31890 54514 31902
rect 54462 31826 54514 31838
rect 55470 31890 55522 31902
rect 55794 31838 55806 31890
rect 55858 31838 55870 31890
rect 57698 31838 57710 31890
rect 57762 31838 57774 31890
rect 55470 31826 55522 31838
rect 7086 31778 7138 31790
rect 6738 31726 6750 31778
rect 6802 31726 6814 31778
rect 7086 31714 7138 31726
rect 7758 31778 7810 31790
rect 7758 31714 7810 31726
rect 7870 31778 7922 31790
rect 13582 31778 13634 31790
rect 15150 31778 15202 31790
rect 18734 31778 18786 31790
rect 9314 31726 9326 31778
rect 9378 31726 9390 31778
rect 11106 31726 11118 31778
rect 11170 31726 11182 31778
rect 13906 31726 13918 31778
rect 13970 31726 13982 31778
rect 15810 31726 15822 31778
rect 15874 31726 15886 31778
rect 7870 31714 7922 31726
rect 13582 31714 13634 31726
rect 15150 31714 15202 31726
rect 18734 31714 18786 31726
rect 19966 31778 20018 31790
rect 19966 31714 20018 31726
rect 20526 31778 20578 31790
rect 20526 31714 20578 31726
rect 21758 31778 21810 31790
rect 21758 31714 21810 31726
rect 21982 31778 22034 31790
rect 21982 31714 22034 31726
rect 22430 31778 22482 31790
rect 31838 31778 31890 31790
rect 34078 31778 34130 31790
rect 45390 31778 45442 31790
rect 23762 31726 23774 31778
rect 23826 31726 23838 31778
rect 25890 31726 25902 31778
rect 25954 31726 25966 31778
rect 26674 31726 26686 31778
rect 26738 31726 26750 31778
rect 29922 31726 29934 31778
rect 29986 31726 29998 31778
rect 32610 31726 32622 31778
rect 32674 31726 32686 31778
rect 34402 31726 34414 31778
rect 34466 31726 34478 31778
rect 36418 31726 36430 31778
rect 36482 31726 36494 31778
rect 39218 31726 39230 31778
rect 39282 31726 39294 31778
rect 41682 31726 41694 31778
rect 41746 31726 41758 31778
rect 42242 31726 42254 31778
rect 42306 31726 42318 31778
rect 43810 31726 43822 31778
rect 43874 31726 43886 31778
rect 22430 31714 22482 31726
rect 31838 31714 31890 31726
rect 34078 31714 34130 31726
rect 45390 31714 45442 31726
rect 46062 31778 46114 31790
rect 49758 31778 49810 31790
rect 52446 31778 52498 31790
rect 48402 31726 48414 31778
rect 48466 31726 48478 31778
rect 49970 31726 49982 31778
rect 50034 31726 50046 31778
rect 51762 31726 51774 31778
rect 51826 31726 51838 31778
rect 46062 31714 46114 31726
rect 49758 31714 49810 31726
rect 52446 31714 52498 31726
rect 53342 31778 53394 31790
rect 53342 31714 53394 31726
rect 55246 31778 55298 31790
rect 57586 31726 57598 31778
rect 57650 31726 57662 31778
rect 55246 31714 55298 31726
rect 2830 31666 2882 31678
rect 2830 31602 2882 31614
rect 8654 31666 8706 31678
rect 14142 31666 14194 31678
rect 9202 31614 9214 31666
rect 9266 31614 9278 31666
rect 11442 31614 11454 31666
rect 11506 31614 11518 31666
rect 8654 31602 8706 31614
rect 14142 31602 14194 31614
rect 14590 31666 14642 31678
rect 15486 31666 15538 31678
rect 15250 31614 15262 31666
rect 15314 31614 15326 31666
rect 14590 31602 14642 31614
rect 15486 31602 15538 31614
rect 20414 31666 20466 31678
rect 31726 31666 31778 31678
rect 37774 31666 37826 31678
rect 42814 31666 42866 31678
rect 27346 31614 27358 31666
rect 27410 31614 27422 31666
rect 29586 31614 29598 31666
rect 29650 31614 29662 31666
rect 35858 31614 35870 31666
rect 35922 31614 35934 31666
rect 38882 31614 38894 31666
rect 38946 31614 38958 31666
rect 20414 31602 20466 31614
rect 31726 31602 31778 31614
rect 37774 31602 37826 31614
rect 42814 31602 42866 31614
rect 44718 31666 44770 31678
rect 44718 31602 44770 31614
rect 45838 31666 45890 31678
rect 45838 31602 45890 31614
rect 49086 31666 49138 31678
rect 49086 31602 49138 31614
rect 50654 31666 50706 31678
rect 50654 31602 50706 31614
rect 52670 31666 52722 31678
rect 52670 31602 52722 31614
rect 54014 31666 54066 31678
rect 54014 31602 54066 31614
rect 1934 31554 1986 31566
rect 1934 31490 1986 31502
rect 3838 31554 3890 31566
rect 3838 31490 3890 31502
rect 4622 31554 4674 31566
rect 4622 31490 4674 31502
rect 7646 31554 7698 31566
rect 7646 31490 7698 31502
rect 8094 31554 8146 31566
rect 8094 31490 8146 31502
rect 12014 31554 12066 31566
rect 12014 31490 12066 31502
rect 12462 31554 12514 31566
rect 12462 31490 12514 31502
rect 14254 31554 14306 31566
rect 14254 31490 14306 31502
rect 16158 31554 16210 31566
rect 16158 31490 16210 31502
rect 17278 31554 17330 31566
rect 17278 31490 17330 31502
rect 19518 31554 19570 31566
rect 19518 31490 19570 31502
rect 22206 31554 22258 31566
rect 22206 31490 22258 31502
rect 25566 31554 25618 31566
rect 25566 31490 25618 31502
rect 28366 31554 28418 31566
rect 28366 31490 28418 31502
rect 28814 31554 28866 31566
rect 30718 31554 30770 31566
rect 30146 31502 30158 31554
rect 30210 31502 30222 31554
rect 28814 31490 28866 31502
rect 30718 31490 30770 31502
rect 31166 31554 31218 31566
rect 31166 31490 31218 31502
rect 31950 31554 32002 31566
rect 31950 31490 32002 31502
rect 37438 31554 37490 31566
rect 37438 31490 37490 31502
rect 37662 31554 37714 31566
rect 37662 31490 37714 31502
rect 42926 31554 42978 31566
rect 42926 31490 42978 31502
rect 43150 31554 43202 31566
rect 43150 31490 43202 31502
rect 45950 31554 46002 31566
rect 45950 31490 46002 31502
rect 47518 31554 47570 31566
rect 47518 31490 47570 31502
rect 53790 31554 53842 31566
rect 53790 31490 53842 31502
rect 1344 31386 59024 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 59024 31386
rect 1344 31300 59024 31334
rect 2382 31218 2434 31230
rect 2382 31154 2434 31166
rect 2718 31218 2770 31230
rect 2718 31154 2770 31166
rect 12126 31218 12178 31230
rect 12126 31154 12178 31166
rect 12686 31218 12738 31230
rect 12686 31154 12738 31166
rect 13134 31218 13186 31230
rect 13134 31154 13186 31166
rect 13694 31218 13746 31230
rect 13694 31154 13746 31166
rect 17054 31218 17106 31230
rect 17054 31154 17106 31166
rect 17838 31218 17890 31230
rect 17838 31154 17890 31166
rect 18846 31218 18898 31230
rect 18846 31154 18898 31166
rect 21422 31218 21474 31230
rect 21422 31154 21474 31166
rect 21646 31218 21698 31230
rect 21646 31154 21698 31166
rect 23998 31218 24050 31230
rect 23998 31154 24050 31166
rect 25006 31218 25058 31230
rect 35982 31218 36034 31230
rect 35298 31166 35310 31218
rect 35362 31166 35374 31218
rect 25006 31154 25058 31166
rect 35982 31154 36034 31166
rect 38110 31218 38162 31230
rect 38110 31154 38162 31166
rect 40574 31218 40626 31230
rect 40574 31154 40626 31166
rect 43822 31218 43874 31230
rect 43822 31154 43874 31166
rect 44270 31218 44322 31230
rect 44270 31154 44322 31166
rect 44718 31218 44770 31230
rect 44718 31154 44770 31166
rect 47182 31218 47234 31230
rect 47182 31154 47234 31166
rect 47630 31218 47682 31230
rect 52782 31218 52834 31230
rect 48738 31166 48750 31218
rect 48802 31166 48814 31218
rect 47630 31154 47682 31166
rect 52782 31154 52834 31166
rect 54798 31218 54850 31230
rect 54798 31154 54850 31166
rect 55246 31218 55298 31230
rect 55246 31154 55298 31166
rect 16494 31106 16546 31118
rect 21870 31106 21922 31118
rect 32622 31106 32674 31118
rect 7186 31054 7198 31106
rect 7250 31054 7262 31106
rect 19394 31054 19406 31106
rect 19458 31054 19470 31106
rect 29362 31054 29374 31106
rect 29426 31054 29438 31106
rect 16494 31042 16546 31054
rect 21870 31042 21922 31054
rect 32622 31042 32674 31054
rect 32734 31106 32786 31118
rect 39118 31106 39170 31118
rect 33730 31054 33742 31106
rect 33794 31054 33806 31106
rect 35634 31054 35646 31106
rect 35698 31054 35710 31106
rect 32734 31042 32786 31054
rect 39118 31042 39170 31054
rect 39790 31106 39842 31118
rect 39790 31042 39842 31054
rect 40014 31106 40066 31118
rect 40014 31042 40066 31054
rect 42702 31106 42754 31118
rect 42702 31042 42754 31054
rect 48190 31106 48242 31118
rect 48190 31042 48242 31054
rect 49534 31106 49586 31118
rect 49534 31042 49586 31054
rect 49758 31106 49810 31118
rect 49758 31042 49810 31054
rect 51550 31106 51602 31118
rect 51550 31042 51602 31054
rect 52446 31106 52498 31118
rect 52446 31042 52498 31054
rect 52558 31106 52610 31118
rect 52558 31042 52610 31054
rect 8542 30994 8594 31006
rect 3714 30942 3726 30994
rect 3778 30942 3790 30994
rect 4834 30942 4846 30994
rect 4898 30942 4910 30994
rect 5170 30942 5182 30994
rect 5234 30942 5246 30994
rect 6626 30942 6638 30994
rect 6690 30942 6702 30994
rect 7074 30942 7086 30994
rect 7138 30942 7150 30994
rect 8542 30930 8594 30942
rect 8766 30994 8818 31006
rect 8766 30930 8818 30942
rect 8990 30994 9042 31006
rect 8990 30930 9042 30942
rect 9662 30994 9714 31006
rect 9662 30930 9714 30942
rect 10110 30994 10162 31006
rect 10110 30930 10162 30942
rect 10334 30994 10386 31006
rect 10334 30930 10386 30942
rect 10782 30994 10834 31006
rect 10782 30930 10834 30942
rect 11230 30994 11282 31006
rect 11230 30930 11282 30942
rect 11454 30994 11506 31006
rect 15150 30994 15202 31006
rect 13794 30942 13806 30994
rect 13858 30942 13870 30994
rect 11454 30930 11506 30942
rect 15150 30930 15202 30942
rect 15374 30994 15426 31006
rect 25902 30994 25954 31006
rect 19282 30942 19294 30994
rect 19346 30942 19358 30994
rect 20290 30942 20302 30994
rect 20354 30942 20366 30994
rect 15374 30930 15426 30942
rect 25902 30930 25954 30942
rect 26126 30994 26178 31006
rect 26126 30930 26178 30942
rect 27582 30994 27634 31006
rect 31838 30994 31890 31006
rect 36766 30994 36818 31006
rect 43150 30994 43202 31006
rect 28466 30942 28478 30994
rect 28530 30942 28542 30994
rect 34178 30942 34190 30994
rect 34242 30942 34254 30994
rect 34626 30942 34638 30994
rect 34690 30942 34702 30994
rect 34962 30942 34974 30994
rect 35026 30942 35038 30994
rect 36978 30942 36990 30994
rect 37042 30942 37054 30994
rect 41794 30942 41806 30994
rect 41858 30942 41870 30994
rect 27582 30930 27634 30942
rect 31838 30930 31890 30942
rect 36766 30930 36818 30942
rect 43150 30930 43202 30942
rect 43598 30994 43650 31006
rect 45826 30942 45838 30994
rect 45890 30942 45902 30994
rect 50866 30942 50878 30994
rect 50930 30942 50942 30994
rect 43598 30930 43650 30942
rect 1934 30882 1986 30894
rect 8878 30882 8930 30894
rect 7298 30830 7310 30882
rect 7362 30830 7374 30882
rect 1934 30818 1986 30830
rect 8878 30818 8930 30830
rect 10222 30882 10274 30894
rect 10222 30818 10274 30830
rect 11006 30882 11058 30894
rect 18286 30882 18338 30894
rect 20078 30882 20130 30894
rect 22654 30882 22706 30894
rect 13906 30830 13918 30882
rect 13970 30830 13982 30882
rect 19842 30830 19854 30882
rect 19906 30830 19918 30882
rect 21522 30830 21534 30882
rect 21586 30830 21598 30882
rect 11006 30818 11058 30830
rect 18286 30818 18338 30830
rect 20078 30818 20130 30830
rect 22654 30818 22706 30830
rect 23214 30882 23266 30894
rect 23214 30818 23266 30830
rect 23662 30882 23714 30894
rect 23662 30818 23714 30830
rect 24446 30882 24498 30894
rect 24446 30818 24498 30830
rect 25678 30882 25730 30894
rect 25678 30818 25730 30830
rect 30494 30882 30546 30894
rect 30494 30818 30546 30830
rect 37662 30882 37714 30894
rect 39902 30882 39954 30894
rect 43710 30882 43762 30894
rect 53118 30882 53170 30894
rect 39218 30830 39230 30882
rect 39282 30830 39294 30882
rect 42130 30830 42142 30882
rect 42194 30830 42206 30882
rect 46050 30830 46062 30882
rect 46114 30830 46126 30882
rect 49858 30830 49870 30882
rect 49922 30830 49934 30882
rect 51090 30830 51102 30882
rect 51154 30830 51166 30882
rect 37662 30818 37714 30830
rect 39902 30818 39954 30830
rect 43710 30818 43762 30830
rect 53118 30818 53170 30830
rect 56366 30882 56418 30894
rect 56366 30818 56418 30830
rect 56814 30882 56866 30894
rect 56814 30818 56866 30830
rect 57486 30882 57538 30894
rect 57486 30818 57538 30830
rect 26574 30770 26626 30782
rect 3602 30718 3614 30770
rect 3666 30718 3678 30770
rect 15698 30718 15710 30770
rect 15762 30718 15774 30770
rect 17490 30718 17502 30770
rect 17554 30767 17566 30770
rect 18162 30767 18174 30770
rect 17554 30721 18174 30767
rect 17554 30718 17566 30721
rect 18162 30718 18174 30721
rect 18226 30718 18238 30770
rect 26574 30706 26626 30718
rect 29822 30770 29874 30782
rect 29822 30706 29874 30718
rect 30718 30770 30770 30782
rect 32734 30770 32786 30782
rect 31042 30718 31054 30770
rect 31106 30718 31118 30770
rect 30718 30706 30770 30718
rect 32734 30706 32786 30718
rect 38894 30770 38946 30782
rect 48414 30770 48466 30782
rect 44034 30718 44046 30770
rect 44098 30767 44110 30770
rect 44370 30767 44382 30770
rect 44098 30721 44382 30767
rect 44098 30718 44110 30721
rect 44370 30718 44382 30721
rect 44434 30718 44446 30770
rect 46386 30718 46398 30770
rect 46450 30718 46462 30770
rect 38894 30706 38946 30718
rect 48414 30706 48466 30718
rect 57710 30770 57762 30782
rect 57710 30706 57762 30718
rect 58046 30770 58098 30782
rect 58046 30706 58098 30718
rect 1344 30602 59024 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 59024 30602
rect 1344 30516 59024 30550
rect 6862 30434 6914 30446
rect 6862 30370 6914 30382
rect 16830 30434 16882 30446
rect 16830 30370 16882 30382
rect 19630 30434 19682 30446
rect 19630 30370 19682 30382
rect 35534 30434 35586 30446
rect 35534 30370 35586 30382
rect 37886 30434 37938 30446
rect 42018 30382 42030 30434
rect 42082 30431 42094 30434
rect 43586 30431 43598 30434
rect 42082 30385 43598 30431
rect 42082 30382 42094 30385
rect 43586 30382 43598 30385
rect 43650 30382 43662 30434
rect 37886 30370 37938 30382
rect 12574 30322 12626 30334
rect 16606 30322 16658 30334
rect 8418 30270 8430 30322
rect 8482 30270 8494 30322
rect 9762 30270 9774 30322
rect 9826 30270 9838 30322
rect 12002 30270 12014 30322
rect 12066 30270 12078 30322
rect 15250 30270 15262 30322
rect 15314 30270 15326 30322
rect 12574 30258 12626 30270
rect 16606 30258 16658 30270
rect 26014 30322 26066 30334
rect 31726 30322 31778 30334
rect 28354 30270 28366 30322
rect 28418 30270 28430 30322
rect 26014 30258 26066 30270
rect 31726 30258 31778 30270
rect 44046 30322 44098 30334
rect 44046 30258 44098 30270
rect 47406 30322 47458 30334
rect 56590 30322 56642 30334
rect 48402 30270 48414 30322
rect 48466 30270 48478 30322
rect 49858 30270 49870 30322
rect 49922 30270 49934 30322
rect 57362 30270 57374 30322
rect 57426 30270 57438 30322
rect 47406 30258 47458 30270
rect 56590 30258 56642 30270
rect 4622 30210 4674 30222
rect 3042 30158 3054 30210
rect 3106 30158 3118 30210
rect 3266 30158 3278 30210
rect 3330 30158 3342 30210
rect 7198 30210 7250 30222
rect 9550 30210 9602 30222
rect 4622 30146 4674 30158
rect 4958 30154 5010 30166
rect 7970 30158 7982 30210
rect 8034 30158 8046 30210
rect 7198 30146 7250 30158
rect 9550 30146 9602 30158
rect 11006 30210 11058 30222
rect 11006 30146 11058 30158
rect 11118 30210 11170 30222
rect 11118 30146 11170 30158
rect 11902 30210 11954 30222
rect 11902 30146 11954 30158
rect 13694 30210 13746 30222
rect 16382 30210 16434 30222
rect 14354 30158 14366 30210
rect 14418 30158 14430 30210
rect 13694 30146 13746 30158
rect 16382 30146 16434 30158
rect 17278 30210 17330 30222
rect 17278 30146 17330 30158
rect 18174 30210 18226 30222
rect 19182 30210 19234 30222
rect 25230 30210 25282 30222
rect 25902 30210 25954 30222
rect 18386 30158 18398 30210
rect 18450 30158 18462 30210
rect 19394 30158 19406 30210
rect 19458 30158 19470 30210
rect 19730 30158 19742 30210
rect 19794 30158 19806 30210
rect 22642 30158 22654 30210
rect 22706 30158 22718 30210
rect 22978 30158 22990 30210
rect 23042 30158 23054 30210
rect 25330 30158 25342 30210
rect 25394 30158 25406 30210
rect 18174 30146 18226 30158
rect 19182 30146 19234 30158
rect 25230 30146 25282 30158
rect 25902 30146 25954 30158
rect 26798 30210 26850 30222
rect 36094 30210 36146 30222
rect 27794 30158 27806 30210
rect 27858 30158 27870 30210
rect 30370 30158 30382 30210
rect 30434 30158 30446 30210
rect 32386 30158 32398 30210
rect 32450 30158 32462 30210
rect 33282 30158 33294 30210
rect 33346 30158 33358 30210
rect 33618 30158 33630 30210
rect 33682 30158 33694 30210
rect 34066 30158 34078 30210
rect 34130 30158 34142 30210
rect 35858 30158 35870 30210
rect 35922 30158 35934 30210
rect 26798 30146 26850 30158
rect 36094 30146 36146 30158
rect 36206 30210 36258 30222
rect 36206 30146 36258 30158
rect 36766 30210 36818 30222
rect 42254 30210 42306 30222
rect 39442 30158 39454 30210
rect 39506 30158 39518 30210
rect 36766 30146 36818 30158
rect 42254 30146 42306 30158
rect 46398 30210 46450 30222
rect 46398 30146 46450 30158
rect 46846 30210 46898 30222
rect 52670 30210 52722 30222
rect 50082 30158 50094 30210
rect 50146 30158 50158 30210
rect 46846 30146 46898 30158
rect 52670 30146 52722 30158
rect 53678 30210 53730 30222
rect 53678 30146 53730 30158
rect 54126 30210 54178 30222
rect 54126 30146 54178 30158
rect 55470 30210 55522 30222
rect 55470 30146 55522 30158
rect 55694 30210 55746 30222
rect 57250 30158 57262 30210
rect 57314 30158 57326 30210
rect 55694 30146 55746 30158
rect 2370 30046 2382 30098
rect 2434 30046 2446 30098
rect 4958 30090 5010 30102
rect 9214 30098 9266 30110
rect 17726 30098 17778 30110
rect 25118 30098 25170 30110
rect 6290 30046 6302 30098
rect 6354 30046 6366 30098
rect 6514 30046 6526 30098
rect 6578 30046 6590 30098
rect 11666 30046 11678 30098
rect 11730 30046 11742 30098
rect 14130 30046 14142 30098
rect 14194 30046 14206 30098
rect 24210 30046 24222 30098
rect 24274 30046 24286 30098
rect 9214 30034 9266 30046
rect 17726 30034 17778 30046
rect 25118 30034 25170 30046
rect 25678 30098 25730 30110
rect 37550 30098 37602 30110
rect 43486 30098 43538 30110
rect 27570 30046 27582 30098
rect 27634 30046 27646 30098
rect 30706 30046 30718 30098
rect 30770 30046 30782 30098
rect 39218 30046 39230 30098
rect 39282 30046 39294 30098
rect 40562 30046 40574 30098
rect 40626 30046 40638 30098
rect 25678 30034 25730 30046
rect 37550 30034 37602 30046
rect 43486 30034 43538 30046
rect 48078 30098 48130 30110
rect 48078 30034 48130 30046
rect 49198 30098 49250 30110
rect 49198 30034 49250 30046
rect 50766 30098 50818 30110
rect 50766 30034 50818 30046
rect 53454 30098 53506 30110
rect 53454 30034 53506 30046
rect 58158 30098 58210 30110
rect 58158 30034 58210 30046
rect 1822 29986 1874 29998
rect 1822 29922 1874 29934
rect 4846 29986 4898 29998
rect 4846 29922 4898 29934
rect 10446 29986 10498 29998
rect 10446 29922 10498 29934
rect 11454 29986 11506 29998
rect 11454 29922 11506 29934
rect 12910 29986 12962 29998
rect 12910 29922 12962 29934
rect 17950 29986 18002 29998
rect 17950 29922 18002 29934
rect 18062 29986 18114 29998
rect 18062 29922 18114 29934
rect 19966 29986 20018 29998
rect 19966 29922 20018 29934
rect 20414 29986 20466 29998
rect 20414 29922 20466 29934
rect 20862 29986 20914 29998
rect 20862 29922 20914 29934
rect 21534 29986 21586 29998
rect 21534 29922 21586 29934
rect 22094 29986 22146 29998
rect 22094 29922 22146 29934
rect 29598 29986 29650 29998
rect 29598 29922 29650 29934
rect 35982 29986 36034 29998
rect 35982 29922 36034 29934
rect 37774 29986 37826 29998
rect 41246 29986 41298 29998
rect 40450 29934 40462 29986
rect 40514 29934 40526 29986
rect 37774 29922 37826 29934
rect 41246 29922 41298 29934
rect 41694 29986 41746 29998
rect 41694 29922 41746 29934
rect 42590 29986 42642 29998
rect 42590 29922 42642 29934
rect 43038 29986 43090 29998
rect 43038 29922 43090 29934
rect 46062 29986 46114 29998
rect 46062 29922 46114 29934
rect 47294 29986 47346 29998
rect 47294 29922 47346 29934
rect 47518 29986 47570 29998
rect 47518 29922 47570 29934
rect 48302 29986 48354 29998
rect 48302 29922 48354 29934
rect 51214 29986 51266 29998
rect 51214 29922 51266 29934
rect 53790 29986 53842 29998
rect 53790 29922 53842 29934
rect 54910 29986 54962 29998
rect 56018 29934 56030 29986
rect 56082 29934 56094 29986
rect 54910 29922 54962 29934
rect 1344 29818 59024 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 59024 29818
rect 1344 29732 59024 29766
rect 3502 29650 3554 29662
rect 3502 29586 3554 29598
rect 4286 29650 4338 29662
rect 4286 29586 4338 29598
rect 6078 29650 6130 29662
rect 6078 29586 6130 29598
rect 9886 29650 9938 29662
rect 12126 29650 12178 29662
rect 11330 29598 11342 29650
rect 11394 29598 11406 29650
rect 9886 29586 9938 29598
rect 12126 29586 12178 29598
rect 12686 29650 12738 29662
rect 12686 29586 12738 29598
rect 14590 29650 14642 29662
rect 14590 29586 14642 29598
rect 15262 29650 15314 29662
rect 15262 29586 15314 29598
rect 19518 29650 19570 29662
rect 19518 29586 19570 29598
rect 22430 29650 22482 29662
rect 22430 29586 22482 29598
rect 25678 29650 25730 29662
rect 25678 29586 25730 29598
rect 25790 29650 25842 29662
rect 25790 29586 25842 29598
rect 25902 29650 25954 29662
rect 32734 29650 32786 29662
rect 32050 29598 32062 29650
rect 32114 29598 32126 29650
rect 25902 29586 25954 29598
rect 32734 29586 32786 29598
rect 33854 29650 33906 29662
rect 33854 29586 33906 29598
rect 34974 29650 35026 29662
rect 34974 29586 35026 29598
rect 35870 29650 35922 29662
rect 35870 29586 35922 29598
rect 36430 29650 36482 29662
rect 36430 29586 36482 29598
rect 38894 29650 38946 29662
rect 38894 29586 38946 29598
rect 45166 29650 45218 29662
rect 45166 29586 45218 29598
rect 46286 29650 46338 29662
rect 46286 29586 46338 29598
rect 46398 29650 46450 29662
rect 46398 29586 46450 29598
rect 46958 29650 47010 29662
rect 46958 29586 47010 29598
rect 47742 29650 47794 29662
rect 47742 29586 47794 29598
rect 57822 29650 57874 29662
rect 57822 29586 57874 29598
rect 10782 29538 10834 29550
rect 2706 29486 2718 29538
rect 2770 29486 2782 29538
rect 5282 29486 5294 29538
rect 5346 29486 5358 29538
rect 8866 29486 8878 29538
rect 8930 29486 8942 29538
rect 10782 29474 10834 29486
rect 11678 29538 11730 29550
rect 11678 29474 11730 29486
rect 13246 29538 13298 29550
rect 17950 29538 18002 29550
rect 14018 29486 14030 29538
rect 14082 29486 14094 29538
rect 13246 29474 13298 29486
rect 17950 29474 18002 29486
rect 18174 29538 18226 29550
rect 18174 29474 18226 29486
rect 19294 29538 19346 29550
rect 27134 29538 27186 29550
rect 20402 29486 20414 29538
rect 20466 29486 20478 29538
rect 24546 29486 24558 29538
rect 24610 29486 24622 29538
rect 19294 29474 19346 29486
rect 27134 29474 27186 29486
rect 27246 29538 27298 29550
rect 33630 29538 33682 29550
rect 29138 29486 29150 29538
rect 29202 29486 29214 29538
rect 30370 29486 30382 29538
rect 30434 29486 30446 29538
rect 32498 29486 32510 29538
rect 32562 29486 32574 29538
rect 27246 29474 27298 29486
rect 33630 29474 33682 29486
rect 44382 29538 44434 29550
rect 44382 29474 44434 29486
rect 53006 29538 53058 29550
rect 53006 29474 53058 29486
rect 57486 29538 57538 29550
rect 57486 29474 57538 29486
rect 4622 29426 4674 29438
rect 9774 29426 9826 29438
rect 5394 29374 5406 29426
rect 5458 29374 5470 29426
rect 6738 29374 6750 29426
rect 6802 29374 6814 29426
rect 7858 29374 7870 29426
rect 7922 29374 7934 29426
rect 4622 29362 4674 29374
rect 9774 29362 9826 29374
rect 11342 29426 11394 29438
rect 11342 29362 11394 29374
rect 13806 29426 13858 29438
rect 15150 29426 15202 29438
rect 14354 29374 14366 29426
rect 14418 29374 14430 29426
rect 13806 29362 13858 29374
rect 15150 29362 15202 29374
rect 16158 29426 16210 29438
rect 26910 29426 26962 29438
rect 31950 29426 32002 29438
rect 34750 29426 34802 29438
rect 20290 29374 20302 29426
rect 20354 29374 20366 29426
rect 21298 29374 21310 29426
rect 21362 29374 21374 29426
rect 23426 29374 23438 29426
rect 23490 29374 23502 29426
rect 26114 29374 26126 29426
rect 26178 29374 26190 29426
rect 26450 29374 26462 29426
rect 26514 29374 26526 29426
rect 28130 29374 28142 29426
rect 28194 29374 28206 29426
rect 28466 29374 28478 29426
rect 28530 29374 28542 29426
rect 30818 29374 30830 29426
rect 30882 29374 30894 29426
rect 31154 29374 31166 29426
rect 31218 29374 31230 29426
rect 34514 29374 34526 29426
rect 34578 29374 34590 29426
rect 16158 29362 16210 29374
rect 26910 29362 26962 29374
rect 31950 29362 32002 29374
rect 34750 29362 34802 29374
rect 35086 29426 35138 29438
rect 35086 29362 35138 29374
rect 35758 29426 35810 29438
rect 35758 29362 35810 29374
rect 36094 29426 36146 29438
rect 39790 29426 39842 29438
rect 37762 29374 37774 29426
rect 37826 29374 37838 29426
rect 36094 29362 36146 29374
rect 39790 29362 39842 29374
rect 40014 29426 40066 29438
rect 40014 29362 40066 29374
rect 40238 29426 40290 29438
rect 40238 29362 40290 29374
rect 40462 29426 40514 29438
rect 40462 29362 40514 29374
rect 40686 29426 40738 29438
rect 40686 29362 40738 29374
rect 41694 29426 41746 29438
rect 52110 29426 52162 29438
rect 57710 29426 57762 29438
rect 41906 29374 41918 29426
rect 41970 29374 41982 29426
rect 43474 29374 43486 29426
rect 43538 29374 43550 29426
rect 52434 29374 52446 29426
rect 52498 29374 52510 29426
rect 53890 29374 53902 29426
rect 53954 29374 53966 29426
rect 41694 29362 41746 29374
rect 52110 29362 52162 29374
rect 57710 29362 57762 29374
rect 58046 29426 58098 29438
rect 58046 29362 58098 29374
rect 11006 29314 11058 29326
rect 2706 29262 2718 29314
rect 2770 29262 2782 29314
rect 8306 29262 8318 29314
rect 8370 29262 8382 29314
rect 11006 29250 11058 29262
rect 16494 29314 16546 29326
rect 16494 29250 16546 29262
rect 16942 29314 16994 29326
rect 16942 29250 16994 29262
rect 18846 29314 18898 29326
rect 21086 29314 21138 29326
rect 29822 29314 29874 29326
rect 19618 29262 19630 29314
rect 19682 29262 19694 29314
rect 20514 29262 20526 29314
rect 20578 29262 20590 29314
rect 23538 29262 23550 29314
rect 23602 29262 23614 29314
rect 28578 29262 28590 29314
rect 28642 29262 28654 29314
rect 18846 29250 18898 29262
rect 21086 29250 21138 29262
rect 29822 29250 29874 29262
rect 34862 29314 34914 29326
rect 42590 29314 42642 29326
rect 37538 29262 37550 29314
rect 37602 29262 37614 29314
rect 40562 29262 40574 29314
rect 40626 29262 40638 29314
rect 34862 29250 34914 29262
rect 42590 29250 42642 29262
rect 44046 29314 44098 29326
rect 44046 29250 44098 29262
rect 45726 29314 45778 29326
rect 45726 29250 45778 29262
rect 46174 29314 46226 29326
rect 54574 29314 54626 29326
rect 54114 29262 54126 29314
rect 54178 29262 54190 29314
rect 46174 29250 46226 29262
rect 54574 29250 54626 29262
rect 55134 29314 55186 29326
rect 55134 29250 55186 29262
rect 55358 29314 55410 29326
rect 55358 29250 55410 29262
rect 56142 29314 56194 29326
rect 56142 29250 56194 29262
rect 56702 29314 56754 29326
rect 56702 29250 56754 29262
rect 9886 29202 9938 29214
rect 9886 29138 9938 29150
rect 11230 29202 11282 29214
rect 15262 29202 15314 29214
rect 14354 29150 14366 29202
rect 14418 29150 14430 29202
rect 11230 29138 11282 29150
rect 15262 29138 15314 29150
rect 18286 29202 18338 29214
rect 18286 29138 18338 29150
rect 33966 29202 34018 29214
rect 43150 29202 43202 29214
rect 38322 29150 38334 29202
rect 38386 29150 38398 29202
rect 33966 29138 34018 29150
rect 43150 29138 43202 29150
rect 43486 29202 43538 29214
rect 43486 29138 43538 29150
rect 55694 29202 55746 29214
rect 55694 29138 55746 29150
rect 1344 29034 59024 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 59024 29034
rect 1344 28948 59024 28982
rect 3950 28866 4002 28878
rect 3950 28802 4002 28814
rect 10334 28866 10386 28878
rect 10334 28802 10386 28814
rect 18846 28866 18898 28878
rect 18846 28802 18898 28814
rect 28030 28866 28082 28878
rect 28030 28802 28082 28814
rect 34750 28866 34802 28878
rect 40014 28866 40066 28878
rect 36418 28814 36430 28866
rect 36482 28863 36494 28866
rect 36642 28863 36654 28866
rect 36482 28817 36654 28863
rect 36482 28814 36494 28817
rect 36642 28814 36654 28817
rect 36706 28814 36718 28866
rect 34750 28802 34802 28814
rect 40014 28802 40066 28814
rect 48078 28866 48130 28878
rect 48078 28802 48130 28814
rect 52334 28866 52386 28878
rect 52658 28814 52670 28866
rect 52722 28814 52734 28866
rect 52334 28802 52386 28814
rect 2046 28754 2098 28766
rect 4510 28754 4562 28766
rect 3154 28702 3166 28754
rect 3218 28702 3230 28754
rect 2046 28690 2098 28702
rect 4510 28690 4562 28702
rect 5854 28754 5906 28766
rect 5854 28690 5906 28702
rect 6414 28754 6466 28766
rect 6414 28690 6466 28702
rect 10894 28754 10946 28766
rect 10894 28690 10946 28702
rect 11790 28754 11842 28766
rect 11790 28690 11842 28702
rect 13694 28754 13746 28766
rect 13694 28690 13746 28702
rect 14926 28754 14978 28766
rect 25230 28754 25282 28766
rect 16930 28702 16942 28754
rect 16994 28702 17006 28754
rect 23538 28702 23550 28754
rect 23602 28702 23614 28754
rect 24546 28702 24558 28754
rect 24610 28702 24622 28754
rect 14926 28690 14978 28702
rect 25230 28690 25282 28702
rect 25790 28754 25842 28766
rect 25790 28690 25842 28702
rect 35870 28754 35922 28766
rect 35870 28690 35922 28702
rect 36654 28754 36706 28766
rect 36654 28690 36706 28702
rect 37438 28754 37490 28766
rect 37438 28690 37490 28702
rect 37886 28754 37938 28766
rect 37886 28690 37938 28702
rect 38334 28754 38386 28766
rect 38334 28690 38386 28702
rect 38782 28754 38834 28766
rect 38782 28690 38834 28702
rect 40350 28754 40402 28766
rect 40350 28690 40402 28702
rect 40798 28754 40850 28766
rect 40798 28690 40850 28702
rect 43934 28754 43986 28766
rect 43934 28690 43986 28702
rect 45390 28754 45442 28766
rect 45390 28690 45442 28702
rect 45838 28754 45890 28766
rect 45838 28690 45890 28702
rect 46286 28754 46338 28766
rect 46286 28690 46338 28702
rect 47070 28754 47122 28766
rect 47070 28690 47122 28702
rect 49310 28754 49362 28766
rect 49310 28690 49362 28702
rect 54350 28754 54402 28766
rect 57822 28754 57874 28766
rect 55122 28702 55134 28754
rect 55186 28702 55198 28754
rect 54350 28690 54402 28702
rect 57822 28690 57874 28702
rect 4958 28642 5010 28654
rect 9102 28642 9154 28654
rect 3042 28590 3054 28642
rect 3106 28590 3118 28642
rect 8306 28590 8318 28642
rect 8370 28590 8382 28642
rect 4958 28578 5010 28590
rect 9102 28578 9154 28590
rect 9550 28642 9602 28654
rect 12686 28642 12738 28654
rect 10658 28590 10670 28642
rect 10722 28590 10734 28642
rect 9550 28578 9602 28590
rect 12686 28578 12738 28590
rect 12910 28642 12962 28654
rect 19070 28642 19122 28654
rect 14130 28590 14142 28642
rect 14194 28590 14206 28642
rect 15362 28590 15374 28642
rect 15426 28590 15438 28642
rect 17154 28590 17166 28642
rect 17218 28590 17230 28642
rect 17490 28590 17502 28642
rect 17554 28590 17566 28642
rect 12910 28578 12962 28590
rect 19070 28578 19122 28590
rect 19294 28642 19346 28654
rect 19294 28578 19346 28590
rect 20526 28642 20578 28654
rect 20526 28578 20578 28590
rect 20974 28642 21026 28654
rect 26238 28642 26290 28654
rect 21970 28590 21982 28642
rect 22034 28590 22046 28642
rect 23650 28590 23662 28642
rect 23714 28590 23726 28642
rect 20974 28578 21026 28590
rect 26238 28578 26290 28590
rect 27694 28642 27746 28654
rect 27694 28578 27746 28590
rect 27806 28642 27858 28654
rect 35086 28642 35138 28654
rect 30146 28590 30158 28642
rect 30210 28590 30222 28642
rect 31378 28590 31390 28642
rect 31442 28590 31454 28642
rect 31602 28590 31614 28642
rect 31666 28590 31678 28642
rect 32274 28590 32286 28642
rect 32338 28590 32350 28642
rect 27806 28578 27858 28590
rect 35086 28578 35138 28590
rect 35982 28642 36034 28654
rect 35982 28578 36034 28590
rect 42926 28642 42978 28654
rect 42926 28578 42978 28590
rect 43486 28642 43538 28654
rect 49870 28642 49922 28654
rect 47170 28590 47182 28642
rect 47234 28590 47246 28642
rect 48290 28590 48302 28642
rect 48354 28590 48366 28642
rect 43486 28578 43538 28590
rect 49870 28578 49922 28590
rect 50094 28642 50146 28654
rect 52110 28642 52162 28654
rect 50418 28590 50430 28642
rect 50482 28590 50494 28642
rect 50094 28578 50146 28590
rect 52110 28578 52162 28590
rect 53342 28642 53394 28654
rect 57934 28642 57986 28654
rect 55010 28590 55022 28642
rect 55074 28590 55086 28642
rect 56354 28590 56366 28642
rect 56418 28590 56430 28642
rect 58258 28590 58270 28642
rect 58322 28590 58334 28642
rect 53342 28578 53394 28590
rect 57934 28578 57986 28590
rect 9662 28530 9714 28542
rect 7074 28478 7086 28530
rect 7138 28478 7150 28530
rect 9662 28466 9714 28478
rect 12350 28530 12402 28542
rect 18622 28530 18674 28542
rect 27022 28530 27074 28542
rect 36094 28530 36146 28542
rect 14466 28478 14478 28530
rect 14530 28478 14542 28530
rect 14914 28478 14926 28530
rect 14978 28478 14990 28530
rect 22194 28478 22206 28530
rect 22258 28478 22270 28530
rect 28578 28478 28590 28530
rect 28642 28478 28654 28530
rect 29922 28478 29934 28530
rect 29986 28478 29998 28530
rect 30930 28478 30942 28530
rect 30994 28478 31006 28530
rect 32834 28478 32846 28530
rect 32898 28478 32910 28530
rect 34178 28478 34190 28530
rect 34242 28478 34254 28530
rect 34514 28478 34526 28530
rect 34578 28478 34590 28530
rect 12350 28466 12402 28478
rect 18622 28466 18674 28478
rect 27022 28466 27074 28478
rect 36094 28466 36146 28478
rect 39454 28530 39506 28542
rect 39454 28466 39506 28478
rect 39678 28530 39730 28542
rect 39678 28466 39730 28478
rect 41582 28530 41634 28542
rect 41582 28466 41634 28478
rect 41918 28530 41970 28542
rect 41918 28466 41970 28478
rect 43710 28530 43762 28542
rect 43710 28466 43762 28478
rect 44046 28530 44098 28542
rect 44046 28466 44098 28478
rect 57150 28530 57202 28542
rect 57150 28466 57202 28478
rect 57710 28530 57762 28542
rect 57710 28466 57762 28478
rect 9774 28418 9826 28430
rect 7970 28366 7982 28418
rect 8034 28366 8046 28418
rect 9774 28354 9826 28366
rect 10782 28418 10834 28430
rect 10782 28354 10834 28366
rect 11006 28418 11058 28430
rect 11006 28354 11058 28366
rect 12574 28418 12626 28430
rect 19742 28418 19794 28430
rect 33182 28418 33234 28430
rect 17826 28366 17838 28418
rect 17890 28366 17902 28418
rect 30146 28366 30158 28418
rect 30210 28366 30222 28418
rect 32498 28366 32510 28418
rect 32562 28366 32574 28418
rect 12574 28354 12626 28366
rect 19742 28354 19794 28366
rect 33182 28354 33234 28366
rect 39902 28418 39954 28430
rect 39902 28354 39954 28366
rect 41694 28418 41746 28430
rect 41694 28354 41746 28366
rect 42366 28418 42418 28430
rect 42366 28354 42418 28366
rect 44606 28418 44658 28430
rect 44606 28354 44658 28366
rect 48638 28418 48690 28430
rect 48638 28354 48690 28366
rect 1344 28250 59024 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 59024 28250
rect 1344 28164 59024 28198
rect 5294 28082 5346 28094
rect 5294 28018 5346 28030
rect 6078 28082 6130 28094
rect 6078 28018 6130 28030
rect 13246 28082 13298 28094
rect 13246 28018 13298 28030
rect 13806 28082 13858 28094
rect 13806 28018 13858 28030
rect 14254 28082 14306 28094
rect 16606 28082 16658 28094
rect 15698 28030 15710 28082
rect 15762 28030 15774 28082
rect 14254 28018 14306 28030
rect 16606 28018 16658 28030
rect 20862 28082 20914 28094
rect 20862 28018 20914 28030
rect 22318 28082 22370 28094
rect 22318 28018 22370 28030
rect 23214 28082 23266 28094
rect 23214 28018 23266 28030
rect 23662 28082 23714 28094
rect 23662 28018 23714 28030
rect 24110 28082 24162 28094
rect 24110 28018 24162 28030
rect 25006 28082 25058 28094
rect 25006 28018 25058 28030
rect 29374 28082 29426 28094
rect 29374 28018 29426 28030
rect 32734 28082 32786 28094
rect 32734 28018 32786 28030
rect 34190 28082 34242 28094
rect 34190 28018 34242 28030
rect 38110 28082 38162 28094
rect 38110 28018 38162 28030
rect 41918 28082 41970 28094
rect 41918 28018 41970 28030
rect 18510 27970 18562 27982
rect 4162 27918 4174 27970
rect 4226 27918 4238 27970
rect 8978 27918 8990 27970
rect 9042 27918 9054 27970
rect 14690 27918 14702 27970
rect 14754 27918 14766 27970
rect 18510 27906 18562 27918
rect 25902 27970 25954 27982
rect 33630 27970 33682 27982
rect 30258 27918 30270 27970
rect 30322 27918 30334 27970
rect 31826 27918 31838 27970
rect 31890 27918 31902 27970
rect 25902 27906 25954 27918
rect 33630 27906 33682 27918
rect 36318 27970 36370 27982
rect 45614 27970 45666 27982
rect 48638 27970 48690 27982
rect 36978 27918 36990 27970
rect 37042 27918 37054 27970
rect 37650 27918 37662 27970
rect 37714 27918 37726 27970
rect 47394 27918 47406 27970
rect 47458 27918 47470 27970
rect 49858 27918 49870 27970
rect 49922 27918 49934 27970
rect 36318 27906 36370 27918
rect 45614 27906 45666 27918
rect 48638 27906 48690 27918
rect 9774 27858 9826 27870
rect 19854 27858 19906 27870
rect 22766 27858 22818 27870
rect 2482 27806 2494 27858
rect 2546 27806 2558 27858
rect 3042 27806 3054 27858
rect 3106 27806 3118 27858
rect 6962 27806 6974 27858
rect 7026 27806 7038 27858
rect 8418 27806 8430 27858
rect 8482 27806 8494 27858
rect 9986 27806 9998 27858
rect 10050 27806 10062 27858
rect 11890 27806 11902 27858
rect 11954 27806 11966 27858
rect 15138 27806 15150 27858
rect 15202 27806 15214 27858
rect 15586 27806 15598 27858
rect 15650 27806 15662 27858
rect 20290 27806 20302 27858
rect 20354 27806 20366 27858
rect 9774 27794 9826 27806
rect 19854 27794 19906 27806
rect 22766 27794 22818 27806
rect 24558 27858 24610 27870
rect 35422 27858 35474 27870
rect 27682 27806 27694 27858
rect 27746 27806 27758 27858
rect 28018 27806 28030 27858
rect 28082 27806 28094 27858
rect 29922 27806 29934 27858
rect 29986 27806 29998 27858
rect 32162 27806 32174 27858
rect 32226 27806 32238 27858
rect 35634 27806 35646 27858
rect 35698 27806 35710 27858
rect 37090 27806 37102 27858
rect 37154 27806 37166 27858
rect 39554 27806 39566 27858
rect 39618 27806 39630 27858
rect 43026 27806 43038 27858
rect 43090 27806 43102 27858
rect 44146 27806 44158 27858
rect 44210 27806 44222 27858
rect 45938 27806 45950 27858
rect 46002 27806 46014 27858
rect 46498 27806 46510 27858
rect 46562 27806 46574 27858
rect 51090 27806 51102 27858
rect 51154 27806 51166 27858
rect 52658 27806 52670 27858
rect 52722 27806 52734 27858
rect 24558 27794 24610 27806
rect 35422 27794 35474 27806
rect 1934 27746 1986 27758
rect 17054 27746 17106 27758
rect 8082 27694 8094 27746
rect 8146 27694 8158 27746
rect 1934 27682 1986 27694
rect 17054 27682 17106 27694
rect 18062 27746 18114 27758
rect 19966 27746 20018 27758
rect 26462 27746 26514 27758
rect 40014 27746 40066 27758
rect 18834 27694 18846 27746
rect 18898 27694 18910 27746
rect 21298 27694 21310 27746
rect 21362 27694 21374 27746
rect 26002 27694 26014 27746
rect 26066 27694 26078 27746
rect 28578 27694 28590 27746
rect 28642 27694 28654 27746
rect 39106 27694 39118 27746
rect 39170 27694 39182 27746
rect 18062 27682 18114 27694
rect 19966 27682 20018 27694
rect 26462 27682 26514 27694
rect 40014 27682 40066 27694
rect 40462 27746 40514 27758
rect 40462 27682 40514 27694
rect 41470 27746 41522 27758
rect 48190 27746 48242 27758
rect 51774 27746 51826 27758
rect 53342 27746 53394 27758
rect 43138 27694 43150 27746
rect 43202 27694 43214 27746
rect 44930 27694 44942 27746
rect 44994 27694 45006 27746
rect 49634 27694 49646 27746
rect 49698 27694 49710 27746
rect 52434 27694 52446 27746
rect 52498 27694 52510 27746
rect 41470 27682 41522 27694
rect 48190 27682 48242 27694
rect 51774 27682 51826 27694
rect 53342 27682 53394 27694
rect 25678 27634 25730 27646
rect 10098 27582 10110 27634
rect 10162 27582 10174 27634
rect 25678 27570 25730 27582
rect 33854 27634 33906 27646
rect 33854 27570 33906 27582
rect 45950 27634 46002 27646
rect 45950 27570 46002 27582
rect 1344 27466 59024 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 59024 27466
rect 1344 27380 59024 27414
rect 14590 27298 14642 27310
rect 45614 27298 45666 27310
rect 22978 27246 22990 27298
rect 23042 27246 23054 27298
rect 14590 27234 14642 27246
rect 45614 27234 45666 27246
rect 48414 27298 48466 27310
rect 48414 27234 48466 27246
rect 50654 27298 50706 27310
rect 50654 27234 50706 27246
rect 8430 27186 8482 27198
rect 10334 27186 10386 27198
rect 4162 27134 4174 27186
rect 4226 27134 4238 27186
rect 5730 27134 5742 27186
rect 5794 27134 5806 27186
rect 9426 27134 9438 27186
rect 9490 27134 9502 27186
rect 8430 27122 8482 27134
rect 10334 27122 10386 27134
rect 12126 27186 12178 27198
rect 12126 27122 12178 27134
rect 20862 27186 20914 27198
rect 27134 27186 27186 27198
rect 29486 27186 29538 27198
rect 23986 27134 23998 27186
rect 24050 27134 24062 27186
rect 26002 27134 26014 27186
rect 26066 27134 26078 27186
rect 28690 27134 28702 27186
rect 28754 27134 28766 27186
rect 20862 27122 20914 27134
rect 27134 27122 27186 27134
rect 29486 27122 29538 27134
rect 29934 27186 29986 27198
rect 41358 27186 41410 27198
rect 38882 27134 38894 27186
rect 38946 27134 38958 27186
rect 29934 27122 29986 27134
rect 41358 27122 41410 27134
rect 41806 27186 41858 27198
rect 41806 27122 41858 27134
rect 42702 27186 42754 27198
rect 42702 27122 42754 27134
rect 43598 27186 43650 27198
rect 43598 27122 43650 27134
rect 46174 27186 46226 27198
rect 46174 27122 46226 27134
rect 48974 27186 49026 27198
rect 48974 27122 49026 27134
rect 49534 27186 49586 27198
rect 50430 27186 50482 27198
rect 49746 27134 49758 27186
rect 49810 27134 49822 27186
rect 49534 27122 49586 27134
rect 50430 27122 50482 27134
rect 50878 27186 50930 27198
rect 51202 27134 51214 27186
rect 51266 27134 51278 27186
rect 57362 27134 57374 27186
rect 57426 27134 57438 27186
rect 50878 27122 50930 27134
rect 11230 27074 11282 27086
rect 3042 27022 3054 27074
rect 3106 27022 3118 27074
rect 3378 27022 3390 27074
rect 3442 27022 3454 27074
rect 6738 27022 6750 27074
rect 6802 27022 6814 27074
rect 7298 27022 7310 27074
rect 7362 27022 7374 27074
rect 11230 27010 11282 27022
rect 11454 27074 11506 27086
rect 11454 27010 11506 27022
rect 12014 27074 12066 27086
rect 15374 27074 15426 27086
rect 13906 27022 13918 27074
rect 13970 27022 13982 27074
rect 12014 27010 12066 27022
rect 15374 27010 15426 27022
rect 17950 27074 18002 27086
rect 27022 27074 27074 27086
rect 36206 27074 36258 27086
rect 18498 27022 18510 27074
rect 18562 27022 18574 27074
rect 22194 27022 22206 27074
rect 22258 27022 22270 27074
rect 24210 27022 24222 27074
rect 24274 27022 24286 27074
rect 25778 27022 25790 27074
rect 25842 27022 25854 27074
rect 28130 27022 28142 27074
rect 28194 27022 28206 27074
rect 30930 27022 30942 27074
rect 30994 27022 31006 27074
rect 32498 27022 32510 27074
rect 32562 27022 32574 27074
rect 34178 27022 34190 27074
rect 34242 27022 34254 27074
rect 34738 27022 34750 27074
rect 34802 27022 34814 27074
rect 17950 27010 18002 27022
rect 27022 27010 27074 27022
rect 36206 27010 36258 27022
rect 36318 27074 36370 27086
rect 36318 27010 36370 27022
rect 36542 27074 36594 27086
rect 36542 27010 36594 27022
rect 37774 27074 37826 27086
rect 40574 27074 40626 27086
rect 39218 27022 39230 27074
rect 39282 27022 39294 27074
rect 37774 27010 37826 27022
rect 40574 27010 40626 27022
rect 40910 27074 40962 27086
rect 40910 27010 40962 27022
rect 45838 27074 45890 27086
rect 45838 27010 45890 27022
rect 46062 27074 46114 27086
rect 46062 27010 46114 27022
rect 47518 27074 47570 27086
rect 47518 27010 47570 27022
rect 47742 27074 47794 27086
rect 47742 27010 47794 27022
rect 51102 27074 51154 27086
rect 51102 27010 51154 27022
rect 52782 27074 52834 27086
rect 52782 27010 52834 27022
rect 53678 27074 53730 27086
rect 58034 27022 58046 27074
rect 58098 27022 58110 27074
rect 53678 27010 53730 27022
rect 4958 26962 5010 26974
rect 4958 26898 5010 26910
rect 10894 26962 10946 26974
rect 10894 26898 10946 26910
rect 12462 26962 12514 26974
rect 12462 26898 12514 26910
rect 15822 26962 15874 26974
rect 18958 26962 19010 26974
rect 24894 26962 24946 26974
rect 16370 26910 16382 26962
rect 16434 26910 16446 26962
rect 21858 26910 21870 26962
rect 21922 26910 21934 26962
rect 15822 26898 15874 26910
rect 18958 26898 19010 26910
rect 24894 26898 24946 26910
rect 26462 26962 26514 26974
rect 26462 26898 26514 26910
rect 27246 26962 27298 26974
rect 36654 26962 36706 26974
rect 42254 26962 42306 26974
rect 28242 26910 28254 26962
rect 28306 26910 28318 26962
rect 31266 26910 31278 26962
rect 31330 26910 31342 26962
rect 32386 26910 32398 26962
rect 32450 26910 32462 26962
rect 39442 26910 39454 26962
rect 39506 26910 39518 26962
rect 27246 26898 27298 26910
rect 36654 26898 36706 26910
rect 42254 26898 42306 26910
rect 43150 26962 43202 26974
rect 43150 26898 43202 26910
rect 44046 26962 44098 26974
rect 44046 26898 44098 26910
rect 47182 26962 47234 26974
rect 47182 26898 47234 26910
rect 48302 26962 48354 26974
rect 48302 26898 48354 26910
rect 51326 26962 51378 26974
rect 51326 26898 51378 26910
rect 51998 26962 52050 26974
rect 51998 26898 52050 26910
rect 53454 26962 53506 26974
rect 53454 26898 53506 26910
rect 54014 26962 54066 26974
rect 54014 26898 54066 26910
rect 57150 26962 57202 26974
rect 57150 26898 57202 26910
rect 1934 26850 1986 26862
rect 1934 26786 1986 26798
rect 7982 26850 8034 26862
rect 7982 26786 8034 26798
rect 8990 26850 9042 26862
rect 8990 26786 9042 26798
rect 11006 26850 11058 26862
rect 11006 26786 11058 26798
rect 12238 26850 12290 26862
rect 27470 26850 27522 26862
rect 36430 26850 36482 26862
rect 19842 26798 19854 26850
rect 19906 26798 19918 26850
rect 32498 26798 32510 26850
rect 32562 26798 32574 26850
rect 12238 26786 12290 26798
rect 27470 26786 27522 26798
rect 36430 26786 36482 26798
rect 40798 26850 40850 26862
rect 40798 26786 40850 26798
rect 44494 26850 44546 26862
rect 44494 26786 44546 26798
rect 46286 26850 46338 26862
rect 46286 26786 46338 26798
rect 48414 26850 48466 26862
rect 48414 26786 48466 26798
rect 49758 26850 49810 26862
rect 49758 26786 49810 26798
rect 53678 26850 53730 26862
rect 53678 26786 53730 26798
rect 1344 26682 59024 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 59024 26682
rect 1344 26596 59024 26630
rect 1934 26514 1986 26526
rect 1934 26450 1986 26462
rect 2942 26514 2994 26526
rect 2942 26450 2994 26462
rect 3726 26514 3778 26526
rect 3726 26450 3778 26462
rect 10334 26514 10386 26526
rect 10334 26450 10386 26462
rect 20862 26514 20914 26526
rect 20862 26450 20914 26462
rect 23886 26514 23938 26526
rect 23886 26450 23938 26462
rect 24558 26514 24610 26526
rect 28590 26514 28642 26526
rect 26226 26462 26238 26514
rect 26290 26462 26302 26514
rect 24558 26450 24610 26462
rect 28590 26450 28642 26462
rect 30830 26514 30882 26526
rect 30830 26450 30882 26462
rect 32174 26514 32226 26526
rect 32174 26450 32226 26462
rect 32958 26514 33010 26526
rect 32958 26450 33010 26462
rect 35198 26514 35250 26526
rect 35198 26450 35250 26462
rect 35310 26514 35362 26526
rect 35310 26450 35362 26462
rect 37326 26514 37378 26526
rect 37326 26450 37378 26462
rect 37774 26514 37826 26526
rect 37774 26450 37826 26462
rect 38110 26514 38162 26526
rect 38110 26450 38162 26462
rect 38558 26514 38610 26526
rect 38558 26450 38610 26462
rect 40462 26514 40514 26526
rect 40462 26450 40514 26462
rect 41806 26514 41858 26526
rect 41806 26450 41858 26462
rect 43710 26514 43762 26526
rect 43710 26450 43762 26462
rect 45390 26514 45442 26526
rect 45390 26450 45442 26462
rect 46958 26514 47010 26526
rect 46958 26450 47010 26462
rect 47406 26514 47458 26526
rect 47406 26450 47458 26462
rect 50430 26514 50482 26526
rect 50430 26450 50482 26462
rect 52110 26514 52162 26526
rect 52110 26450 52162 26462
rect 54462 26514 54514 26526
rect 54462 26450 54514 26462
rect 56478 26514 56530 26526
rect 56478 26450 56530 26462
rect 56590 26514 56642 26526
rect 56590 26450 56642 26462
rect 11678 26402 11730 26414
rect 4834 26350 4846 26402
rect 4898 26350 4910 26402
rect 11678 26338 11730 26350
rect 14030 26402 14082 26414
rect 23662 26402 23714 26414
rect 21746 26350 21758 26402
rect 21810 26350 21822 26402
rect 22754 26350 22766 26402
rect 22818 26350 22830 26402
rect 14030 26338 14082 26350
rect 23662 26338 23714 26350
rect 24894 26402 24946 26414
rect 24894 26338 24946 26350
rect 25678 26402 25730 26414
rect 25678 26338 25730 26350
rect 29486 26402 29538 26414
rect 29486 26338 29538 26350
rect 30046 26402 30098 26414
rect 30046 26338 30098 26350
rect 33966 26402 34018 26414
rect 33966 26338 34018 26350
rect 34974 26402 35026 26414
rect 43598 26402 43650 26414
rect 39218 26350 39230 26402
rect 39282 26350 39294 26402
rect 34974 26338 35026 26350
rect 43598 26338 43650 26350
rect 46062 26402 46114 26414
rect 46062 26338 46114 26350
rect 54574 26402 54626 26414
rect 54574 26338 54626 26350
rect 56254 26402 56306 26414
rect 56254 26338 56306 26350
rect 2382 26290 2434 26302
rect 2382 26226 2434 26238
rect 4174 26290 4226 26302
rect 10670 26290 10722 26302
rect 11230 26290 11282 26302
rect 5394 26238 5406 26290
rect 5458 26238 5470 26290
rect 5954 26238 5966 26290
rect 6018 26238 6030 26290
rect 8642 26238 8654 26290
rect 8706 26238 8718 26290
rect 10994 26238 11006 26290
rect 11058 26238 11070 26290
rect 4174 26226 4226 26238
rect 10670 26226 10722 26238
rect 11230 26226 11282 26238
rect 12574 26290 12626 26302
rect 12574 26226 12626 26238
rect 14142 26290 14194 26302
rect 23550 26290 23602 26302
rect 27134 26290 27186 26302
rect 15362 26238 15374 26290
rect 15426 26238 15438 26290
rect 18722 26238 18734 26290
rect 18786 26238 18798 26290
rect 21970 26238 21982 26290
rect 22034 26238 22046 26290
rect 26898 26238 26910 26290
rect 26962 26238 26974 26290
rect 14142 26226 14194 26238
rect 23550 26226 23602 26238
rect 27134 26226 27186 26238
rect 27358 26290 27410 26302
rect 28254 26290 28306 26302
rect 27570 26238 27582 26290
rect 27634 26238 27646 26290
rect 27358 26226 27410 26238
rect 28254 26226 28306 26238
rect 28366 26290 28418 26302
rect 28366 26226 28418 26238
rect 28702 26290 28754 26302
rect 33742 26290 33794 26302
rect 29698 26238 29710 26290
rect 29762 26238 29774 26290
rect 28702 26226 28754 26238
rect 33742 26226 33794 26238
rect 33854 26290 33906 26302
rect 33854 26226 33906 26238
rect 34078 26290 34130 26302
rect 34078 26226 34130 26238
rect 34190 26290 34242 26302
rect 34190 26226 34242 26238
rect 35422 26290 35474 26302
rect 41694 26290 41746 26302
rect 39554 26238 39566 26290
rect 39618 26238 39630 26290
rect 40114 26238 40126 26290
rect 40178 26238 40190 26290
rect 35422 26226 35474 26238
rect 41694 26226 41746 26238
rect 41918 26290 41970 26302
rect 41918 26226 41970 26238
rect 43150 26290 43202 26302
rect 43150 26226 43202 26238
rect 43822 26290 43874 26302
rect 43822 26226 43874 26238
rect 45614 26290 45666 26302
rect 45614 26226 45666 26238
rect 48302 26290 48354 26302
rect 56702 26290 56754 26302
rect 52882 26238 52894 26290
rect 52946 26238 52958 26290
rect 48302 26226 48354 26238
rect 56702 26226 56754 26238
rect 57598 26290 57650 26302
rect 57922 26238 57934 26290
rect 57986 26238 57998 26290
rect 57598 26226 57650 26238
rect 3278 26178 3330 26190
rect 9774 26178 9826 26190
rect 7522 26126 7534 26178
rect 7586 26126 7598 26178
rect 8530 26126 8542 26178
rect 8594 26126 8606 26178
rect 3278 26114 3330 26126
rect 9774 26114 9826 26126
rect 11454 26178 11506 26190
rect 11454 26114 11506 26126
rect 11566 26178 11618 26190
rect 28478 26178 28530 26190
rect 31278 26178 31330 26190
rect 12898 26126 12910 26178
rect 12962 26126 12974 26178
rect 15250 26126 15262 26178
rect 15314 26126 15326 26178
rect 18610 26126 18622 26178
rect 18674 26126 18686 26178
rect 20066 26126 20078 26178
rect 20130 26126 20142 26178
rect 27458 26126 27470 26178
rect 27522 26126 27534 26178
rect 29362 26126 29374 26178
rect 29426 26126 29438 26178
rect 11566 26114 11618 26126
rect 28478 26114 28530 26126
rect 31278 26114 31330 26126
rect 31726 26178 31778 26190
rect 31726 26114 31778 26126
rect 35870 26178 35922 26190
rect 35870 26114 35922 26126
rect 36430 26178 36482 26190
rect 36430 26114 36482 26126
rect 36878 26178 36930 26190
rect 42142 26178 42194 26190
rect 39890 26126 39902 26178
rect 39954 26126 39966 26178
rect 36878 26114 36930 26126
rect 42142 26114 42194 26126
rect 42366 26178 42418 26190
rect 42366 26114 42418 26126
rect 44270 26178 44322 26190
rect 44270 26114 44322 26126
rect 44718 26178 44770 26190
rect 44718 26114 44770 26126
rect 45502 26178 45554 26190
rect 45502 26114 45554 26126
rect 46510 26178 46562 26190
rect 46510 26114 46562 26126
rect 47854 26178 47906 26190
rect 47854 26114 47906 26126
rect 48750 26178 48802 26190
rect 48750 26114 48802 26126
rect 49422 26178 49474 26190
rect 49422 26114 49474 26126
rect 49870 26178 49922 26190
rect 57486 26178 57538 26190
rect 53442 26126 53454 26178
rect 53506 26126 53518 26178
rect 49870 26114 49922 26126
rect 57486 26114 57538 26126
rect 16494 26066 16546 26078
rect 12786 26014 12798 26066
rect 12850 26014 12862 26066
rect 16494 26002 16546 26014
rect 25902 26066 25954 26078
rect 25902 26002 25954 26014
rect 30270 26066 30322 26078
rect 30270 26002 30322 26014
rect 30382 26066 30434 26078
rect 42590 26066 42642 26078
rect 54350 26066 54402 26078
rect 31154 26014 31166 26066
rect 31218 26063 31230 26066
rect 31714 26063 31726 26066
rect 31218 26017 31726 26063
rect 31218 26014 31230 26017
rect 31714 26014 31726 26017
rect 31778 26014 31790 26066
rect 35970 26014 35982 26066
rect 36034 26063 36046 26066
rect 36418 26063 36430 26066
rect 36034 26017 36430 26063
rect 36034 26014 36046 26017
rect 36418 26014 36430 26017
rect 36482 26063 36494 26066
rect 36866 26063 36878 26066
rect 36482 26017 36878 26063
rect 36482 26014 36494 26017
rect 36866 26014 36878 26017
rect 36930 26014 36942 26066
rect 44034 26014 44046 26066
rect 44098 26063 44110 26066
rect 44706 26063 44718 26066
rect 44098 26017 44718 26063
rect 44098 26014 44110 26017
rect 44706 26014 44718 26017
rect 44770 26014 44782 26066
rect 45826 26014 45838 26066
rect 45890 26063 45902 26066
rect 46498 26063 46510 26066
rect 45890 26017 46510 26063
rect 45890 26014 45902 26017
rect 46498 26014 46510 26017
rect 46562 26014 46574 26066
rect 47506 26014 47518 26066
rect 47570 26063 47582 26066
rect 47842 26063 47854 26066
rect 47570 26017 47854 26063
rect 47570 26014 47582 26017
rect 47842 26014 47854 26017
rect 47906 26014 47918 26066
rect 53666 26014 53678 26066
rect 53730 26014 53742 26066
rect 30382 26002 30434 26014
rect 42590 26002 42642 26014
rect 54350 26002 54402 26014
rect 1344 25898 59024 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 59024 25898
rect 1344 25812 59024 25846
rect 22094 25730 22146 25742
rect 43822 25730 43874 25742
rect 8978 25678 8990 25730
rect 9042 25727 9054 25730
rect 9538 25727 9550 25730
rect 9042 25681 9550 25727
rect 9042 25678 9054 25681
rect 9538 25678 9550 25681
rect 9602 25678 9614 25730
rect 22418 25678 22430 25730
rect 22482 25678 22494 25730
rect 22094 25666 22146 25678
rect 43822 25666 43874 25678
rect 2046 25618 2098 25630
rect 2046 25554 2098 25566
rect 2942 25618 2994 25630
rect 5854 25618 5906 25630
rect 8766 25618 8818 25630
rect 4050 25566 4062 25618
rect 4114 25566 4126 25618
rect 6738 25566 6750 25618
rect 6802 25566 6814 25618
rect 7858 25566 7870 25618
rect 7922 25566 7934 25618
rect 2942 25554 2994 25566
rect 5854 25554 5906 25566
rect 8766 25554 8818 25566
rect 9214 25618 9266 25630
rect 9214 25554 9266 25566
rect 9662 25618 9714 25630
rect 9662 25554 9714 25566
rect 11678 25618 11730 25630
rect 11678 25554 11730 25566
rect 13022 25618 13074 25630
rect 13022 25554 13074 25566
rect 13806 25618 13858 25630
rect 13806 25554 13858 25566
rect 14142 25618 14194 25630
rect 16942 25618 16994 25630
rect 21870 25618 21922 25630
rect 15250 25566 15262 25618
rect 15314 25566 15326 25618
rect 19058 25566 19070 25618
rect 19122 25566 19134 25618
rect 20066 25566 20078 25618
rect 20130 25566 20142 25618
rect 14142 25554 14194 25566
rect 16942 25554 16994 25566
rect 21870 25554 21922 25566
rect 22990 25618 23042 25630
rect 22990 25554 23042 25566
rect 23550 25618 23602 25630
rect 26910 25618 26962 25630
rect 26114 25566 26126 25618
rect 26178 25566 26190 25618
rect 23550 25554 23602 25566
rect 26910 25554 26962 25566
rect 33182 25618 33234 25630
rect 36542 25618 36594 25630
rect 33954 25566 33966 25618
rect 34018 25566 34030 25618
rect 33182 25554 33234 25566
rect 36542 25554 36594 25566
rect 37438 25618 37490 25630
rect 37438 25554 37490 25566
rect 38446 25618 38498 25630
rect 38446 25554 38498 25566
rect 38782 25618 38834 25630
rect 38782 25554 38834 25566
rect 39678 25618 39730 25630
rect 41470 25618 41522 25630
rect 43150 25618 43202 25630
rect 51326 25618 51378 25630
rect 41010 25566 41022 25618
rect 41074 25566 41086 25618
rect 42354 25566 42366 25618
rect 42418 25566 42430 25618
rect 48850 25566 48862 25618
rect 48914 25566 48926 25618
rect 54338 25566 54350 25618
rect 54402 25566 54414 25618
rect 55794 25566 55806 25618
rect 55858 25566 55870 25618
rect 57138 25566 57150 25618
rect 57202 25566 57214 25618
rect 39678 25554 39730 25566
rect 41470 25554 41522 25566
rect 43150 25554 43202 25566
rect 51326 25554 51378 25566
rect 10110 25506 10162 25518
rect 6402 25454 6414 25506
rect 6466 25454 6478 25506
rect 10110 25442 10162 25454
rect 10558 25506 10610 25518
rect 10558 25442 10610 25454
rect 11790 25506 11842 25518
rect 11790 25442 11842 25454
rect 12574 25506 12626 25518
rect 32846 25506 32898 25518
rect 43934 25506 43986 25518
rect 50542 25506 50594 25518
rect 15362 25454 15374 25506
rect 15426 25454 15438 25506
rect 18162 25454 18174 25506
rect 18226 25454 18238 25506
rect 18386 25454 18398 25506
rect 18450 25454 18462 25506
rect 24098 25454 24110 25506
rect 24162 25454 24174 25506
rect 24658 25454 24670 25506
rect 24722 25454 24734 25506
rect 27346 25454 27358 25506
rect 27410 25454 27422 25506
rect 32162 25454 32174 25506
rect 32226 25454 32238 25506
rect 34178 25454 34190 25506
rect 34242 25454 34254 25506
rect 40674 25454 40686 25506
rect 40738 25454 40750 25506
rect 42802 25454 42814 25506
rect 42866 25454 42878 25506
rect 45826 25454 45838 25506
rect 45890 25454 45902 25506
rect 46834 25454 46846 25506
rect 46898 25454 46910 25506
rect 47618 25454 47630 25506
rect 47682 25454 47694 25506
rect 49074 25454 49086 25506
rect 49138 25454 49150 25506
rect 12574 25442 12626 25454
rect 32846 25442 32898 25454
rect 43934 25442 43986 25454
rect 50542 25442 50594 25454
rect 50766 25506 50818 25518
rect 56926 25506 56978 25518
rect 53890 25454 53902 25506
rect 53954 25454 53966 25506
rect 55682 25454 55694 25506
rect 55746 25454 55758 25506
rect 57810 25454 57822 25506
rect 57874 25454 57886 25506
rect 50766 25442 50818 25454
rect 56926 25442 56978 25454
rect 10782 25394 10834 25406
rect 4050 25342 4062 25394
rect 4114 25342 4126 25394
rect 10782 25330 10834 25342
rect 11342 25394 11394 25406
rect 30382 25394 30434 25406
rect 34862 25394 34914 25406
rect 16258 25342 16270 25394
rect 16322 25342 16334 25394
rect 28242 25342 28254 25394
rect 28306 25342 28318 25394
rect 32050 25342 32062 25394
rect 32114 25342 32126 25394
rect 11342 25330 11394 25342
rect 30382 25330 30434 25342
rect 34862 25330 34914 25342
rect 35534 25394 35586 25406
rect 35534 25330 35586 25342
rect 37886 25394 37938 25406
rect 37886 25330 37938 25342
rect 45502 25394 45554 25406
rect 49758 25394 49810 25406
rect 47954 25342 47966 25394
rect 48018 25342 48030 25394
rect 45502 25330 45554 25342
rect 49758 25330 49810 25342
rect 50318 25394 50370 25406
rect 50318 25330 50370 25342
rect 50878 25394 50930 25406
rect 50878 25330 50930 25342
rect 53454 25394 53506 25406
rect 53454 25330 53506 25342
rect 56030 25394 56082 25406
rect 56030 25330 56082 25342
rect 2382 25282 2434 25294
rect 2382 25218 2434 25230
rect 4846 25282 4898 25294
rect 4846 25218 4898 25230
rect 7422 25282 7474 25294
rect 7422 25218 7474 25230
rect 10446 25282 10498 25294
rect 10446 25218 10498 25230
rect 11566 25282 11618 25294
rect 11566 25218 11618 25230
rect 11902 25282 11954 25294
rect 11902 25218 11954 25230
rect 20526 25282 20578 25294
rect 20526 25218 20578 25230
rect 29822 25282 29874 25294
rect 29822 25218 29874 25230
rect 31166 25282 31218 25294
rect 31166 25218 31218 25230
rect 35758 25282 35810 25294
rect 35758 25218 35810 25230
rect 35870 25282 35922 25294
rect 35870 25218 35922 25230
rect 35982 25282 36034 25294
rect 35982 25218 36034 25230
rect 39230 25282 39282 25294
rect 39230 25218 39282 25230
rect 44046 25282 44098 25294
rect 44046 25218 44098 25230
rect 44606 25282 44658 25294
rect 44606 25218 44658 25230
rect 45614 25282 45666 25294
rect 46834 25230 46846 25282
rect 46898 25230 46910 25282
rect 47842 25230 47854 25282
rect 47906 25230 47918 25282
rect 45614 25218 45666 25230
rect 1344 25114 59024 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 59024 25114
rect 1344 25028 59024 25062
rect 2270 24946 2322 24958
rect 2270 24882 2322 24894
rect 2718 24946 2770 24958
rect 2718 24882 2770 24894
rect 3726 24946 3778 24958
rect 3726 24882 3778 24894
rect 9886 24946 9938 24958
rect 9886 24882 9938 24894
rect 11902 24946 11954 24958
rect 11902 24882 11954 24894
rect 15710 24946 15762 24958
rect 15710 24882 15762 24894
rect 16606 24946 16658 24958
rect 16606 24882 16658 24894
rect 17054 24946 17106 24958
rect 30382 24946 30434 24958
rect 19842 24894 19854 24946
rect 19906 24894 19918 24946
rect 17054 24882 17106 24894
rect 30382 24882 30434 24894
rect 30830 24946 30882 24958
rect 30830 24882 30882 24894
rect 32062 24946 32114 24958
rect 34862 24946 34914 24958
rect 34738 24894 34750 24946
rect 34802 24894 34814 24946
rect 32062 24882 32114 24894
rect 34862 24882 34914 24894
rect 36094 24946 36146 24958
rect 36094 24882 36146 24894
rect 36654 24946 36706 24958
rect 36654 24882 36706 24894
rect 40014 24946 40066 24958
rect 40014 24882 40066 24894
rect 40462 24946 40514 24958
rect 40462 24882 40514 24894
rect 41470 24946 41522 24958
rect 41470 24882 41522 24894
rect 44382 24946 44434 24958
rect 44382 24882 44434 24894
rect 45054 24946 45106 24958
rect 45054 24882 45106 24894
rect 47742 24946 47794 24958
rect 47742 24882 47794 24894
rect 48414 24946 48466 24958
rect 48414 24882 48466 24894
rect 48638 24946 48690 24958
rect 48638 24882 48690 24894
rect 49982 24946 50034 24958
rect 49982 24882 50034 24894
rect 50094 24946 50146 24958
rect 57474 24894 57486 24946
rect 57538 24894 57550 24946
rect 50094 24882 50146 24894
rect 8878 24834 8930 24846
rect 12238 24834 12290 24846
rect 18734 24834 18786 24846
rect 29486 24834 29538 24846
rect 5730 24782 5742 24834
rect 5794 24782 5806 24834
rect 10434 24782 10446 24834
rect 10498 24782 10510 24834
rect 10994 24782 11006 24834
rect 11058 24782 11070 24834
rect 13234 24782 13246 24834
rect 13298 24782 13310 24834
rect 21970 24782 21982 24834
rect 22034 24782 22046 24834
rect 24434 24782 24446 24834
rect 24498 24782 24510 24834
rect 26338 24782 26350 24834
rect 26402 24782 26414 24834
rect 27570 24782 27582 24834
rect 27634 24782 27646 24834
rect 8878 24770 8930 24782
rect 12238 24770 12290 24782
rect 18734 24770 18786 24782
rect 29486 24770 29538 24782
rect 29934 24834 29986 24846
rect 35870 24834 35922 24846
rect 52782 24834 52834 24846
rect 33954 24782 33966 24834
rect 34018 24782 34030 24834
rect 47170 24782 47182 24834
rect 47234 24782 47246 24834
rect 29934 24770 29986 24782
rect 35870 24770 35922 24782
rect 52782 24770 52834 24782
rect 55582 24834 55634 24846
rect 55582 24770 55634 24782
rect 55694 24834 55746 24846
rect 55694 24770 55746 24782
rect 6974 24722 7026 24734
rect 11566 24722 11618 24734
rect 4722 24670 4734 24722
rect 4786 24670 4798 24722
rect 7074 24670 7086 24722
rect 7138 24670 7150 24722
rect 6974 24658 7026 24670
rect 11566 24658 11618 24670
rect 11902 24722 11954 24734
rect 28366 24722 28418 24734
rect 14130 24670 14142 24722
rect 14194 24670 14206 24722
rect 14690 24670 14702 24722
rect 14754 24670 14766 24722
rect 18050 24670 18062 24722
rect 18114 24670 18126 24722
rect 20850 24670 20862 24722
rect 20914 24670 20926 24722
rect 21410 24670 21422 24722
rect 21474 24670 21486 24722
rect 23090 24670 23102 24722
rect 23154 24670 23166 24722
rect 23762 24670 23774 24722
rect 23826 24670 23838 24722
rect 26226 24670 26238 24722
rect 26290 24670 26302 24722
rect 11902 24658 11954 24670
rect 28366 24658 28418 24670
rect 31278 24722 31330 24734
rect 35646 24722 35698 24734
rect 34178 24670 34190 24722
rect 34242 24670 34254 24722
rect 34514 24670 34526 24722
rect 34578 24670 34590 24722
rect 31278 24658 31330 24670
rect 35646 24658 35698 24670
rect 36318 24722 36370 24734
rect 43038 24722 43090 24734
rect 45390 24722 45442 24734
rect 48750 24722 48802 24734
rect 37426 24670 37438 24722
rect 37490 24670 37502 24722
rect 38770 24670 38782 24722
rect 38834 24670 38846 24722
rect 43250 24670 43262 24722
rect 43314 24670 43326 24722
rect 47058 24670 47070 24722
rect 47122 24670 47134 24722
rect 36318 24658 36370 24670
rect 43038 24658 43090 24670
rect 45390 24658 45442 24670
rect 48750 24658 48802 24670
rect 53006 24722 53058 24734
rect 53006 24658 53058 24670
rect 53342 24722 53394 24734
rect 53342 24658 53394 24670
rect 57822 24722 57874 24734
rect 57822 24658 57874 24670
rect 1934 24610 1986 24622
rect 1934 24546 1986 24558
rect 3166 24610 3218 24622
rect 16158 24610 16210 24622
rect 19294 24610 19346 24622
rect 4946 24558 4958 24610
rect 5010 24558 5022 24610
rect 18386 24558 18398 24610
rect 18450 24558 18462 24610
rect 3166 24546 3218 24558
rect 16158 24546 16210 24558
rect 19294 24546 19346 24558
rect 25790 24610 25842 24622
rect 25790 24546 25842 24558
rect 32510 24610 32562 24622
rect 42366 24610 42418 24622
rect 37314 24558 37326 24610
rect 37378 24558 37390 24610
rect 32510 24546 32562 24558
rect 42366 24546 42418 24558
rect 43934 24610 43986 24622
rect 43934 24546 43986 24558
rect 53230 24610 53282 24622
rect 53230 24546 53282 24558
rect 58046 24610 58098 24622
rect 58046 24546 58098 24558
rect 10222 24498 10274 24510
rect 2034 24446 2046 24498
rect 2098 24495 2110 24498
rect 2706 24495 2718 24498
rect 2098 24449 2718 24495
rect 2098 24446 2110 24449
rect 2706 24446 2718 24449
rect 2770 24495 2782 24498
rect 3266 24495 3278 24498
rect 2770 24449 3278 24495
rect 2770 24446 2782 24449
rect 3266 24446 3278 24449
rect 3330 24446 3342 24498
rect 10222 24434 10274 24446
rect 19518 24498 19570 24510
rect 19518 24434 19570 24446
rect 28590 24498 28642 24510
rect 46062 24498 46114 24510
rect 28914 24446 28926 24498
rect 28978 24446 28990 24498
rect 39442 24446 39454 24498
rect 39506 24446 39518 24498
rect 40002 24446 40014 24498
rect 40066 24495 40078 24498
rect 40450 24495 40462 24498
rect 40066 24449 40462 24495
rect 40066 24446 40078 24449
rect 40450 24446 40462 24449
rect 40514 24446 40526 24498
rect 44146 24446 44158 24498
rect 44210 24495 44222 24498
rect 44818 24495 44830 24498
rect 44210 24449 44830 24495
rect 44210 24446 44222 24449
rect 44818 24446 44830 24449
rect 44882 24446 44894 24498
rect 28590 24434 28642 24446
rect 46062 24434 46114 24446
rect 46398 24498 46450 24510
rect 46398 24434 46450 24446
rect 50206 24498 50258 24510
rect 50206 24434 50258 24446
rect 55582 24498 55634 24510
rect 55582 24434 55634 24446
rect 1344 24330 59024 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 59024 24330
rect 1344 24244 59024 24278
rect 11790 24162 11842 24174
rect 41134 24162 41186 24174
rect 3378 24110 3390 24162
rect 3442 24159 3454 24162
rect 4498 24159 4510 24162
rect 3442 24113 4510 24159
rect 3442 24110 3454 24113
rect 4498 24110 4510 24113
rect 4562 24110 4574 24162
rect 32386 24110 32398 24162
rect 32450 24110 32462 24162
rect 11790 24098 11842 24110
rect 41134 24098 41186 24110
rect 1822 24050 1874 24062
rect 1822 23986 1874 23998
rect 2382 24050 2434 24062
rect 2382 23986 2434 23998
rect 2718 24050 2770 24062
rect 2718 23986 2770 23998
rect 3278 24050 3330 24062
rect 3278 23986 3330 23998
rect 3726 24050 3778 24062
rect 3726 23986 3778 23998
rect 4062 24050 4114 24062
rect 4062 23986 4114 23998
rect 4510 24050 4562 24062
rect 12462 24050 12514 24062
rect 7634 23998 7646 24050
rect 7698 23998 7710 24050
rect 4510 23986 4562 23998
rect 12462 23986 12514 23998
rect 13022 24050 13074 24062
rect 18286 24050 18338 24062
rect 15138 23998 15150 24050
rect 15202 23998 15214 24050
rect 13022 23986 13074 23998
rect 18286 23986 18338 23998
rect 18734 24050 18786 24062
rect 18734 23986 18786 23998
rect 19182 24050 19234 24062
rect 19182 23986 19234 23998
rect 19518 24050 19570 24062
rect 19518 23986 19570 23998
rect 22094 24050 22146 24062
rect 22094 23986 22146 23998
rect 23662 24050 23714 24062
rect 33406 24050 33458 24062
rect 26786 23998 26798 24050
rect 26850 23998 26862 24050
rect 28466 23998 28478 24050
rect 28530 23998 28542 24050
rect 23662 23986 23714 23998
rect 33406 23986 33458 23998
rect 33854 24050 33906 24062
rect 33854 23986 33906 23998
rect 34750 24050 34802 24062
rect 34750 23986 34802 23998
rect 37774 24050 37826 24062
rect 37774 23986 37826 23998
rect 39006 24050 39058 24062
rect 39006 23986 39058 23998
rect 39566 24050 39618 24062
rect 39566 23986 39618 23998
rect 39902 24050 39954 24062
rect 39902 23986 39954 23998
rect 40462 24050 40514 24062
rect 40462 23986 40514 23998
rect 44382 24050 44434 24062
rect 46958 24050 47010 24062
rect 45602 23998 45614 24050
rect 45666 23998 45678 24050
rect 48514 23998 48526 24050
rect 48578 23998 48590 24050
rect 54674 23998 54686 24050
rect 54738 23998 54750 24050
rect 44382 23986 44434 23998
rect 46958 23986 47010 23998
rect 8654 23938 8706 23950
rect 21758 23938 21810 23950
rect 6738 23886 6750 23938
rect 6802 23886 6814 23938
rect 7074 23886 7086 23938
rect 7138 23886 7150 23938
rect 8754 23886 8766 23938
rect 8818 23886 8830 23938
rect 11218 23886 11230 23938
rect 11282 23886 11294 23938
rect 11442 23886 11454 23938
rect 11506 23886 11518 23938
rect 13906 23886 13918 23938
rect 13970 23886 13982 23938
rect 14578 23886 14590 23938
rect 14642 23886 14654 23938
rect 20178 23886 20190 23938
rect 20242 23886 20254 23938
rect 20626 23886 20638 23938
rect 20690 23886 20702 23938
rect 8654 23874 8706 23886
rect 21758 23874 21810 23886
rect 21870 23938 21922 23950
rect 21870 23874 21922 23886
rect 22206 23938 22258 23950
rect 37550 23938 37602 23950
rect 25442 23886 25454 23938
rect 25506 23886 25518 23938
rect 26002 23886 26014 23938
rect 26066 23886 26078 23938
rect 27458 23886 27470 23938
rect 27522 23886 27534 23938
rect 28018 23886 28030 23938
rect 28082 23886 28094 23938
rect 29586 23886 29598 23938
rect 29650 23886 29662 23938
rect 30930 23886 30942 23938
rect 30994 23886 31006 23938
rect 31938 23886 31950 23938
rect 32002 23886 32014 23938
rect 36082 23886 36094 23938
rect 36146 23886 36158 23938
rect 22206 23874 22258 23886
rect 37550 23874 37602 23886
rect 37998 23938 38050 23950
rect 37998 23874 38050 23886
rect 38334 23938 38386 23950
rect 38334 23874 38386 23886
rect 40910 23938 40962 23950
rect 40910 23874 40962 23886
rect 42926 23938 42978 23950
rect 42926 23874 42978 23886
rect 43150 23938 43202 23950
rect 45826 23886 45838 23938
rect 45890 23886 45902 23938
rect 50194 23886 50206 23938
rect 50258 23886 50270 23938
rect 54114 23886 54126 23938
rect 54178 23886 54190 23938
rect 54450 23886 54462 23938
rect 54514 23886 54526 23938
rect 56354 23886 56366 23938
rect 56418 23886 56430 23938
rect 57250 23886 57262 23938
rect 57314 23886 57326 23938
rect 43150 23874 43202 23886
rect 4958 23826 5010 23838
rect 4958 23762 5010 23774
rect 10558 23826 10610 23838
rect 10558 23762 10610 23774
rect 11678 23826 11730 23838
rect 11678 23762 11730 23774
rect 17614 23826 17666 23838
rect 17614 23762 17666 23774
rect 23774 23826 23826 23838
rect 36766 23826 36818 23838
rect 25106 23774 25118 23826
rect 25170 23774 25182 23826
rect 28354 23774 28366 23826
rect 28418 23774 28430 23826
rect 32162 23774 32174 23826
rect 32226 23774 32238 23826
rect 34962 23774 34974 23826
rect 35026 23774 35038 23826
rect 23774 23762 23826 23774
rect 36766 23762 36818 23774
rect 38222 23826 38274 23838
rect 42478 23826 42530 23838
rect 41458 23774 41470 23826
rect 41522 23774 41534 23826
rect 38222 23762 38274 23774
rect 42478 23762 42530 23774
rect 42702 23826 42754 23838
rect 42702 23762 42754 23774
rect 46510 23826 46562 23838
rect 50654 23826 50706 23838
rect 57934 23826 57986 23838
rect 49074 23774 49086 23826
rect 49138 23774 49150 23826
rect 55122 23774 55134 23826
rect 55186 23774 55198 23826
rect 56130 23774 56142 23826
rect 56194 23774 56206 23826
rect 46510 23762 46562 23774
rect 50654 23762 50706 23774
rect 57934 23762 57986 23774
rect 16382 23714 16434 23726
rect 16382 23650 16434 23662
rect 16830 23714 16882 23726
rect 16830 23650 16882 23662
rect 20750 23714 20802 23726
rect 20750 23650 20802 23662
rect 22990 23714 23042 23726
rect 22990 23650 23042 23662
rect 23550 23714 23602 23726
rect 23550 23650 23602 23662
rect 38446 23714 38498 23726
rect 38446 23650 38498 23662
rect 47518 23714 47570 23726
rect 47518 23650 47570 23662
rect 1344 23546 59024 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 59024 23546
rect 1344 23460 59024 23494
rect 2046 23378 2098 23390
rect 2046 23314 2098 23326
rect 2830 23378 2882 23390
rect 2830 23314 2882 23326
rect 3838 23378 3890 23390
rect 3838 23314 3890 23326
rect 5630 23378 5682 23390
rect 5630 23314 5682 23326
rect 5966 23378 6018 23390
rect 5966 23314 6018 23326
rect 9662 23378 9714 23390
rect 9662 23314 9714 23326
rect 11790 23378 11842 23390
rect 11790 23314 11842 23326
rect 12126 23378 12178 23390
rect 12126 23314 12178 23326
rect 13470 23378 13522 23390
rect 13470 23314 13522 23326
rect 14030 23378 14082 23390
rect 14030 23314 14082 23326
rect 14478 23378 14530 23390
rect 14478 23314 14530 23326
rect 14926 23378 14978 23390
rect 14926 23314 14978 23326
rect 17950 23378 18002 23390
rect 17950 23314 18002 23326
rect 19854 23378 19906 23390
rect 30606 23378 30658 23390
rect 26562 23326 26574 23378
rect 26626 23326 26638 23378
rect 19854 23314 19906 23326
rect 30606 23314 30658 23326
rect 32062 23378 32114 23390
rect 32062 23314 32114 23326
rect 32398 23378 32450 23390
rect 32398 23314 32450 23326
rect 33630 23378 33682 23390
rect 39902 23378 39954 23390
rect 36194 23326 36206 23378
rect 36258 23326 36270 23378
rect 33630 23314 33682 23326
rect 39902 23314 39954 23326
rect 40014 23378 40066 23390
rect 40014 23314 40066 23326
rect 46398 23378 46450 23390
rect 46398 23314 46450 23326
rect 55694 23378 55746 23390
rect 55694 23314 55746 23326
rect 56142 23378 56194 23390
rect 56142 23314 56194 23326
rect 4622 23266 4674 23278
rect 4622 23202 4674 23214
rect 5070 23266 5122 23278
rect 5070 23202 5122 23214
rect 8990 23266 9042 23278
rect 8990 23202 9042 23214
rect 10894 23266 10946 23278
rect 10894 23202 10946 23214
rect 12798 23266 12850 23278
rect 12798 23202 12850 23214
rect 18510 23266 18562 23278
rect 18510 23202 18562 23214
rect 22318 23266 22370 23278
rect 22318 23202 22370 23214
rect 24670 23266 24722 23278
rect 24670 23202 24722 23214
rect 24782 23266 24834 23278
rect 32174 23266 32226 23278
rect 26114 23214 26126 23266
rect 26178 23214 26190 23266
rect 24782 23202 24834 23214
rect 32174 23202 32226 23214
rect 35086 23266 35138 23278
rect 35086 23202 35138 23214
rect 36766 23266 36818 23278
rect 36766 23202 36818 23214
rect 36990 23266 37042 23278
rect 51102 23266 51154 23278
rect 37202 23214 37214 23266
rect 37266 23263 37278 23266
rect 37538 23263 37550 23266
rect 37266 23217 37550 23263
rect 37266 23214 37278 23217
rect 37538 23214 37550 23217
rect 37602 23214 37614 23266
rect 36990 23202 37042 23214
rect 51102 23202 51154 23214
rect 51326 23266 51378 23278
rect 51326 23202 51378 23214
rect 11230 23154 11282 23166
rect 6626 23102 6638 23154
rect 6690 23102 6702 23154
rect 8082 23102 8094 23154
rect 8146 23102 8158 23154
rect 11230 23090 11282 23102
rect 12910 23154 12962 23166
rect 12910 23090 12962 23102
rect 15486 23154 15538 23166
rect 17838 23154 17890 23166
rect 30942 23154 30994 23166
rect 31390 23154 31442 23166
rect 34638 23154 34690 23166
rect 16706 23102 16718 23154
rect 16770 23102 16782 23154
rect 16930 23102 16942 23154
rect 16994 23102 17006 23154
rect 21298 23102 21310 23154
rect 21362 23102 21374 23154
rect 26002 23102 26014 23154
rect 26066 23102 26078 23154
rect 27458 23102 27470 23154
rect 27522 23102 27534 23154
rect 30706 23102 30718 23154
rect 30770 23102 30782 23154
rect 31154 23102 31166 23154
rect 31218 23102 31230 23154
rect 32610 23102 32622 23154
rect 32674 23102 32686 23154
rect 15486 23090 15538 23102
rect 17838 23090 17890 23102
rect 30942 23090 30994 23102
rect 31390 23090 31442 23102
rect 34638 23090 34690 23102
rect 34750 23154 34802 23166
rect 34750 23090 34802 23102
rect 35870 23154 35922 23166
rect 40126 23154 40178 23166
rect 38210 23102 38222 23154
rect 38274 23102 38286 23154
rect 39666 23102 39678 23154
rect 39730 23102 39742 23154
rect 35870 23090 35922 23102
rect 40126 23090 40178 23102
rect 40238 23154 40290 23166
rect 40238 23090 40290 23102
rect 41694 23154 41746 23166
rect 42590 23154 42642 23166
rect 42018 23102 42030 23154
rect 42082 23102 42094 23154
rect 41694 23090 41746 23102
rect 42590 23090 42642 23102
rect 43262 23154 43314 23166
rect 44830 23154 44882 23166
rect 50990 23154 51042 23166
rect 53342 23154 53394 23166
rect 43474 23102 43486 23154
rect 43538 23102 43550 23154
rect 45042 23102 45054 23154
rect 45106 23102 45118 23154
rect 47170 23102 47182 23154
rect 47234 23102 47246 23154
rect 52658 23102 52670 23154
rect 52722 23102 52734 23154
rect 54338 23102 54350 23154
rect 54402 23102 54414 23154
rect 43262 23090 43314 23102
rect 44830 23090 44882 23102
rect 50990 23090 51042 23102
rect 53342 23090 53394 23102
rect 2382 23042 2434 23054
rect 2382 22978 2434 22990
rect 3278 23042 3330 23054
rect 3278 22978 3330 22990
rect 4174 23042 4226 23054
rect 10110 23042 10162 23054
rect 6962 22990 6974 23042
rect 7026 22990 7038 23042
rect 8642 22990 8654 23042
rect 8706 22990 8718 23042
rect 4174 22978 4226 22990
rect 10110 22978 10162 22990
rect 16046 23042 16098 23054
rect 16046 22978 16098 22990
rect 18958 23042 19010 23054
rect 18958 22978 19010 22990
rect 19518 23042 19570 23054
rect 19518 22978 19570 22990
rect 20414 23042 20466 23054
rect 23102 23042 23154 23054
rect 20738 22990 20750 23042
rect 20802 22990 20814 23042
rect 20414 22978 20466 22990
rect 23102 22978 23154 22990
rect 23662 23042 23714 23054
rect 33966 23042 34018 23054
rect 29250 22990 29262 23042
rect 29314 22990 29326 23042
rect 32162 22990 32174 23042
rect 32226 22990 32238 23042
rect 23662 22978 23714 22990
rect 33966 22978 34018 22990
rect 35646 23042 35698 23054
rect 38782 23042 38834 23054
rect 37090 22990 37102 23042
rect 37154 22990 37166 23042
rect 38434 22990 38446 23042
rect 38498 22990 38510 23042
rect 35646 22978 35698 22990
rect 38782 22978 38834 22990
rect 40798 23042 40850 23054
rect 40798 22978 40850 22990
rect 44158 23042 44210 23054
rect 44158 22978 44210 22990
rect 45726 23042 45778 23054
rect 47854 23042 47906 23054
rect 47058 22990 47070 23042
rect 47122 22990 47134 23042
rect 45726 22978 45778 22990
rect 47854 22978 47906 22990
rect 48302 23042 48354 23054
rect 48302 22978 48354 22990
rect 53454 23042 53506 23054
rect 54450 22990 54462 23042
rect 54514 22990 54526 23042
rect 53454 22978 53506 22990
rect 12798 22930 12850 22942
rect 1922 22878 1934 22930
rect 1986 22927 1998 22930
rect 2370 22927 2382 22930
rect 1986 22881 2382 22927
rect 1986 22878 1998 22881
rect 2370 22878 2382 22881
rect 2434 22927 2446 22930
rect 2930 22927 2942 22930
rect 2434 22881 2942 22927
rect 2434 22878 2446 22881
rect 2930 22878 2942 22881
rect 2994 22927 3006 22930
rect 3266 22927 3278 22930
rect 2994 22881 3278 22927
rect 2994 22878 3006 22881
rect 3266 22878 3278 22881
rect 3330 22927 3342 22930
rect 4946 22927 4958 22930
rect 3330 22881 4958 22927
rect 3330 22878 3342 22881
rect 4946 22878 4958 22881
rect 5010 22878 5022 22930
rect 11554 22878 11566 22930
rect 11618 22927 11630 22930
rect 11890 22927 11902 22930
rect 11618 22881 11902 22927
rect 11618 22878 11630 22881
rect 11890 22878 11902 22881
rect 11954 22927 11966 22930
rect 12114 22927 12126 22930
rect 11954 22881 12126 22927
rect 11954 22878 11966 22881
rect 12114 22878 12126 22881
rect 12178 22878 12190 22930
rect 12798 22866 12850 22878
rect 17950 22930 18002 22942
rect 17950 22866 18002 22878
rect 24782 22930 24834 22942
rect 24782 22866 24834 22878
rect 34974 22930 35026 22942
rect 54674 22878 54686 22930
rect 54738 22878 54750 22930
rect 34974 22866 35026 22878
rect 1344 22762 59024 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 59024 22762
rect 1344 22676 59024 22710
rect 30158 22594 30210 22606
rect 46734 22594 46786 22606
rect 3490 22542 3502 22594
rect 3554 22591 3566 22594
rect 3714 22591 3726 22594
rect 3554 22545 3726 22591
rect 3554 22542 3566 22545
rect 3714 22542 3726 22545
rect 3778 22542 3790 22594
rect 4386 22542 4398 22594
rect 4450 22591 4462 22594
rect 4946 22591 4958 22594
rect 4450 22545 4958 22591
rect 4450 22542 4462 22545
rect 4946 22542 4958 22545
rect 5010 22542 5022 22594
rect 41122 22542 41134 22594
rect 41186 22591 41198 22594
rect 41906 22591 41918 22594
rect 41186 22545 41918 22591
rect 41186 22542 41198 22545
rect 41906 22542 41918 22545
rect 41970 22542 41982 22594
rect 30158 22530 30210 22542
rect 46734 22530 46786 22542
rect 2158 22482 2210 22494
rect 2158 22418 2210 22430
rect 2606 22482 2658 22494
rect 2606 22418 2658 22430
rect 3502 22482 3554 22494
rect 3502 22418 3554 22430
rect 4062 22482 4114 22494
rect 4062 22418 4114 22430
rect 4398 22482 4450 22494
rect 4398 22418 4450 22430
rect 5966 22482 6018 22494
rect 10222 22482 10274 22494
rect 8194 22430 8206 22482
rect 8258 22430 8270 22482
rect 9538 22430 9550 22482
rect 9602 22430 9614 22482
rect 5966 22418 6018 22430
rect 10222 22418 10274 22430
rect 10670 22482 10722 22494
rect 10670 22418 10722 22430
rect 11566 22482 11618 22494
rect 11566 22418 11618 22430
rect 14814 22482 14866 22494
rect 14814 22418 14866 22430
rect 15598 22482 15650 22494
rect 21646 22482 21698 22494
rect 22542 22482 22594 22494
rect 17266 22430 17278 22482
rect 17330 22430 17342 22482
rect 18722 22430 18734 22482
rect 18786 22430 18798 22482
rect 21970 22430 21982 22482
rect 22034 22430 22046 22482
rect 15598 22418 15650 22430
rect 21646 22418 21698 22430
rect 22542 22418 22594 22430
rect 23550 22482 23602 22494
rect 27358 22482 27410 22494
rect 25778 22430 25790 22482
rect 25842 22430 25854 22482
rect 23550 22418 23602 22430
rect 27358 22418 27410 22430
rect 28478 22482 28530 22494
rect 28478 22418 28530 22430
rect 29710 22482 29762 22494
rect 29710 22418 29762 22430
rect 30382 22482 30434 22494
rect 30382 22418 30434 22430
rect 31614 22482 31666 22494
rect 31614 22418 31666 22430
rect 32286 22482 32338 22494
rect 32286 22418 32338 22430
rect 32622 22482 32674 22494
rect 32622 22418 32674 22430
rect 34862 22482 34914 22494
rect 34862 22418 34914 22430
rect 35646 22482 35698 22494
rect 35646 22418 35698 22430
rect 36094 22482 36146 22494
rect 36094 22418 36146 22430
rect 37438 22482 37490 22494
rect 37438 22418 37490 22430
rect 39342 22482 39394 22494
rect 39342 22418 39394 22430
rect 41918 22482 41970 22494
rect 41918 22418 41970 22430
rect 42814 22482 42866 22494
rect 42814 22418 42866 22430
rect 43262 22482 43314 22494
rect 43262 22418 43314 22430
rect 43934 22482 43986 22494
rect 43934 22418 43986 22430
rect 48190 22482 48242 22494
rect 56354 22430 56366 22482
rect 56418 22430 56430 22482
rect 48190 22418 48242 22430
rect 4846 22370 4898 22382
rect 12798 22370 12850 22382
rect 7858 22318 7870 22370
rect 7922 22318 7934 22370
rect 4846 22306 4898 22318
rect 12798 22306 12850 22318
rect 13918 22370 13970 22382
rect 20190 22370 20242 22382
rect 17042 22318 17054 22370
rect 17106 22318 17118 22370
rect 18386 22318 18398 22370
rect 18450 22318 18462 22370
rect 13918 22306 13970 22318
rect 20190 22306 20242 22318
rect 20862 22370 20914 22382
rect 20862 22306 20914 22318
rect 22990 22370 23042 22382
rect 27582 22370 27634 22382
rect 24210 22318 24222 22370
rect 24274 22318 24286 22370
rect 25890 22318 25902 22370
rect 25954 22318 25966 22370
rect 22990 22306 23042 22318
rect 27582 22306 27634 22318
rect 30606 22370 30658 22382
rect 30606 22306 30658 22318
rect 30830 22370 30882 22382
rect 30830 22306 30882 22318
rect 33518 22370 33570 22382
rect 33966 22370 34018 22382
rect 33842 22318 33854 22370
rect 33906 22318 33918 22370
rect 33518 22306 33570 22318
rect 33966 22306 34018 22318
rect 44494 22370 44546 22382
rect 44494 22306 44546 22318
rect 44830 22370 44882 22382
rect 44830 22306 44882 22318
rect 45502 22370 45554 22382
rect 45502 22306 45554 22318
rect 46062 22370 46114 22382
rect 50530 22318 50542 22370
rect 50594 22318 50606 22370
rect 50978 22318 50990 22370
rect 51042 22318 51054 22370
rect 54002 22318 54014 22370
rect 54066 22318 54078 22370
rect 54450 22318 54462 22370
rect 54514 22318 54526 22370
rect 57250 22318 57262 22370
rect 57314 22318 57326 22370
rect 46062 22306 46114 22318
rect 6414 22258 6466 22270
rect 6414 22194 6466 22206
rect 7422 22258 7474 22270
rect 7422 22194 7474 22206
rect 11118 22258 11170 22270
rect 11118 22194 11170 22206
rect 13806 22258 13858 22270
rect 13806 22194 13858 22206
rect 16382 22258 16434 22270
rect 16382 22194 16434 22206
rect 17950 22258 18002 22270
rect 40126 22258 40178 22270
rect 24770 22206 24782 22258
rect 24834 22206 24846 22258
rect 27906 22206 27918 22258
rect 27970 22206 27982 22258
rect 17950 22194 18002 22206
rect 40126 22194 40178 22206
rect 40574 22258 40626 22270
rect 40574 22194 40626 22206
rect 47742 22258 47794 22270
rect 47742 22194 47794 22206
rect 51214 22258 51266 22270
rect 51214 22194 51266 22206
rect 51774 22258 51826 22270
rect 51774 22194 51826 22206
rect 51998 22258 52050 22270
rect 51998 22194 52050 22206
rect 52222 22258 52274 22270
rect 52222 22194 52274 22206
rect 52334 22258 52386 22270
rect 55122 22206 55134 22258
rect 55186 22206 55198 22258
rect 56018 22206 56030 22258
rect 56082 22206 56094 22258
rect 52334 22194 52386 22206
rect 1822 22146 1874 22158
rect 1822 22082 1874 22094
rect 3054 22146 3106 22158
rect 3054 22082 3106 22094
rect 6862 22146 6914 22158
rect 6862 22082 6914 22094
rect 9102 22146 9154 22158
rect 9102 22082 9154 22094
rect 12126 22146 12178 22158
rect 12126 22082 12178 22094
rect 12238 22146 12290 22158
rect 12238 22082 12290 22094
rect 12350 22146 12402 22158
rect 12350 22082 12402 22094
rect 13582 22146 13634 22158
rect 13582 22082 13634 22094
rect 15150 22146 15202 22158
rect 15150 22082 15202 22094
rect 19518 22146 19570 22158
rect 19518 22082 19570 22094
rect 19630 22146 19682 22158
rect 19630 22082 19682 22094
rect 19742 22146 19794 22158
rect 19742 22082 19794 22094
rect 20526 22146 20578 22158
rect 20526 22082 20578 22094
rect 20750 22146 20802 22158
rect 20750 22082 20802 22094
rect 23438 22146 23490 22158
rect 23438 22082 23490 22094
rect 23662 22146 23714 22158
rect 23662 22082 23714 22094
rect 28814 22146 28866 22158
rect 28814 22082 28866 22094
rect 30718 22146 30770 22158
rect 30718 22082 30770 22094
rect 34078 22146 34130 22158
rect 34078 22082 34130 22094
rect 34190 22146 34242 22158
rect 34190 22082 34242 22094
rect 35198 22146 35250 22158
rect 35198 22082 35250 22094
rect 36542 22146 36594 22158
rect 36542 22082 36594 22094
rect 37886 22146 37938 22158
rect 37886 22082 37938 22094
rect 38334 22146 38386 22158
rect 38334 22082 38386 22094
rect 38782 22146 38834 22158
rect 38782 22082 38834 22094
rect 40350 22146 40402 22158
rect 40350 22082 40402 22094
rect 40686 22146 40738 22158
rect 40686 22082 40738 22094
rect 41022 22146 41074 22158
rect 41022 22082 41074 22094
rect 41470 22146 41522 22158
rect 41470 22082 41522 22094
rect 42366 22146 42418 22158
rect 42366 22082 42418 22094
rect 44606 22146 44658 22158
rect 44606 22082 44658 22094
rect 45950 22146 46002 22158
rect 45950 22082 46002 22094
rect 46174 22146 46226 22158
rect 46174 22082 46226 22094
rect 46846 22146 46898 22158
rect 46846 22082 46898 22094
rect 46958 22146 47010 22158
rect 46958 22082 47010 22094
rect 47630 22146 47682 22158
rect 47630 22082 47682 22094
rect 48638 22146 48690 22158
rect 48638 22082 48690 22094
rect 58158 22146 58210 22158
rect 58158 22082 58210 22094
rect 1344 21978 59024 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 59024 21978
rect 1344 21892 59024 21926
rect 2158 21810 2210 21822
rect 2158 21746 2210 21758
rect 2718 21810 2770 21822
rect 2718 21746 2770 21758
rect 3502 21810 3554 21822
rect 3502 21746 3554 21758
rect 5406 21810 5458 21822
rect 5406 21746 5458 21758
rect 7310 21810 7362 21822
rect 7310 21746 7362 21758
rect 8990 21810 9042 21822
rect 8990 21746 9042 21758
rect 9998 21810 10050 21822
rect 9998 21746 10050 21758
rect 11454 21810 11506 21822
rect 11454 21746 11506 21758
rect 14478 21810 14530 21822
rect 14478 21746 14530 21758
rect 17838 21810 17890 21822
rect 17838 21746 17890 21758
rect 17950 21810 18002 21822
rect 17950 21746 18002 21758
rect 18622 21810 18674 21822
rect 18622 21746 18674 21758
rect 25678 21810 25730 21822
rect 25678 21746 25730 21758
rect 29150 21810 29202 21822
rect 29150 21746 29202 21758
rect 29486 21810 29538 21822
rect 29486 21746 29538 21758
rect 30382 21810 30434 21822
rect 30382 21746 30434 21758
rect 30830 21810 30882 21822
rect 30830 21746 30882 21758
rect 34862 21810 34914 21822
rect 34862 21746 34914 21758
rect 35310 21810 35362 21822
rect 35310 21746 35362 21758
rect 37214 21810 37266 21822
rect 37214 21746 37266 21758
rect 37774 21810 37826 21822
rect 37774 21746 37826 21758
rect 38222 21810 38274 21822
rect 38222 21746 38274 21758
rect 40574 21810 40626 21822
rect 40574 21746 40626 21758
rect 43374 21810 43426 21822
rect 43374 21746 43426 21758
rect 47406 21810 47458 21822
rect 51650 21758 51662 21810
rect 51714 21758 51726 21810
rect 54114 21758 54126 21810
rect 54178 21758 54190 21810
rect 47406 21746 47458 21758
rect 1822 21698 1874 21710
rect 1822 21634 1874 21646
rect 5854 21698 5906 21710
rect 5854 21634 5906 21646
rect 6190 21698 6242 21710
rect 10558 21698 10610 21710
rect 7970 21646 7982 21698
rect 8034 21646 8046 21698
rect 6190 21634 6242 21646
rect 10558 21634 10610 21646
rect 16606 21698 16658 21710
rect 16606 21634 16658 21646
rect 16942 21698 16994 21710
rect 16942 21634 16994 21646
rect 20526 21698 20578 21710
rect 20526 21634 20578 21646
rect 23102 21698 23154 21710
rect 23102 21634 23154 21646
rect 24558 21698 24610 21710
rect 24558 21634 24610 21646
rect 28926 21698 28978 21710
rect 28926 21634 28978 21646
rect 30606 21698 30658 21710
rect 30606 21634 30658 21646
rect 32510 21698 32562 21710
rect 32510 21634 32562 21646
rect 32734 21698 32786 21710
rect 32734 21634 32786 21646
rect 36318 21698 36370 21710
rect 36318 21634 36370 21646
rect 43486 21698 43538 21710
rect 48302 21698 48354 21710
rect 45042 21646 45054 21698
rect 45106 21646 45118 21698
rect 43486 21634 43538 21646
rect 48302 21634 48354 21646
rect 48414 21698 48466 21710
rect 48414 21634 48466 21646
rect 50542 21698 50594 21710
rect 50542 21634 50594 21646
rect 53566 21698 53618 21710
rect 53566 21634 53618 21646
rect 3054 21586 3106 21598
rect 3054 21522 3106 21534
rect 4846 21586 4898 21598
rect 4846 21522 4898 21534
rect 6638 21586 6690 21598
rect 10334 21586 10386 21598
rect 7858 21534 7870 21586
rect 7922 21534 7934 21586
rect 6638 21522 6690 21534
rect 10334 21522 10386 21534
rect 10670 21586 10722 21598
rect 10670 21522 10722 21534
rect 12238 21586 12290 21598
rect 15822 21586 15874 21598
rect 12898 21534 12910 21586
rect 12962 21534 12974 21586
rect 13234 21534 13246 21586
rect 13298 21534 13310 21586
rect 15586 21534 15598 21586
rect 15650 21534 15662 21586
rect 12238 21522 12290 21534
rect 15822 21522 15874 21534
rect 18062 21586 18114 21598
rect 18062 21522 18114 21534
rect 18846 21586 18898 21598
rect 18846 21522 18898 21534
rect 19294 21586 19346 21598
rect 24446 21586 24498 21598
rect 20066 21534 20078 21586
rect 20130 21534 20142 21586
rect 20290 21534 20302 21586
rect 20354 21534 20366 21586
rect 21298 21534 21310 21586
rect 21362 21534 21374 21586
rect 22194 21534 22206 21586
rect 22258 21534 22270 21586
rect 19294 21522 19346 21534
rect 24446 21522 24498 21534
rect 24670 21586 24722 21598
rect 29374 21586 29426 21598
rect 35870 21586 35922 21598
rect 26338 21534 26350 21586
rect 26402 21534 26414 21586
rect 26674 21534 26686 21586
rect 26738 21534 26750 21586
rect 33842 21534 33854 21586
rect 33906 21534 33918 21586
rect 24670 21522 24722 21534
rect 29374 21522 29426 21534
rect 35870 21522 35922 21534
rect 36094 21586 36146 21598
rect 36094 21522 36146 21534
rect 36542 21586 36594 21598
rect 36542 21522 36594 21534
rect 37102 21586 37154 21598
rect 37102 21522 37154 21534
rect 37438 21586 37490 21598
rect 39790 21586 39842 21598
rect 39218 21534 39230 21586
rect 39282 21534 39294 21586
rect 37438 21522 37490 21534
rect 39790 21522 39842 21534
rect 41470 21586 41522 21598
rect 41470 21522 41522 21534
rect 43150 21586 43202 21598
rect 45726 21586 45778 21598
rect 47182 21586 47234 21598
rect 43810 21534 43822 21586
rect 43874 21534 43886 21586
rect 45938 21534 45950 21586
rect 46002 21534 46014 21586
rect 43150 21522 43202 21534
rect 45726 21522 45778 21534
rect 47182 21522 47234 21534
rect 47294 21586 47346 21598
rect 47294 21522 47346 21534
rect 47854 21586 47906 21598
rect 47854 21522 47906 21534
rect 49646 21586 49698 21598
rect 51102 21586 51154 21598
rect 49858 21534 49870 21586
rect 49922 21534 49934 21586
rect 49646 21522 49698 21534
rect 51102 21522 51154 21534
rect 53790 21586 53842 21598
rect 53790 21522 53842 21534
rect 55358 21586 55410 21598
rect 55358 21522 55410 21534
rect 57486 21586 57538 21598
rect 57486 21522 57538 21534
rect 57710 21586 57762 21598
rect 58494 21586 58546 21598
rect 58034 21534 58046 21586
rect 58098 21534 58110 21586
rect 57710 21522 57762 21534
rect 58494 21522 58546 21534
rect 3950 21474 4002 21486
rect 3950 21410 4002 21422
rect 4398 21474 4450 21486
rect 11790 21474 11842 21486
rect 14926 21474 14978 21486
rect 8530 21422 8542 21474
rect 8594 21422 8606 21474
rect 12562 21422 12574 21474
rect 12626 21422 12638 21474
rect 4398 21410 4450 21422
rect 11790 21410 11842 21422
rect 14926 21410 14978 21422
rect 18734 21474 18786 21486
rect 18734 21410 18786 21422
rect 22318 21474 22370 21486
rect 28366 21474 28418 21486
rect 23538 21422 23550 21474
rect 23602 21422 23614 21474
rect 27794 21422 27806 21474
rect 27858 21422 27870 21474
rect 22318 21410 22370 21422
rect 28366 21410 28418 21422
rect 29262 21474 29314 21486
rect 29262 21410 29314 21422
rect 30494 21474 30546 21486
rect 30494 21410 30546 21422
rect 31614 21474 31666 21486
rect 34414 21474 34466 21486
rect 32834 21422 32846 21474
rect 32898 21422 32910 21474
rect 33954 21422 33966 21474
rect 34018 21422 34030 21474
rect 31614 21410 31666 21422
rect 34414 21410 34466 21422
rect 36654 21474 36706 21486
rect 36654 21410 36706 21422
rect 41918 21474 41970 21486
rect 41918 21410 41970 21422
rect 42590 21474 42642 21486
rect 44494 21474 44546 21486
rect 43922 21422 43934 21474
rect 43986 21422 43998 21474
rect 42590 21410 42642 21422
rect 44494 21410 44546 21422
rect 44718 21474 44770 21486
rect 44718 21410 44770 21422
rect 46622 21474 46674 21486
rect 52110 21474 52162 21486
rect 47842 21422 47854 21474
rect 47906 21471 47918 21474
rect 48066 21471 48078 21474
rect 47906 21425 48078 21471
rect 47906 21422 47918 21425
rect 48066 21422 48078 21425
rect 48130 21422 48142 21474
rect 46622 21410 46674 21422
rect 52110 21410 52162 21422
rect 55582 21474 55634 21486
rect 55582 21410 55634 21422
rect 56702 21474 56754 21486
rect 56702 21410 56754 21422
rect 57598 21474 57650 21486
rect 57598 21410 57650 21422
rect 20638 21362 20690 21374
rect 38894 21362 38946 21374
rect 3490 21310 3502 21362
rect 3554 21359 3566 21362
rect 4162 21359 4174 21362
rect 3554 21313 4174 21359
rect 3554 21310 3566 21313
rect 4162 21310 4174 21313
rect 4226 21310 4238 21362
rect 11778 21310 11790 21362
rect 11842 21359 11854 21362
rect 12002 21359 12014 21362
rect 11842 21313 12014 21359
rect 11842 21310 11854 21313
rect 12002 21310 12014 21313
rect 12066 21310 12078 21362
rect 22194 21310 22206 21362
rect 22258 21310 22270 21362
rect 20638 21298 20690 21310
rect 38894 21298 38946 21310
rect 39230 21362 39282 21374
rect 39230 21298 39282 21310
rect 48414 21362 48466 21374
rect 48414 21298 48466 21310
rect 51326 21362 51378 21374
rect 56142 21362 56194 21374
rect 55010 21310 55022 21362
rect 55074 21310 55086 21362
rect 51326 21298 51378 21310
rect 56142 21298 56194 21310
rect 56478 21362 56530 21374
rect 56478 21298 56530 21310
rect 1344 21194 59024 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 59024 21194
rect 1344 21108 59024 21142
rect 12910 21026 12962 21038
rect 3938 20974 3950 21026
rect 4002 21023 4014 21026
rect 4498 21023 4510 21026
rect 4002 20977 4510 21023
rect 4002 20974 4014 20977
rect 4498 20974 4510 20977
rect 4562 20974 4574 21026
rect 12910 20962 12962 20974
rect 13694 21026 13746 21038
rect 13694 20962 13746 20974
rect 21870 21026 21922 21038
rect 21870 20962 21922 20974
rect 23326 21026 23378 21038
rect 31614 21026 31666 21038
rect 30930 20974 30942 21026
rect 30994 20974 31006 21026
rect 23326 20962 23378 20974
rect 31614 20962 31666 20974
rect 31950 21026 32002 21038
rect 40686 21026 40738 21038
rect 34738 20974 34750 21026
rect 34802 20974 34814 21026
rect 39106 20974 39118 21026
rect 39170 21023 39182 21026
rect 39890 21023 39902 21026
rect 39170 20977 39902 21023
rect 39170 20974 39182 20977
rect 39890 20974 39902 20977
rect 39954 20974 39966 21026
rect 31950 20962 32002 20974
rect 40686 20962 40738 20974
rect 2270 20914 2322 20926
rect 2270 20850 2322 20862
rect 2718 20914 2770 20926
rect 2718 20850 2770 20862
rect 3166 20914 3218 20926
rect 3166 20850 3218 20862
rect 4062 20914 4114 20926
rect 4062 20850 4114 20862
rect 4510 20914 4562 20926
rect 4510 20850 4562 20862
rect 4958 20914 5010 20926
rect 4958 20850 5010 20862
rect 5630 20914 5682 20926
rect 5630 20850 5682 20862
rect 6078 20914 6130 20926
rect 15822 20914 15874 20926
rect 7522 20862 7534 20914
rect 7586 20862 7598 20914
rect 9762 20862 9774 20914
rect 9826 20862 9838 20914
rect 6078 20850 6130 20862
rect 15822 20850 15874 20862
rect 17166 20914 17218 20926
rect 17166 20850 17218 20862
rect 18062 20914 18114 20926
rect 18062 20850 18114 20862
rect 19070 20914 19122 20926
rect 25902 20914 25954 20926
rect 20178 20862 20190 20914
rect 20242 20862 20254 20914
rect 24322 20862 24334 20914
rect 24386 20862 24398 20914
rect 19070 20850 19122 20862
rect 25902 20850 25954 20862
rect 26574 20914 26626 20926
rect 26574 20850 26626 20862
rect 26686 20914 26738 20926
rect 36766 20914 36818 20926
rect 36082 20862 36094 20914
rect 36146 20862 36158 20914
rect 26686 20850 26738 20862
rect 36766 20850 36818 20862
rect 39902 20914 39954 20926
rect 39902 20850 39954 20862
rect 43038 20914 43090 20926
rect 43038 20850 43090 20862
rect 45726 20914 45778 20926
rect 49310 20914 49362 20926
rect 46386 20862 46398 20914
rect 46450 20862 46462 20914
rect 50530 20862 50542 20914
rect 50594 20862 50606 20914
rect 57362 20862 57374 20914
rect 57426 20862 57438 20914
rect 45726 20850 45778 20862
rect 49310 20850 49362 20862
rect 11790 20802 11842 20814
rect 7298 20750 7310 20802
rect 7362 20750 7374 20802
rect 9426 20750 9438 20802
rect 9490 20750 9502 20802
rect 11790 20738 11842 20750
rect 15150 20802 15202 20814
rect 17726 20802 17778 20814
rect 21758 20802 21810 20814
rect 16482 20750 16494 20802
rect 16546 20750 16558 20802
rect 19506 20750 19518 20802
rect 19570 20750 19582 20802
rect 15150 20738 15202 20750
rect 17726 20738 17778 20750
rect 21758 20738 21810 20750
rect 22094 20802 22146 20814
rect 22094 20738 22146 20750
rect 26910 20802 26962 20814
rect 27806 20802 27858 20814
rect 27346 20750 27358 20802
rect 27410 20750 27422 20802
rect 26910 20738 26962 20750
rect 27806 20738 27858 20750
rect 28366 20802 28418 20814
rect 28366 20738 28418 20750
rect 28590 20802 28642 20814
rect 32510 20802 32562 20814
rect 34078 20802 34130 20814
rect 35758 20802 35810 20814
rect 37886 20802 37938 20814
rect 30258 20750 30270 20802
rect 30322 20750 30334 20802
rect 32946 20750 32958 20802
rect 33010 20750 33022 20802
rect 33618 20750 33630 20802
rect 33682 20750 33694 20802
rect 34178 20750 34190 20802
rect 34242 20750 34254 20802
rect 35522 20750 35534 20802
rect 35586 20750 35598 20802
rect 37538 20750 37550 20802
rect 37602 20750 37614 20802
rect 28590 20738 28642 20750
rect 32510 20738 32562 20750
rect 34078 20738 34130 20750
rect 35758 20738 35810 20750
rect 37886 20738 37938 20750
rect 38110 20802 38162 20814
rect 42366 20802 42418 20814
rect 41010 20750 41022 20802
rect 41074 20750 41086 20802
rect 42018 20750 42030 20802
rect 42082 20750 42094 20802
rect 38110 20738 38162 20750
rect 42366 20738 42418 20750
rect 42590 20802 42642 20814
rect 54350 20802 54402 20814
rect 46498 20750 46510 20802
rect 46562 20750 46574 20802
rect 47842 20750 47854 20802
rect 47906 20750 47918 20802
rect 50866 20750 50878 20802
rect 50930 20750 50942 20802
rect 56354 20750 56366 20802
rect 56418 20750 56430 20802
rect 57250 20750 57262 20802
rect 57314 20750 57326 20802
rect 42590 20738 42642 20750
rect 54350 20738 54402 20750
rect 6638 20690 6690 20702
rect 6638 20626 6690 20638
rect 8990 20690 9042 20702
rect 12798 20690 12850 20702
rect 10882 20638 10894 20690
rect 10946 20638 10958 20690
rect 11554 20638 11566 20690
rect 11618 20638 11630 20690
rect 8990 20626 9042 20638
rect 12798 20626 12850 20638
rect 13918 20690 13970 20702
rect 23214 20690 23266 20702
rect 22642 20638 22654 20690
rect 22706 20638 22718 20690
rect 13918 20626 13970 20638
rect 23214 20626 23266 20638
rect 23998 20690 24050 20702
rect 23998 20626 24050 20638
rect 25006 20690 25058 20702
rect 25006 20626 25058 20638
rect 26462 20690 26514 20702
rect 28814 20690 28866 20702
rect 40462 20690 40514 20702
rect 27122 20638 27134 20690
rect 27186 20638 27198 20690
rect 28130 20638 28142 20690
rect 28194 20638 28206 20690
rect 29810 20638 29822 20690
rect 29874 20638 29886 20690
rect 26462 20626 26514 20638
rect 28814 20626 28866 20638
rect 40462 20626 40514 20638
rect 48638 20690 48690 20702
rect 48638 20626 48690 20638
rect 51326 20690 51378 20702
rect 51326 20626 51378 20638
rect 54686 20690 54738 20702
rect 56702 20690 56754 20702
rect 56018 20638 56030 20690
rect 56082 20638 56094 20690
rect 54686 20626 54738 20638
rect 56702 20626 56754 20638
rect 1934 20578 1986 20590
rect 1934 20514 1986 20526
rect 3614 20578 3666 20590
rect 3614 20514 3666 20526
rect 8430 20578 8482 20590
rect 12238 20578 12290 20590
rect 11666 20526 11678 20578
rect 11730 20526 11742 20578
rect 8430 20514 8482 20526
rect 12238 20514 12290 20526
rect 13806 20578 13858 20590
rect 13806 20514 13858 20526
rect 14814 20578 14866 20590
rect 14814 20514 14866 20526
rect 16270 20578 16322 20590
rect 16270 20514 16322 20526
rect 18510 20578 18562 20590
rect 18510 20514 18562 20526
rect 23326 20578 23378 20590
rect 23326 20514 23378 20526
rect 24222 20578 24274 20590
rect 24222 20514 24274 20526
rect 25454 20578 25506 20590
rect 25454 20514 25506 20526
rect 28366 20578 28418 20590
rect 28366 20514 28418 20526
rect 31838 20578 31890 20590
rect 31838 20514 31890 20526
rect 35982 20578 36034 20590
rect 35982 20514 36034 20526
rect 36094 20578 36146 20590
rect 36094 20514 36146 20526
rect 37998 20578 38050 20590
rect 37998 20514 38050 20526
rect 38558 20578 38610 20590
rect 38558 20514 38610 20526
rect 39006 20578 39058 20590
rect 39006 20514 39058 20526
rect 39454 20578 39506 20590
rect 39454 20514 39506 20526
rect 42478 20578 42530 20590
rect 42478 20514 42530 20526
rect 53790 20578 53842 20590
rect 53790 20514 53842 20526
rect 54462 20578 54514 20590
rect 54462 20514 54514 20526
rect 1344 20410 59024 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 59024 20410
rect 1344 20324 59024 20358
rect 2718 20242 2770 20254
rect 2718 20178 2770 20190
rect 5294 20242 5346 20254
rect 5294 20178 5346 20190
rect 5854 20242 5906 20254
rect 5854 20178 5906 20190
rect 7870 20242 7922 20254
rect 7870 20178 7922 20190
rect 17838 20242 17890 20254
rect 17838 20178 17890 20190
rect 20526 20242 20578 20254
rect 20526 20178 20578 20190
rect 21422 20242 21474 20254
rect 21422 20178 21474 20190
rect 23662 20242 23714 20254
rect 23662 20178 23714 20190
rect 23886 20242 23938 20254
rect 23886 20178 23938 20190
rect 24446 20242 24498 20254
rect 31838 20242 31890 20254
rect 30818 20190 30830 20242
rect 30882 20190 30894 20242
rect 24446 20178 24498 20190
rect 31838 20178 31890 20190
rect 40014 20242 40066 20254
rect 40014 20178 40066 20190
rect 40910 20242 40962 20254
rect 40910 20178 40962 20190
rect 46062 20242 46114 20254
rect 46062 20178 46114 20190
rect 47854 20242 47906 20254
rect 47854 20178 47906 20190
rect 48302 20242 48354 20254
rect 48302 20178 48354 20190
rect 56478 20242 56530 20254
rect 56478 20178 56530 20190
rect 4510 20130 4562 20142
rect 4510 20066 4562 20078
rect 4958 20130 5010 20142
rect 4958 20066 5010 20078
rect 6190 20130 6242 20142
rect 6190 20066 6242 20078
rect 11678 20130 11730 20142
rect 11678 20066 11730 20078
rect 14478 20130 14530 20142
rect 14478 20066 14530 20078
rect 18286 20130 18338 20142
rect 18286 20066 18338 20078
rect 18846 20130 18898 20142
rect 18846 20066 18898 20078
rect 21310 20130 21362 20142
rect 21310 20066 21362 20078
rect 21646 20130 21698 20142
rect 21646 20066 21698 20078
rect 22094 20130 22146 20142
rect 22094 20066 22146 20078
rect 23550 20130 23602 20142
rect 23550 20066 23602 20078
rect 25006 20130 25058 20142
rect 25006 20066 25058 20078
rect 27246 20130 27298 20142
rect 27246 20066 27298 20078
rect 27806 20130 27858 20142
rect 27806 20066 27858 20078
rect 28030 20130 28082 20142
rect 32062 20130 32114 20142
rect 30146 20078 30158 20130
rect 30210 20078 30222 20130
rect 28030 20066 28082 20078
rect 32062 20066 32114 20078
rect 32734 20130 32786 20142
rect 32734 20066 32786 20078
rect 35870 20130 35922 20142
rect 35870 20066 35922 20078
rect 36542 20130 36594 20142
rect 36542 20066 36594 20078
rect 36766 20130 36818 20142
rect 56590 20130 56642 20142
rect 37538 20078 37550 20130
rect 37602 20078 37614 20130
rect 39106 20078 39118 20130
rect 39170 20078 39182 20130
rect 53442 20078 53454 20130
rect 53506 20078 53518 20130
rect 54786 20078 54798 20130
rect 54850 20078 54862 20130
rect 36766 20066 36818 20078
rect 56590 20066 56642 20078
rect 57486 20130 57538 20142
rect 57486 20066 57538 20078
rect 3054 20018 3106 20030
rect 3054 19954 3106 19966
rect 3502 20018 3554 20030
rect 3502 19954 3554 19966
rect 7086 20018 7138 20030
rect 7086 19954 7138 19966
rect 7198 20018 7250 20030
rect 7198 19954 7250 19966
rect 7646 20018 7698 20030
rect 12014 20018 12066 20030
rect 10658 19966 10670 20018
rect 10722 19966 10734 20018
rect 7646 19954 7698 19966
rect 12014 19954 12066 19966
rect 12574 20018 12626 20030
rect 16494 20018 16546 20030
rect 13234 19966 13246 20018
rect 13298 19966 13310 20018
rect 12574 19954 12626 19966
rect 16494 19954 16546 19966
rect 19742 20018 19794 20030
rect 19742 19954 19794 19966
rect 28702 20018 28754 20030
rect 28702 19954 28754 19966
rect 28926 20018 28978 20030
rect 31726 20018 31778 20030
rect 36430 20018 36482 20030
rect 56254 20018 56306 20030
rect 57822 20018 57874 20030
rect 29810 19966 29822 20018
rect 29874 19966 29886 20018
rect 30930 19966 30942 20018
rect 30994 19966 31006 20018
rect 33842 19966 33854 20018
rect 33906 19966 33918 20018
rect 34850 19966 34862 20018
rect 34914 19966 34926 20018
rect 42242 19966 42254 20018
rect 42306 19966 42318 20018
rect 56018 19966 56030 20018
rect 56082 19966 56094 20018
rect 57586 19966 57598 20018
rect 57650 19966 57662 20018
rect 28926 19954 28978 19966
rect 31726 19954 31778 19966
rect 36430 19954 36482 19966
rect 56254 19954 56306 19966
rect 57822 19954 57874 19966
rect 1822 19906 1874 19918
rect 1822 19842 1874 19854
rect 2270 19906 2322 19918
rect 2270 19842 2322 19854
rect 3950 19906 4002 19918
rect 3950 19842 4002 19854
rect 6862 19906 6914 19918
rect 6862 19842 6914 19854
rect 8206 19906 8258 19918
rect 8206 19842 8258 19854
rect 8990 19906 9042 19918
rect 8990 19842 9042 19854
rect 9998 19906 10050 19918
rect 15262 19906 15314 19918
rect 10770 19854 10782 19906
rect 10834 19854 10846 19906
rect 13346 19854 13358 19906
rect 13410 19854 13422 19906
rect 9998 19842 10050 19854
rect 15262 19842 15314 19854
rect 15598 19906 15650 19918
rect 15598 19842 15650 19854
rect 16046 19906 16098 19918
rect 16046 19842 16098 19854
rect 17054 19906 17106 19918
rect 17054 19842 17106 19854
rect 19182 19906 19234 19918
rect 19182 19842 19234 19854
rect 23102 19906 23154 19918
rect 23102 19842 23154 19854
rect 25678 19906 25730 19918
rect 26462 19906 26514 19918
rect 37438 19906 37490 19918
rect 26002 19854 26014 19906
rect 26066 19854 26078 19906
rect 28130 19854 28142 19906
rect 28194 19854 28206 19906
rect 32834 19854 32846 19906
rect 32898 19854 32910 19906
rect 34178 19854 34190 19906
rect 34242 19854 34254 19906
rect 34626 19854 34638 19906
rect 34690 19854 34702 19906
rect 25678 19842 25730 19854
rect 26462 19842 26514 19854
rect 37438 19842 37490 19854
rect 39454 19906 39506 19918
rect 39454 19842 39506 19854
rect 40350 19906 40402 19918
rect 42926 19906 42978 19918
rect 42466 19854 42478 19906
rect 42530 19854 42542 19906
rect 40350 19842 40402 19854
rect 42926 19842 42978 19854
rect 52222 19906 52274 19918
rect 55022 19906 55074 19918
rect 52882 19854 52894 19906
rect 52946 19854 52958 19906
rect 52222 19842 52274 19854
rect 55022 19842 55074 19854
rect 55470 19906 55522 19918
rect 56578 19854 56590 19906
rect 56642 19854 56654 19906
rect 55470 19842 55522 19854
rect 22206 19794 22258 19806
rect 32510 19794 32562 19806
rect 16034 19742 16046 19794
rect 16098 19791 16110 19794
rect 16706 19791 16718 19794
rect 16098 19745 16718 19791
rect 16098 19742 16110 19745
rect 16706 19742 16718 19745
rect 16770 19742 16782 19794
rect 29250 19742 29262 19794
rect 29314 19742 29326 19794
rect 34962 19742 34974 19794
rect 35026 19742 35038 19794
rect 22206 19730 22258 19742
rect 32510 19730 32562 19742
rect 1344 19626 59024 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 59024 19626
rect 1344 19540 59024 19574
rect 19070 19458 19122 19470
rect 46062 19458 46114 19470
rect 6850 19406 6862 19458
rect 6914 19455 6926 19458
rect 7410 19455 7422 19458
rect 6914 19409 7422 19455
rect 6914 19406 6926 19409
rect 7410 19406 7422 19409
rect 7474 19406 7486 19458
rect 12786 19406 12798 19458
rect 12850 19455 12862 19458
rect 13122 19455 13134 19458
rect 12850 19409 13134 19455
rect 12850 19406 12862 19409
rect 13122 19406 13134 19409
rect 13186 19406 13198 19458
rect 19282 19406 19294 19458
rect 19346 19455 19358 19458
rect 20514 19455 20526 19458
rect 19346 19409 20526 19455
rect 19346 19406 19358 19409
rect 20514 19406 20526 19409
rect 20578 19455 20590 19458
rect 20850 19455 20862 19458
rect 20578 19409 20862 19455
rect 20578 19406 20590 19409
rect 20850 19406 20862 19409
rect 20914 19406 20926 19458
rect 30370 19406 30382 19458
rect 30434 19455 30446 19458
rect 30706 19455 30718 19458
rect 30434 19409 30718 19455
rect 30434 19406 30446 19409
rect 30706 19406 30718 19409
rect 30770 19406 30782 19458
rect 33842 19406 33854 19458
rect 33906 19455 33918 19458
rect 34066 19455 34078 19458
rect 33906 19409 34078 19455
rect 33906 19406 33918 19409
rect 34066 19406 34078 19409
rect 34130 19455 34142 19458
rect 34850 19455 34862 19458
rect 34130 19409 34862 19455
rect 34130 19406 34142 19409
rect 34850 19406 34862 19409
rect 34914 19406 34926 19458
rect 39106 19455 39118 19458
rect 38673 19409 39118 19455
rect 19070 19394 19122 19406
rect 2382 19346 2434 19358
rect 2382 19282 2434 19294
rect 5070 19346 5122 19358
rect 5070 19282 5122 19294
rect 5854 19346 5906 19358
rect 5854 19282 5906 19294
rect 6302 19346 6354 19358
rect 6302 19282 6354 19294
rect 6750 19346 6802 19358
rect 6750 19282 6802 19294
rect 7086 19346 7138 19358
rect 7086 19282 7138 19294
rect 7534 19346 7586 19358
rect 7534 19282 7586 19294
rect 7982 19346 8034 19358
rect 7982 19282 8034 19294
rect 8990 19346 9042 19358
rect 8990 19282 9042 19294
rect 10558 19346 10610 19358
rect 10558 19282 10610 19294
rect 11006 19346 11058 19358
rect 11006 19282 11058 19294
rect 11454 19346 11506 19358
rect 11454 19282 11506 19294
rect 12126 19346 12178 19358
rect 12126 19282 12178 19294
rect 12574 19346 12626 19358
rect 12574 19282 12626 19294
rect 14366 19346 14418 19358
rect 14366 19282 14418 19294
rect 19406 19346 19458 19358
rect 19406 19282 19458 19294
rect 20414 19346 20466 19358
rect 20414 19282 20466 19294
rect 23774 19346 23826 19358
rect 27134 19346 27186 19358
rect 26450 19294 26462 19346
rect 26514 19294 26526 19346
rect 23774 19282 23826 19294
rect 27134 19282 27186 19294
rect 27582 19346 27634 19358
rect 27582 19282 27634 19294
rect 28366 19346 28418 19358
rect 28366 19282 28418 19294
rect 28814 19346 28866 19358
rect 28814 19282 28866 19294
rect 30382 19346 30434 19358
rect 30382 19282 30434 19294
rect 31166 19346 31218 19358
rect 31166 19282 31218 19294
rect 32958 19346 33010 19358
rect 32958 19282 33010 19294
rect 33406 19346 33458 19358
rect 33406 19282 33458 19294
rect 33854 19346 33906 19358
rect 33854 19282 33906 19294
rect 34302 19346 34354 19358
rect 34302 19282 34354 19294
rect 34750 19346 34802 19358
rect 38446 19346 38498 19358
rect 35746 19294 35758 19346
rect 35810 19294 35822 19346
rect 34750 19282 34802 19294
rect 38446 19282 38498 19294
rect 9886 19234 9938 19246
rect 9886 19170 9938 19182
rect 15374 19234 15426 19246
rect 22318 19234 22370 19246
rect 16034 19182 16046 19234
rect 16098 19182 16110 19234
rect 15374 19170 15426 19182
rect 22318 19170 22370 19182
rect 23102 19234 23154 19246
rect 32622 19234 32674 19246
rect 37886 19234 37938 19246
rect 38673 19234 38719 19409
rect 39106 19406 39118 19409
rect 39170 19406 39182 19458
rect 46062 19394 46114 19406
rect 38782 19346 38834 19358
rect 38782 19282 38834 19294
rect 39342 19346 39394 19358
rect 39342 19282 39394 19294
rect 40910 19346 40962 19358
rect 46398 19346 46450 19358
rect 42914 19294 42926 19346
rect 42978 19294 42990 19346
rect 40910 19282 40962 19294
rect 46398 19282 46450 19294
rect 41470 19234 41522 19246
rect 24994 19182 25006 19234
rect 25058 19182 25070 19234
rect 36194 19182 36206 19234
rect 36258 19182 36270 19234
rect 38658 19182 38670 19234
rect 38722 19182 38734 19234
rect 23102 19170 23154 19182
rect 32622 19170 32674 19182
rect 37886 19170 37938 19182
rect 41470 19170 41522 19182
rect 41806 19234 41858 19246
rect 44046 19234 44098 19246
rect 42578 19182 42590 19234
rect 42642 19182 42654 19234
rect 41806 19170 41858 19182
rect 44046 19170 44098 19182
rect 46846 19234 46898 19246
rect 46846 19170 46898 19182
rect 49086 19234 49138 19246
rect 49086 19170 49138 19182
rect 49422 19234 49474 19246
rect 49422 19170 49474 19182
rect 49870 19234 49922 19246
rect 49870 19170 49922 19182
rect 53678 19234 53730 19246
rect 53678 19170 53730 19182
rect 54350 19234 54402 19246
rect 55458 19182 55470 19234
rect 55522 19182 55534 19234
rect 57922 19182 57934 19234
rect 57986 19182 57998 19234
rect 58370 19182 58382 19234
rect 58434 19182 58446 19234
rect 54350 19170 54402 19182
rect 22094 19122 22146 19134
rect 22094 19058 22146 19070
rect 22990 19122 23042 19134
rect 22990 19058 23042 19070
rect 24334 19122 24386 19134
rect 36654 19122 36706 19134
rect 26114 19070 26126 19122
rect 26178 19070 26190 19122
rect 24334 19058 24386 19070
rect 36654 19058 36706 19070
rect 41582 19122 41634 19134
rect 41582 19058 41634 19070
rect 43486 19122 43538 19134
rect 43486 19058 43538 19070
rect 44158 19122 44210 19134
rect 44158 19058 44210 19070
rect 44718 19122 44770 19134
rect 44718 19058 44770 19070
rect 45838 19122 45890 19134
rect 45838 19058 45890 19070
rect 47406 19122 47458 19134
rect 47406 19058 47458 19070
rect 49198 19122 49250 19134
rect 49198 19058 49250 19070
rect 51326 19122 51378 19134
rect 51326 19058 51378 19070
rect 52670 19122 52722 19134
rect 52670 19058 52722 19070
rect 53902 19122 53954 19134
rect 55346 19070 55358 19122
rect 55410 19070 55422 19122
rect 53902 19058 53954 19070
rect 2718 19010 2770 19022
rect 2718 18946 2770 18958
rect 3166 19010 3218 19022
rect 3166 18946 3218 18958
rect 3614 19010 3666 19022
rect 3614 18946 3666 18958
rect 4062 19010 4114 19022
rect 4062 18946 4114 18958
rect 4510 19010 4562 19022
rect 4510 18946 4562 18958
rect 8430 19010 8482 19022
rect 8430 18946 8482 18958
rect 9550 19010 9602 19022
rect 9550 18946 9602 18958
rect 12910 19010 12962 19022
rect 12910 18946 12962 18958
rect 13582 19010 13634 19022
rect 13582 18946 13634 18958
rect 14702 19010 14754 19022
rect 19966 19010 20018 19022
rect 18274 18958 18286 19010
rect 18338 18958 18350 19010
rect 14702 18946 14754 18958
rect 19966 18946 20018 18958
rect 20862 19010 20914 19022
rect 20862 18946 20914 18958
rect 22206 19010 22258 19022
rect 22206 18946 22258 18958
rect 22766 19010 22818 19022
rect 22766 18946 22818 18958
rect 27918 19010 27970 19022
rect 27918 18946 27970 18958
rect 29486 19010 29538 19022
rect 29486 18946 29538 18958
rect 30718 19010 30770 19022
rect 30718 18946 30770 18958
rect 31614 19010 31666 19022
rect 31614 18946 31666 18958
rect 32062 19010 32114 19022
rect 32062 18946 32114 18958
rect 37438 19010 37490 19022
rect 37438 18946 37490 18958
rect 40238 19010 40290 19022
rect 40238 18946 40290 18958
rect 44382 19010 44434 19022
rect 44382 18946 44434 18958
rect 47294 19010 47346 19022
rect 47294 18946 47346 18958
rect 47518 19010 47570 19022
rect 47518 18946 47570 18958
rect 50318 19010 50370 19022
rect 50318 18946 50370 18958
rect 50430 19010 50482 19022
rect 50430 18946 50482 18958
rect 50542 19010 50594 19022
rect 50542 18946 50594 18958
rect 51438 19010 51490 19022
rect 51438 18946 51490 18958
rect 51662 19010 51714 19022
rect 51662 18946 51714 18958
rect 54126 19010 54178 19022
rect 56018 18958 56030 19010
rect 56082 18958 56094 19010
rect 54126 18946 54178 18958
rect 1344 18842 59024 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 59024 18842
rect 1344 18756 59024 18790
rect 4174 18674 4226 18686
rect 4174 18610 4226 18622
rect 10558 18674 10610 18686
rect 10558 18610 10610 18622
rect 11342 18674 11394 18686
rect 11342 18610 11394 18622
rect 17054 18674 17106 18686
rect 25678 18674 25730 18686
rect 21074 18622 21086 18674
rect 21138 18622 21150 18674
rect 17054 18610 17106 18622
rect 25678 18610 25730 18622
rect 27022 18674 27074 18686
rect 27022 18610 27074 18622
rect 27806 18674 27858 18686
rect 27806 18610 27858 18622
rect 33518 18674 33570 18686
rect 33518 18610 33570 18622
rect 35310 18674 35362 18686
rect 35310 18610 35362 18622
rect 37438 18674 37490 18686
rect 37438 18610 37490 18622
rect 39678 18674 39730 18686
rect 39678 18610 39730 18622
rect 40910 18674 40962 18686
rect 40910 18610 40962 18622
rect 42926 18674 42978 18686
rect 42926 18610 42978 18622
rect 43486 18674 43538 18686
rect 43486 18610 43538 18622
rect 57598 18674 57650 18686
rect 57598 18610 57650 18622
rect 57710 18674 57762 18686
rect 57710 18610 57762 18622
rect 3726 18562 3778 18574
rect 3726 18498 3778 18510
rect 7982 18562 8034 18574
rect 7982 18498 8034 18510
rect 16270 18562 16322 18574
rect 23550 18562 23602 18574
rect 22642 18510 22654 18562
rect 22706 18510 22718 18562
rect 16270 18498 16322 18510
rect 23550 18498 23602 18510
rect 23886 18562 23938 18574
rect 23886 18498 23938 18510
rect 25902 18562 25954 18574
rect 25902 18498 25954 18510
rect 26910 18562 26962 18574
rect 26910 18498 26962 18510
rect 27918 18562 27970 18574
rect 27918 18498 27970 18510
rect 29598 18562 29650 18574
rect 30158 18562 30210 18574
rect 34414 18562 34466 18574
rect 29810 18510 29822 18562
rect 29874 18510 29886 18562
rect 32162 18510 32174 18562
rect 32226 18510 32238 18562
rect 29598 18498 29650 18510
rect 30158 18498 30210 18510
rect 34414 18498 34466 18510
rect 34750 18562 34802 18574
rect 34750 18498 34802 18510
rect 38782 18562 38834 18574
rect 38782 18498 38834 18510
rect 39006 18562 39058 18574
rect 39006 18498 39058 18510
rect 41582 18562 41634 18574
rect 57822 18562 57874 18574
rect 52770 18510 52782 18562
rect 52834 18510 52846 18562
rect 54002 18510 54014 18562
rect 54066 18510 54078 18562
rect 41582 18498 41634 18510
rect 57822 18498 57874 18510
rect 3390 18450 3442 18462
rect 3390 18386 3442 18398
rect 5070 18450 5122 18462
rect 8766 18450 8818 18462
rect 5730 18398 5742 18450
rect 5794 18398 5806 18450
rect 5070 18386 5122 18398
rect 8766 18386 8818 18398
rect 10110 18450 10162 18462
rect 10110 18386 10162 18398
rect 12126 18450 12178 18462
rect 12126 18386 12178 18398
rect 12574 18450 12626 18462
rect 12574 18386 12626 18398
rect 13582 18450 13634 18462
rect 17838 18450 17890 18462
rect 24782 18450 24834 18462
rect 14018 18398 14030 18450
rect 14082 18398 14094 18450
rect 21298 18398 21310 18450
rect 21362 18398 21374 18450
rect 24546 18398 24558 18450
rect 24610 18398 24622 18450
rect 13582 18386 13634 18398
rect 17838 18386 17890 18398
rect 24782 18386 24834 18398
rect 24894 18450 24946 18462
rect 24894 18386 24946 18398
rect 26350 18450 26402 18462
rect 26350 18386 26402 18398
rect 27582 18450 27634 18462
rect 27582 18386 27634 18398
rect 28366 18450 28418 18462
rect 28366 18386 28418 18398
rect 31502 18450 31554 18462
rect 34190 18450 34242 18462
rect 32274 18398 32286 18450
rect 32338 18398 32350 18450
rect 31502 18386 31554 18398
rect 34190 18386 34242 18398
rect 36094 18450 36146 18462
rect 36094 18386 36146 18398
rect 37102 18450 37154 18462
rect 37102 18386 37154 18398
rect 38558 18450 38610 18462
rect 38558 18386 38610 18398
rect 39118 18450 39170 18462
rect 39118 18386 39170 18398
rect 40238 18450 40290 18462
rect 40238 18386 40290 18398
rect 43598 18450 43650 18462
rect 43598 18386 43650 18398
rect 43710 18450 43762 18462
rect 43710 18386 43762 18398
rect 44158 18450 44210 18462
rect 46510 18450 46562 18462
rect 45602 18398 45614 18450
rect 45666 18398 45678 18450
rect 44158 18386 44210 18398
rect 46510 18386 46562 18398
rect 47854 18450 47906 18462
rect 48066 18398 48078 18450
rect 48130 18398 48142 18450
rect 49970 18398 49982 18450
rect 50034 18398 50046 18450
rect 51650 18398 51662 18450
rect 51714 18398 51726 18450
rect 52098 18398 52110 18450
rect 52162 18398 52174 18450
rect 54898 18398 54910 18450
rect 54962 18398 54974 18450
rect 57922 18398 57934 18450
rect 57986 18398 57998 18450
rect 47854 18386 47906 18398
rect 4622 18338 4674 18350
rect 4622 18274 4674 18286
rect 11678 18338 11730 18350
rect 11678 18274 11730 18286
rect 18398 18338 18450 18350
rect 18398 18274 18450 18286
rect 18734 18338 18786 18350
rect 18734 18274 18786 18286
rect 19182 18338 19234 18350
rect 19182 18274 19234 18286
rect 19630 18338 19682 18350
rect 19630 18274 19682 18286
rect 20078 18338 20130 18350
rect 25790 18338 25842 18350
rect 22866 18286 22878 18338
rect 22930 18286 22942 18338
rect 20078 18274 20130 18286
rect 25790 18274 25842 18286
rect 28814 18338 28866 18350
rect 30382 18338 30434 18350
rect 29474 18286 29486 18338
rect 29538 18286 29550 18338
rect 28814 18274 28866 18286
rect 30382 18274 30434 18286
rect 31054 18338 31106 18350
rect 34638 18338 34690 18350
rect 32722 18286 32734 18338
rect 32786 18286 32798 18338
rect 31054 18274 31106 18286
rect 34638 18274 34690 18286
rect 35758 18338 35810 18350
rect 35758 18274 35810 18286
rect 36542 18338 36594 18350
rect 36542 18274 36594 18286
rect 37886 18338 37938 18350
rect 37886 18274 37938 18286
rect 44494 18338 44546 18350
rect 48750 18338 48802 18350
rect 46050 18286 46062 18338
rect 46114 18286 46126 18338
rect 50082 18286 50094 18338
rect 50146 18286 50158 18338
rect 52210 18286 52222 18338
rect 52274 18286 52286 18338
rect 53442 18286 53454 18338
rect 53506 18286 53518 18338
rect 56018 18286 56030 18338
rect 56082 18286 56094 18338
rect 44494 18274 44546 18286
rect 48750 18274 48802 18286
rect 27134 18226 27186 18238
rect 11106 18174 11118 18226
rect 11170 18223 11182 18226
rect 11330 18223 11342 18226
rect 11170 18177 11342 18223
rect 11170 18174 11182 18177
rect 11330 18174 11342 18177
rect 11394 18223 11406 18226
rect 11666 18223 11678 18226
rect 11394 18177 11678 18223
rect 11394 18174 11406 18177
rect 11666 18174 11678 18177
rect 11730 18174 11742 18226
rect 17714 18174 17726 18226
rect 17778 18223 17790 18226
rect 18498 18223 18510 18226
rect 17778 18177 18510 18223
rect 17778 18174 17790 18177
rect 18498 18174 18510 18177
rect 18562 18174 18574 18226
rect 18722 18174 18734 18226
rect 18786 18223 18798 18226
rect 20178 18223 20190 18226
rect 18786 18177 20190 18223
rect 18786 18174 18798 18177
rect 20178 18174 20190 18177
rect 20242 18174 20254 18226
rect 27134 18162 27186 18174
rect 30494 18226 30546 18238
rect 41806 18226 41858 18238
rect 34962 18174 34974 18226
rect 35026 18223 35038 18226
rect 36530 18223 36542 18226
rect 35026 18177 36542 18223
rect 35026 18174 35038 18177
rect 36530 18174 36542 18177
rect 36594 18174 36606 18226
rect 30494 18162 30546 18174
rect 41806 18162 41858 18174
rect 42142 18226 42194 18238
rect 58270 18226 58322 18238
rect 50306 18174 50318 18226
rect 50370 18174 50382 18226
rect 42142 18162 42194 18174
rect 58270 18162 58322 18174
rect 1344 18058 59024 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 59024 18058
rect 1344 17972 59024 18006
rect 13022 17890 13074 17902
rect 22990 17890 23042 17902
rect 30830 17890 30882 17902
rect 13570 17838 13582 17890
rect 13634 17887 13646 17890
rect 15362 17887 15374 17890
rect 13634 17841 15374 17887
rect 13634 17838 13646 17841
rect 15362 17838 15374 17841
rect 15426 17838 15438 17890
rect 23762 17838 23774 17890
rect 23826 17887 23838 17890
rect 24434 17887 24446 17890
rect 23826 17841 24446 17887
rect 23826 17838 23838 17841
rect 24434 17838 24446 17841
rect 24498 17838 24510 17890
rect 27570 17838 27582 17890
rect 27634 17887 27646 17890
rect 28018 17887 28030 17890
rect 27634 17841 28030 17887
rect 27634 17838 27646 17841
rect 28018 17838 28030 17841
rect 28082 17838 28094 17890
rect 13022 17826 13074 17838
rect 22990 17826 23042 17838
rect 30830 17826 30882 17838
rect 33070 17890 33122 17902
rect 33070 17826 33122 17838
rect 37662 17890 37714 17902
rect 37662 17826 37714 17838
rect 37998 17890 38050 17902
rect 37998 17826 38050 17838
rect 48974 17890 49026 17902
rect 48974 17826 49026 17838
rect 50094 17890 50146 17902
rect 50094 17826 50146 17838
rect 4062 17778 4114 17790
rect 4062 17714 4114 17726
rect 4510 17778 4562 17790
rect 4510 17714 4562 17726
rect 4958 17778 5010 17790
rect 4958 17714 5010 17726
rect 5742 17778 5794 17790
rect 5742 17714 5794 17726
rect 6526 17778 6578 17790
rect 6526 17714 6578 17726
rect 7086 17778 7138 17790
rect 7086 17714 7138 17726
rect 7870 17778 7922 17790
rect 7870 17714 7922 17726
rect 8430 17778 8482 17790
rect 8430 17714 8482 17726
rect 14142 17778 14194 17790
rect 14142 17714 14194 17726
rect 19630 17778 19682 17790
rect 19630 17714 19682 17726
rect 19966 17778 20018 17790
rect 19966 17714 20018 17726
rect 20526 17778 20578 17790
rect 20526 17714 20578 17726
rect 20974 17778 21026 17790
rect 20974 17714 21026 17726
rect 23774 17778 23826 17790
rect 23774 17714 23826 17726
rect 24894 17778 24946 17790
rect 24894 17714 24946 17726
rect 25342 17778 25394 17790
rect 25342 17714 25394 17726
rect 26574 17778 26626 17790
rect 26574 17714 26626 17726
rect 27582 17778 27634 17790
rect 27582 17714 27634 17726
rect 28590 17778 28642 17790
rect 40910 17778 40962 17790
rect 38882 17726 38894 17778
rect 38946 17726 38958 17778
rect 28590 17714 28642 17726
rect 40910 17714 40962 17726
rect 41358 17778 41410 17790
rect 44494 17778 44546 17790
rect 49982 17778 50034 17790
rect 53454 17778 53506 17790
rect 43810 17726 43822 17778
rect 43874 17726 43886 17778
rect 46610 17726 46622 17778
rect 46674 17726 46686 17778
rect 51314 17726 51326 17778
rect 51378 17726 51390 17778
rect 41358 17714 41410 17726
rect 44494 17714 44546 17726
rect 49982 17714 50034 17726
rect 53454 17714 53506 17726
rect 53790 17778 53842 17790
rect 53790 17714 53842 17726
rect 9550 17666 9602 17678
rect 13582 17666 13634 17678
rect 9874 17614 9886 17666
rect 9938 17614 9950 17666
rect 9550 17602 9602 17614
rect 13582 17602 13634 17614
rect 15486 17666 15538 17678
rect 19182 17666 19234 17678
rect 16146 17614 16158 17666
rect 16210 17614 16222 17666
rect 15486 17602 15538 17614
rect 19182 17602 19234 17614
rect 22094 17666 22146 17678
rect 22094 17602 22146 17614
rect 22542 17666 22594 17678
rect 22542 17602 22594 17614
rect 23102 17666 23154 17678
rect 23102 17602 23154 17614
rect 24446 17666 24498 17678
rect 24446 17602 24498 17614
rect 25678 17666 25730 17678
rect 25678 17602 25730 17614
rect 26350 17666 26402 17678
rect 26350 17602 26402 17614
rect 26686 17666 26738 17678
rect 26686 17602 26738 17614
rect 33406 17666 33458 17678
rect 33406 17602 33458 17614
rect 34190 17666 34242 17678
rect 35870 17666 35922 17678
rect 34514 17614 34526 17666
rect 34578 17614 34590 17666
rect 34190 17602 34242 17614
rect 35870 17602 35922 17614
rect 36094 17666 36146 17678
rect 40238 17666 40290 17678
rect 36306 17614 36318 17666
rect 36370 17614 36382 17666
rect 38770 17614 38782 17666
rect 38834 17614 38846 17666
rect 36094 17602 36146 17614
rect 40238 17602 40290 17614
rect 42590 17666 42642 17678
rect 48862 17666 48914 17678
rect 51998 17666 52050 17678
rect 42802 17614 42814 17666
rect 42866 17614 42878 17666
rect 43698 17614 43710 17666
rect 43762 17614 43774 17666
rect 46498 17614 46510 17666
rect 46562 17614 46574 17666
rect 51426 17614 51438 17666
rect 51490 17614 51502 17666
rect 55458 17614 55470 17666
rect 55522 17614 55534 17666
rect 57026 17614 57038 17666
rect 57090 17614 57102 17666
rect 57362 17614 57374 17666
rect 57426 17614 57438 17666
rect 42590 17602 42642 17614
rect 48862 17602 48914 17614
rect 51998 17602 52050 17614
rect 25902 17554 25954 17566
rect 25902 17490 25954 17502
rect 27022 17554 27074 17566
rect 35086 17554 35138 17566
rect 30034 17502 30046 17554
rect 30098 17502 30110 17554
rect 30594 17502 30606 17554
rect 30658 17502 30670 17554
rect 32274 17502 32286 17554
rect 32338 17502 32350 17554
rect 32722 17502 32734 17554
rect 32786 17502 32798 17554
rect 27022 17490 27074 17502
rect 35086 17490 35138 17502
rect 35646 17554 35698 17566
rect 35646 17490 35698 17502
rect 36766 17554 36818 17566
rect 36766 17490 36818 17502
rect 39678 17554 39730 17566
rect 39678 17490 39730 17502
rect 42926 17554 42978 17566
rect 42926 17490 42978 17502
rect 47406 17554 47458 17566
rect 47406 17490 47458 17502
rect 48974 17554 49026 17566
rect 55682 17502 55694 17554
rect 55746 17502 55758 17554
rect 48974 17490 49026 17502
rect 6078 17442 6130 17454
rect 6078 17378 6130 17390
rect 7422 17442 7474 17454
rect 7422 17378 7474 17390
rect 8990 17442 9042 17454
rect 14590 17442 14642 17454
rect 12226 17390 12238 17442
rect 12290 17390 12302 17442
rect 8990 17378 9042 17390
rect 14590 17378 14642 17390
rect 15038 17442 15090 17454
rect 21870 17442 21922 17454
rect 18498 17390 18510 17442
rect 18562 17390 18574 17442
rect 15038 17378 15090 17390
rect 21870 17378 21922 17390
rect 21982 17442 22034 17454
rect 21982 17378 22034 17390
rect 28142 17442 28194 17454
rect 28142 17378 28194 17390
rect 28702 17442 28754 17454
rect 28702 17378 28754 17390
rect 31166 17442 31218 17454
rect 31166 17378 31218 17390
rect 35982 17442 36034 17454
rect 35982 17378 36034 17390
rect 37886 17442 37938 17454
rect 37886 17378 37938 17390
rect 40350 17442 40402 17454
rect 40350 17378 40402 17390
rect 40574 17442 40626 17454
rect 56914 17390 56926 17442
rect 56978 17390 56990 17442
rect 40574 17378 40626 17390
rect 1344 17274 59024 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 59024 17274
rect 1344 17188 59024 17222
rect 4622 17106 4674 17118
rect 4622 17042 4674 17054
rect 5070 17106 5122 17118
rect 9102 17106 9154 17118
rect 8530 17054 8542 17106
rect 8594 17054 8606 17106
rect 5070 17042 5122 17054
rect 9102 17042 9154 17054
rect 9774 17106 9826 17118
rect 9774 17042 9826 17054
rect 10222 17106 10274 17118
rect 10222 17042 10274 17054
rect 10670 17106 10722 17118
rect 15710 17106 15762 17118
rect 12114 17054 12126 17106
rect 12178 17054 12190 17106
rect 10670 17042 10722 17054
rect 15710 17042 15762 17054
rect 16158 17106 16210 17118
rect 16158 17042 16210 17054
rect 16606 17106 16658 17118
rect 16606 17042 16658 17054
rect 17726 17106 17778 17118
rect 17726 17042 17778 17054
rect 18062 17106 18114 17118
rect 18062 17042 18114 17054
rect 19182 17106 19234 17118
rect 19182 17042 19234 17054
rect 19854 17106 19906 17118
rect 19854 17042 19906 17054
rect 20526 17106 20578 17118
rect 20526 17042 20578 17054
rect 20974 17106 21026 17118
rect 20974 17042 21026 17054
rect 21422 17106 21474 17118
rect 21422 17042 21474 17054
rect 22990 17106 23042 17118
rect 22990 17042 23042 17054
rect 23550 17106 23602 17118
rect 23550 17042 23602 17054
rect 23998 17106 24050 17118
rect 23998 17042 24050 17054
rect 25006 17106 25058 17118
rect 25006 17042 25058 17054
rect 26238 17106 26290 17118
rect 26238 17042 26290 17054
rect 28366 17106 28418 17118
rect 28366 17042 28418 17054
rect 29374 17106 29426 17118
rect 29374 17042 29426 17054
rect 29934 17106 29986 17118
rect 29934 17042 29986 17054
rect 30046 17106 30098 17118
rect 30046 17042 30098 17054
rect 31054 17106 31106 17118
rect 31054 17042 31106 17054
rect 31390 17106 31442 17118
rect 31390 17042 31442 17054
rect 31838 17106 31890 17118
rect 31838 17042 31890 17054
rect 32734 17106 32786 17118
rect 32734 17042 32786 17054
rect 33854 17106 33906 17118
rect 33854 17042 33906 17054
rect 34078 17106 34130 17118
rect 34078 17042 34130 17054
rect 34750 17106 34802 17118
rect 34750 17042 34802 17054
rect 38894 17106 38946 17118
rect 38894 17042 38946 17054
rect 39566 17106 39618 17118
rect 39566 17042 39618 17054
rect 40350 17106 40402 17118
rect 40350 17042 40402 17054
rect 40574 17106 40626 17118
rect 40574 17042 40626 17054
rect 41470 17106 41522 17118
rect 41470 17042 41522 17054
rect 41918 17106 41970 17118
rect 41918 17042 41970 17054
rect 43038 17106 43090 17118
rect 43038 17042 43090 17054
rect 43150 17106 43202 17118
rect 43150 17042 43202 17054
rect 43262 17106 43314 17118
rect 43262 17042 43314 17054
rect 44382 17106 44434 17118
rect 44382 17042 44434 17054
rect 45166 17106 45218 17118
rect 45166 17042 45218 17054
rect 45614 17106 45666 17118
rect 45614 17042 45666 17054
rect 53790 17106 53842 17118
rect 53790 17042 53842 17054
rect 58270 17106 58322 17118
rect 58270 17042 58322 17054
rect 17054 16994 17106 17006
rect 17054 16930 17106 16942
rect 18846 16994 18898 17006
rect 18846 16930 18898 16942
rect 21870 16994 21922 17006
rect 21870 16930 21922 16942
rect 22206 16994 22258 17006
rect 22206 16930 22258 16942
rect 24446 16994 24498 17006
rect 24446 16930 24498 16942
rect 32622 16994 32674 17006
rect 32622 16930 32674 16942
rect 34190 16994 34242 17006
rect 34190 16930 34242 16942
rect 35646 16994 35698 17006
rect 35646 16930 35698 16942
rect 36542 16994 36594 17006
rect 36542 16930 36594 16942
rect 38334 16994 38386 17006
rect 38334 16930 38386 16942
rect 40126 16994 40178 17006
rect 40126 16930 40178 16942
rect 44718 16994 44770 17006
rect 44718 16930 44770 16942
rect 53902 16994 53954 17006
rect 57822 16994 57874 17006
rect 58382 16994 58434 17006
rect 56354 16942 56366 16994
rect 56418 16942 56430 16994
rect 58146 16942 58158 16994
rect 58210 16942 58222 16994
rect 53902 16930 53954 16942
rect 57822 16930 57874 16942
rect 58382 16930 58434 16942
rect 5406 16882 5458 16894
rect 11230 16882 11282 16894
rect 15038 16882 15090 16894
rect 5954 16830 5966 16882
rect 6018 16830 6030 16882
rect 14466 16830 14478 16882
rect 14530 16830 14542 16882
rect 5406 16818 5458 16830
rect 11230 16818 11282 16830
rect 15038 16818 15090 16830
rect 26686 16882 26738 16894
rect 28702 16882 28754 16894
rect 27234 16830 27246 16882
rect 27298 16830 27310 16882
rect 26686 16818 26738 16830
rect 28702 16818 28754 16830
rect 30158 16882 30210 16894
rect 30158 16818 30210 16830
rect 30606 16882 30658 16894
rect 30606 16818 30658 16830
rect 32958 16882 33010 16894
rect 32958 16818 33010 16830
rect 33742 16882 33794 16894
rect 35534 16882 35586 16894
rect 35298 16830 35310 16882
rect 35362 16830 35374 16882
rect 33742 16818 33794 16830
rect 35534 16818 35586 16830
rect 37438 16882 37490 16894
rect 42814 16882 42866 16894
rect 37874 16830 37886 16882
rect 37938 16830 37950 16882
rect 37438 16818 37490 16830
rect 42814 16818 42866 16830
rect 42926 16882 42978 16894
rect 42926 16818 42978 16830
rect 43822 16882 43874 16894
rect 51998 16882 52050 16894
rect 53342 16882 53394 16894
rect 50082 16830 50094 16882
rect 50146 16830 50158 16882
rect 52322 16830 52334 16882
rect 52386 16830 52398 16882
rect 43822 16818 43874 16830
rect 51998 16818 52050 16830
rect 53342 16818 53394 16830
rect 54014 16882 54066 16894
rect 55234 16830 55246 16882
rect 55298 16830 55310 16882
rect 55570 16830 55582 16882
rect 55634 16830 55646 16882
rect 56242 16830 56254 16882
rect 56306 16830 56318 16882
rect 54014 16818 54066 16830
rect 25678 16770 25730 16782
rect 50766 16770 50818 16782
rect 27458 16718 27470 16770
rect 27522 16718 27534 16770
rect 30594 16718 30606 16770
rect 30658 16718 30670 16770
rect 34178 16718 34190 16770
rect 34242 16718 34254 16770
rect 50306 16718 50318 16770
rect 50370 16718 50382 16770
rect 25678 16706 25730 16718
rect 28366 16658 28418 16670
rect 10322 16606 10334 16658
rect 10386 16655 10398 16658
rect 10882 16655 10894 16658
rect 10386 16609 10894 16655
rect 10386 16606 10398 16609
rect 10882 16606 10894 16609
rect 10946 16606 10958 16658
rect 18946 16606 18958 16658
rect 19010 16655 19022 16658
rect 19506 16655 19518 16658
rect 19010 16609 19518 16655
rect 19010 16606 19022 16609
rect 19506 16606 19518 16609
rect 19570 16606 19582 16658
rect 28366 16594 28418 16606
rect 28478 16658 28530 16670
rect 30609 16655 30655 16718
rect 50766 16706 50818 16718
rect 52894 16770 52946 16782
rect 55906 16718 55918 16770
rect 55970 16718 55982 16770
rect 52894 16706 52946 16718
rect 40686 16658 40738 16670
rect 31266 16655 31278 16658
rect 30609 16609 31278 16655
rect 31266 16606 31278 16609
rect 31330 16606 31342 16658
rect 36082 16606 36094 16658
rect 36146 16606 36158 16658
rect 28478 16594 28530 16606
rect 40686 16594 40738 16606
rect 57486 16658 57538 16670
rect 57486 16594 57538 16606
rect 57598 16658 57650 16670
rect 57598 16594 57650 16606
rect 1344 16490 59024 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 59024 16490
rect 1344 16404 59024 16438
rect 11790 16322 11842 16334
rect 19070 16322 19122 16334
rect 13570 16270 13582 16322
rect 13634 16319 13646 16322
rect 14354 16319 14366 16322
rect 13634 16273 14366 16319
rect 13634 16270 13646 16273
rect 14354 16270 14366 16273
rect 14418 16270 14430 16322
rect 11790 16258 11842 16270
rect 19070 16258 19122 16270
rect 27582 16322 27634 16334
rect 29710 16322 29762 16334
rect 27794 16270 27806 16322
rect 27858 16319 27870 16322
rect 28354 16319 28366 16322
rect 27858 16273 28366 16319
rect 27858 16270 27870 16273
rect 28354 16270 28366 16273
rect 28418 16270 28430 16322
rect 27582 16258 27634 16270
rect 29710 16258 29762 16270
rect 30606 16322 30658 16334
rect 30606 16258 30658 16270
rect 31278 16322 31330 16334
rect 31278 16258 31330 16270
rect 42814 16322 42866 16334
rect 42814 16258 42866 16270
rect 45726 16322 45778 16334
rect 45726 16258 45778 16270
rect 6414 16210 6466 16222
rect 6414 16146 6466 16158
rect 7646 16210 7698 16222
rect 7646 16146 7698 16158
rect 12574 16210 12626 16222
rect 12574 16146 12626 16158
rect 13022 16210 13074 16222
rect 13022 16146 13074 16158
rect 14590 16210 14642 16222
rect 14590 16146 14642 16158
rect 19518 16210 19570 16222
rect 19518 16146 19570 16158
rect 19854 16210 19906 16222
rect 19854 16146 19906 16158
rect 20414 16210 20466 16222
rect 20414 16146 20466 16158
rect 20862 16210 20914 16222
rect 20862 16146 20914 16158
rect 21646 16210 21698 16222
rect 21646 16146 21698 16158
rect 22318 16210 22370 16222
rect 22318 16146 22370 16158
rect 23214 16210 23266 16222
rect 23214 16146 23266 16158
rect 23662 16210 23714 16222
rect 23662 16146 23714 16158
rect 24894 16210 24946 16222
rect 27470 16210 27522 16222
rect 26226 16158 26238 16210
rect 26290 16158 26302 16210
rect 24894 16146 24946 16158
rect 27470 16146 27522 16158
rect 28254 16210 28306 16222
rect 28254 16146 28306 16158
rect 29598 16210 29650 16222
rect 29598 16146 29650 16158
rect 31838 16210 31890 16222
rect 31838 16146 31890 16158
rect 32286 16210 32338 16222
rect 32286 16146 32338 16158
rect 32734 16210 32786 16222
rect 32734 16146 32786 16158
rect 33182 16210 33234 16222
rect 33182 16146 33234 16158
rect 34750 16210 34802 16222
rect 34750 16146 34802 16158
rect 37438 16210 37490 16222
rect 37438 16146 37490 16158
rect 37886 16210 37938 16222
rect 37886 16146 37938 16158
rect 38446 16210 38498 16222
rect 38446 16146 38498 16158
rect 41246 16210 41298 16222
rect 41246 16146 41298 16158
rect 41694 16210 41746 16222
rect 41694 16146 41746 16158
rect 42142 16210 42194 16222
rect 46622 16210 46674 16222
rect 55918 16210 55970 16222
rect 46050 16158 46062 16210
rect 46114 16158 46126 16210
rect 53666 16158 53678 16210
rect 53730 16158 53742 16210
rect 42142 16146 42194 16158
rect 46622 16146 46674 16158
rect 55918 16146 55970 16158
rect 8094 16098 8146 16110
rect 15374 16098 15426 16110
rect 22430 16098 22482 16110
rect 31166 16098 31218 16110
rect 8754 16046 8766 16098
rect 8818 16046 8830 16098
rect 16034 16046 16046 16098
rect 16098 16046 16110 16098
rect 26002 16046 26014 16098
rect 26066 16046 26078 16098
rect 8094 16034 8146 16046
rect 15374 16034 15426 16046
rect 22430 16034 22482 16046
rect 31166 16034 31218 16046
rect 34078 16098 34130 16110
rect 34078 16034 34130 16046
rect 35982 16098 36034 16110
rect 35982 16034 36034 16046
rect 39006 16098 39058 16110
rect 40686 16098 40738 16110
rect 40226 16046 40238 16098
rect 40290 16046 40302 16098
rect 39006 16034 39058 16046
rect 40686 16034 40738 16046
rect 43374 16098 43426 16110
rect 43374 16034 43426 16046
rect 43710 16098 43762 16110
rect 43710 16034 43762 16046
rect 52782 16098 52834 16110
rect 55010 16046 55022 16098
rect 55074 16046 55086 16098
rect 56130 16046 56142 16098
rect 56194 16046 56206 16098
rect 58482 16046 58494 16098
rect 58546 16046 58558 16098
rect 52782 16034 52834 16046
rect 18286 15986 18338 15998
rect 18286 15922 18338 15934
rect 22206 15986 22258 15998
rect 22206 15922 22258 15934
rect 22766 15986 22818 15998
rect 22766 15922 22818 15934
rect 25342 15986 25394 15998
rect 25342 15922 25394 15934
rect 27358 15986 27410 15998
rect 27358 15922 27410 15934
rect 30382 15986 30434 15998
rect 30382 15922 30434 15934
rect 31278 15986 31330 15998
rect 31278 15922 31330 15934
rect 34190 15986 34242 15998
rect 34190 15922 34242 15934
rect 35422 15986 35474 15998
rect 35422 15922 35474 15934
rect 35646 15986 35698 15998
rect 35646 15922 35698 15934
rect 36430 15986 36482 15998
rect 36430 15922 36482 15934
rect 39118 15986 39170 15998
rect 39118 15922 39170 15934
rect 39790 15986 39842 15998
rect 39790 15922 39842 15934
rect 42702 15986 42754 15998
rect 42702 15922 42754 15934
rect 42814 15986 42866 15998
rect 42814 15922 42866 15934
rect 44046 15986 44098 15998
rect 44046 15922 44098 15934
rect 44606 15986 44658 15998
rect 44606 15922 44658 15934
rect 45950 15986 46002 15998
rect 45950 15922 46002 15934
rect 52446 15986 52498 15998
rect 52446 15922 52498 15934
rect 53454 15986 53506 15998
rect 55234 15934 55246 15986
rect 55298 15934 55310 15986
rect 57810 15934 57822 15986
rect 57874 15934 57886 15986
rect 53454 15922 53506 15934
rect 5854 15874 5906 15886
rect 5854 15810 5906 15822
rect 6750 15874 6802 15886
rect 6750 15810 6802 15822
rect 7198 15874 7250 15886
rect 13582 15874 13634 15886
rect 11106 15822 11118 15874
rect 11170 15822 11182 15874
rect 7198 15810 7250 15822
rect 13582 15810 13634 15822
rect 14030 15874 14082 15886
rect 14030 15810 14082 15822
rect 15038 15874 15090 15886
rect 15038 15810 15090 15822
rect 24446 15874 24498 15886
rect 24446 15810 24498 15822
rect 28590 15874 28642 15886
rect 28590 15810 28642 15822
rect 30494 15874 30546 15886
rect 30494 15810 30546 15822
rect 34414 15874 34466 15886
rect 34414 15810 34466 15822
rect 35870 15874 35922 15886
rect 35870 15810 35922 15822
rect 39342 15874 39394 15886
rect 39342 15810 39394 15822
rect 43710 15874 43762 15886
rect 43710 15810 43762 15822
rect 46734 15874 46786 15886
rect 46734 15810 46786 15822
rect 49198 15874 49250 15886
rect 49198 15810 49250 15822
rect 52558 15874 52610 15886
rect 52558 15810 52610 15822
rect 53678 15874 53730 15886
rect 53678 15810 53730 15822
rect 1344 15706 59024 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 59024 15706
rect 1344 15620 59024 15654
rect 10558 15538 10610 15550
rect 10558 15474 10610 15486
rect 11006 15538 11058 15550
rect 11006 15474 11058 15486
rect 18062 15538 18114 15550
rect 18062 15474 18114 15486
rect 19742 15538 19794 15550
rect 19742 15474 19794 15486
rect 24558 15538 24610 15550
rect 24558 15474 24610 15486
rect 26238 15538 26290 15550
rect 26238 15474 26290 15486
rect 26574 15538 26626 15550
rect 26574 15474 26626 15486
rect 27022 15538 27074 15550
rect 27022 15474 27074 15486
rect 28030 15538 28082 15550
rect 28030 15474 28082 15486
rect 28478 15538 28530 15550
rect 28478 15474 28530 15486
rect 28926 15538 28978 15550
rect 28926 15474 28978 15486
rect 29374 15538 29426 15550
rect 29374 15474 29426 15486
rect 30718 15538 30770 15550
rect 30718 15474 30770 15486
rect 31390 15538 31442 15550
rect 31390 15474 31442 15486
rect 32286 15538 32338 15550
rect 32286 15474 32338 15486
rect 33630 15538 33682 15550
rect 33630 15474 33682 15486
rect 34526 15538 34578 15550
rect 34526 15474 34578 15486
rect 35198 15538 35250 15550
rect 35198 15474 35250 15486
rect 38894 15538 38946 15550
rect 43934 15538 43986 15550
rect 42914 15486 42926 15538
rect 42978 15486 42990 15538
rect 38894 15474 38946 15486
rect 43934 15474 43986 15486
rect 45838 15538 45890 15550
rect 45838 15474 45890 15486
rect 48638 15538 48690 15550
rect 48638 15474 48690 15486
rect 49758 15538 49810 15550
rect 55682 15486 55694 15538
rect 55746 15486 55758 15538
rect 49758 15474 49810 15486
rect 17614 15426 17666 15438
rect 5394 15374 5406 15426
rect 5458 15374 5470 15426
rect 16594 15374 16606 15426
rect 16658 15374 16670 15426
rect 17614 15362 17666 15374
rect 22206 15426 22258 15438
rect 22206 15362 22258 15374
rect 23886 15426 23938 15438
rect 23886 15362 23938 15374
rect 24894 15426 24946 15438
rect 24894 15362 24946 15374
rect 31614 15426 31666 15438
rect 31614 15362 31666 15374
rect 37438 15426 37490 15438
rect 37438 15362 37490 15374
rect 37998 15426 38050 15438
rect 37998 15362 38050 15374
rect 39230 15426 39282 15438
rect 39230 15362 39282 15374
rect 40798 15426 40850 15438
rect 40798 15362 40850 15374
rect 41806 15426 41858 15438
rect 41806 15362 41858 15374
rect 42366 15426 42418 15438
rect 42366 15362 42418 15374
rect 43710 15426 43762 15438
rect 43710 15362 43762 15374
rect 45054 15426 45106 15438
rect 45054 15362 45106 15374
rect 45614 15426 45666 15438
rect 45614 15362 45666 15374
rect 45950 15426 46002 15438
rect 45950 15362 46002 15374
rect 46174 15426 46226 15438
rect 46174 15362 46226 15374
rect 47182 15426 47234 15438
rect 47182 15362 47234 15374
rect 49982 15426 50034 15438
rect 57486 15426 57538 15438
rect 52546 15374 52558 15426
rect 52610 15374 52622 15426
rect 56354 15374 56366 15426
rect 56418 15374 56430 15426
rect 49982 15362 50034 15374
rect 57486 15362 57538 15374
rect 18510 15314 18562 15326
rect 23774 15314 23826 15326
rect 8306 15262 8318 15314
rect 8370 15262 8382 15314
rect 11778 15262 11790 15314
rect 11842 15262 11854 15314
rect 21186 15262 21198 15314
rect 21250 15262 21262 15314
rect 21410 15262 21422 15314
rect 21474 15262 21486 15314
rect 22866 15262 22878 15314
rect 22930 15262 22942 15314
rect 18510 15250 18562 15262
rect 23774 15250 23826 15262
rect 25678 15314 25730 15326
rect 25678 15250 25730 15262
rect 27470 15314 27522 15326
rect 30606 15314 30658 15326
rect 30482 15262 30494 15314
rect 30546 15262 30558 15314
rect 27470 15250 27522 15262
rect 30606 15250 30658 15262
rect 30830 15314 30882 15326
rect 30830 15250 30882 15262
rect 31726 15314 31778 15326
rect 31726 15250 31778 15262
rect 33966 15314 34018 15326
rect 33966 15250 34018 15262
rect 35870 15314 35922 15326
rect 35870 15250 35922 15262
rect 35982 15314 36034 15326
rect 35982 15250 36034 15262
rect 36206 15314 36258 15326
rect 36206 15250 36258 15262
rect 36766 15314 36818 15326
rect 36766 15250 36818 15262
rect 37214 15314 37266 15326
rect 39902 15314 39954 15326
rect 42590 15314 42642 15326
rect 38322 15262 38334 15314
rect 38386 15262 38398 15314
rect 40338 15262 40350 15314
rect 40402 15262 40414 15314
rect 37214 15250 37266 15262
rect 39902 15250 39954 15262
rect 42590 15250 42642 15262
rect 43486 15314 43538 15326
rect 43486 15250 43538 15262
rect 49534 15314 49586 15326
rect 49534 15250 49586 15262
rect 49646 15314 49698 15326
rect 54238 15314 54290 15326
rect 57598 15314 57650 15326
rect 52434 15262 52446 15314
rect 52498 15262 52510 15314
rect 52658 15262 52670 15314
rect 52722 15262 52734 15314
rect 53330 15262 53342 15314
rect 53394 15262 53406 15314
rect 54786 15262 54798 15314
rect 54850 15262 54862 15314
rect 55570 15262 55582 15314
rect 55634 15262 55646 15314
rect 56690 15262 56702 15314
rect 56754 15262 56766 15314
rect 57922 15262 57934 15314
rect 57986 15262 57998 15314
rect 49646 15250 49698 15262
rect 54238 15250 54290 15262
rect 57598 15250 57650 15262
rect 9662 15202 9714 15214
rect 9662 15138 9714 15150
rect 19294 15202 19346 15214
rect 19294 15138 19346 15150
rect 21646 15202 21698 15214
rect 32622 15202 32674 15214
rect 22978 15150 22990 15202
rect 23042 15150 23054 15202
rect 21646 15138 21698 15150
rect 32622 15138 32674 15150
rect 37326 15202 37378 15214
rect 37326 15138 37378 15150
rect 43598 15202 43650 15214
rect 48414 15202 48466 15214
rect 47282 15150 47294 15202
rect 47346 15150 47358 15202
rect 43598 15138 43650 15150
rect 48414 15138 48466 15150
rect 30158 15090 30210 15102
rect 30158 15026 30210 15038
rect 36318 15090 36370 15102
rect 36318 15026 36370 15038
rect 38334 15090 38386 15102
rect 38334 15026 38386 15038
rect 46958 15090 47010 15102
rect 46958 15026 47010 15038
rect 48750 15090 48802 15102
rect 48750 15026 48802 15038
rect 54462 15090 54514 15102
rect 54462 15026 54514 15038
rect 1344 14922 59024 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 59024 14922
rect 1344 14836 59024 14870
rect 13022 14754 13074 14766
rect 7186 14702 7198 14754
rect 7250 14751 7262 14754
rect 8194 14751 8206 14754
rect 7250 14705 8206 14751
rect 7250 14702 7262 14705
rect 8194 14702 8206 14705
rect 8258 14702 8270 14754
rect 13022 14690 13074 14702
rect 19070 14754 19122 14766
rect 19070 14690 19122 14702
rect 27694 14754 27746 14766
rect 27694 14690 27746 14702
rect 30158 14754 30210 14766
rect 35086 14754 35138 14766
rect 30594 14702 30606 14754
rect 30658 14751 30670 14754
rect 31602 14751 31614 14754
rect 30658 14705 31614 14751
rect 30658 14702 30670 14705
rect 31602 14702 31614 14705
rect 31666 14702 31678 14754
rect 33842 14702 33854 14754
rect 33906 14702 33918 14754
rect 30158 14690 30210 14702
rect 35086 14690 35138 14702
rect 35422 14754 35474 14766
rect 51886 14754 51938 14766
rect 35634 14702 35646 14754
rect 35698 14751 35710 14754
rect 36418 14751 36430 14754
rect 35698 14705 36430 14751
rect 35698 14702 35710 14705
rect 36418 14702 36430 14705
rect 36482 14702 36494 14754
rect 43138 14702 43150 14754
rect 43202 14751 43214 14754
rect 43474 14751 43486 14754
rect 43202 14705 43486 14751
rect 43202 14702 43214 14705
rect 43474 14702 43486 14705
rect 43538 14702 43550 14754
rect 52210 14702 52222 14754
rect 52274 14702 52286 14754
rect 35422 14690 35474 14702
rect 51886 14690 51938 14702
rect 4958 14642 5010 14654
rect 4958 14578 5010 14590
rect 5630 14642 5682 14654
rect 5630 14578 5682 14590
rect 6414 14642 6466 14654
rect 6414 14578 6466 14590
rect 6862 14642 6914 14654
rect 6862 14578 6914 14590
rect 7310 14642 7362 14654
rect 7310 14578 7362 14590
rect 7758 14642 7810 14654
rect 7758 14578 7810 14590
rect 8766 14642 8818 14654
rect 8766 14578 8818 14590
rect 13694 14642 13746 14654
rect 13694 14578 13746 14590
rect 14030 14642 14082 14654
rect 23886 14642 23938 14654
rect 22754 14590 22766 14642
rect 22818 14590 22830 14642
rect 14030 14578 14082 14590
rect 23886 14578 23938 14590
rect 26574 14642 26626 14654
rect 26574 14578 26626 14590
rect 31054 14642 31106 14654
rect 31054 14578 31106 14590
rect 31390 14642 31442 14654
rect 31390 14578 31442 14590
rect 35982 14642 36034 14654
rect 35982 14578 36034 14590
rect 36766 14642 36818 14654
rect 36766 14578 36818 14590
rect 43150 14642 43202 14654
rect 44718 14642 44770 14654
rect 48862 14642 48914 14654
rect 50318 14642 50370 14654
rect 44258 14590 44270 14642
rect 44322 14590 44334 14642
rect 46498 14590 46510 14642
rect 46562 14590 46574 14642
rect 49634 14590 49646 14642
rect 49698 14590 49710 14642
rect 43150 14578 43202 14590
rect 44718 14578 44770 14590
rect 48862 14578 48914 14590
rect 50318 14578 50370 14590
rect 54686 14642 54738 14654
rect 54686 14578 54738 14590
rect 55582 14642 55634 14654
rect 57262 14642 57314 14654
rect 56466 14590 56478 14642
rect 56530 14590 56542 14642
rect 55582 14578 55634 14590
rect 57262 14578 57314 14590
rect 9550 14530 9602 14542
rect 15374 14530 15426 14542
rect 25118 14530 25170 14542
rect 9986 14478 9998 14530
rect 10050 14478 10062 14530
rect 16034 14478 16046 14530
rect 16098 14478 16110 14530
rect 21858 14478 21870 14530
rect 21922 14478 21934 14530
rect 9550 14466 9602 14478
rect 15374 14466 15426 14478
rect 25118 14466 25170 14478
rect 27134 14530 27186 14542
rect 32734 14530 32786 14542
rect 30482 14478 30494 14530
rect 30546 14478 30558 14530
rect 32498 14478 32510 14530
rect 32562 14478 32574 14530
rect 27134 14466 27186 14478
rect 32734 14466 32786 14478
rect 34078 14530 34130 14542
rect 34078 14466 34130 14478
rect 34526 14530 34578 14542
rect 51662 14530 51714 14542
rect 38322 14478 38334 14530
rect 38386 14478 38398 14530
rect 44034 14478 44046 14530
rect 44098 14478 44110 14530
rect 46834 14478 46846 14530
rect 46898 14478 46910 14530
rect 49970 14478 49982 14530
rect 50034 14478 50046 14530
rect 54226 14478 54238 14530
rect 54290 14478 54302 14530
rect 54450 14478 54462 14530
rect 54514 14478 54526 14530
rect 56242 14478 56254 14530
rect 56306 14478 56318 14530
rect 34526 14466 34578 14478
rect 51662 14466 51714 14478
rect 18286 14418 18338 14430
rect 18286 14354 18338 14366
rect 22766 14418 22818 14430
rect 22766 14354 22818 14366
rect 22990 14418 23042 14430
rect 22990 14354 23042 14366
rect 27582 14418 27634 14430
rect 27582 14354 27634 14366
rect 29710 14418 29762 14430
rect 35310 14418 35362 14430
rect 29922 14366 29934 14418
rect 29986 14366 29998 14418
rect 29710 14354 29762 14366
rect 35310 14354 35362 14366
rect 36318 14418 36370 14430
rect 47406 14418 47458 14430
rect 38098 14366 38110 14418
rect 38162 14366 38174 14418
rect 39554 14366 39566 14418
rect 39618 14366 39630 14418
rect 36318 14354 36370 14366
rect 47406 14354 47458 14366
rect 8206 14306 8258 14318
rect 14478 14306 14530 14318
rect 12450 14254 12462 14306
rect 12514 14254 12526 14306
rect 8206 14242 8258 14254
rect 14478 14242 14530 14254
rect 14926 14306 14978 14318
rect 14926 14242 14978 14254
rect 19406 14306 19458 14318
rect 19406 14242 19458 14254
rect 21646 14306 21698 14318
rect 21646 14242 21698 14254
rect 24222 14306 24274 14318
rect 24222 14242 24274 14254
rect 24782 14306 24834 14318
rect 24782 14242 24834 14254
rect 25902 14306 25954 14318
rect 25902 14242 25954 14254
rect 26462 14306 26514 14318
rect 26462 14242 26514 14254
rect 26686 14306 26738 14318
rect 26686 14242 26738 14254
rect 27694 14306 27746 14318
rect 27694 14242 27746 14254
rect 28366 14306 28418 14318
rect 28366 14242 28418 14254
rect 28814 14306 28866 14318
rect 31838 14306 31890 14318
rect 30034 14254 30046 14306
rect 30098 14254 30110 14306
rect 28814 14242 28866 14254
rect 31838 14242 31890 14254
rect 32846 14306 32898 14318
rect 32846 14242 32898 14254
rect 32958 14306 33010 14318
rect 32958 14242 33010 14254
rect 33070 14306 33122 14318
rect 42030 14306 42082 14318
rect 39666 14254 39678 14306
rect 39730 14254 39742 14306
rect 33070 14242 33122 14254
rect 42030 14242 42082 14254
rect 47854 14306 47906 14318
rect 47854 14242 47906 14254
rect 58494 14306 58546 14318
rect 58494 14242 58546 14254
rect 1344 14138 59024 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 59024 14138
rect 1344 14052 59024 14086
rect 8878 13970 8930 13982
rect 8082 13918 8094 13970
rect 8146 13918 8158 13970
rect 8878 13906 8930 13918
rect 9662 13970 9714 13982
rect 9662 13906 9714 13918
rect 10110 13970 10162 13982
rect 22542 13970 22594 13982
rect 13682 13918 13694 13970
rect 13746 13918 13758 13970
rect 10110 13906 10162 13918
rect 22542 13906 22594 13918
rect 23438 13970 23490 13982
rect 23438 13906 23490 13918
rect 28590 13970 28642 13982
rect 28590 13906 28642 13918
rect 29150 13970 29202 13982
rect 29150 13906 29202 13918
rect 29598 13970 29650 13982
rect 29598 13906 29650 13918
rect 31502 13970 31554 13982
rect 31502 13906 31554 13918
rect 39790 13970 39842 13982
rect 39790 13906 39842 13918
rect 44158 13970 44210 13982
rect 44158 13906 44210 13918
rect 46062 13970 46114 13982
rect 46062 13906 46114 13918
rect 48190 13970 48242 13982
rect 48190 13906 48242 13918
rect 55358 13970 55410 13982
rect 55358 13906 55410 13918
rect 55806 13970 55858 13982
rect 55806 13906 55858 13918
rect 30830 13858 30882 13870
rect 35422 13858 35474 13870
rect 34290 13806 34302 13858
rect 34354 13806 34366 13858
rect 34626 13806 34638 13858
rect 34690 13806 34702 13858
rect 30830 13794 30882 13806
rect 35422 13794 35474 13806
rect 37774 13858 37826 13870
rect 37774 13794 37826 13806
rect 37998 13858 38050 13870
rect 37998 13794 38050 13806
rect 38334 13858 38386 13870
rect 46622 13858 46674 13870
rect 42690 13806 42702 13858
rect 42754 13806 42766 13858
rect 43026 13806 43038 13858
rect 43090 13806 43102 13858
rect 38334 13794 38386 13806
rect 46622 13794 46674 13806
rect 46846 13858 46898 13870
rect 46846 13794 46898 13806
rect 47630 13858 47682 13870
rect 47630 13794 47682 13806
rect 47742 13858 47794 13870
rect 52658 13806 52670 13858
rect 52722 13806 52734 13858
rect 53778 13806 53790 13858
rect 53842 13806 53854 13858
rect 47742 13794 47794 13806
rect 5406 13746 5458 13758
rect 10558 13746 10610 13758
rect 16270 13746 16322 13758
rect 4274 13694 4286 13746
rect 4338 13694 4350 13746
rect 5730 13694 5742 13746
rect 5794 13694 5806 13746
rect 11218 13694 11230 13746
rect 11282 13694 11294 13746
rect 5406 13682 5458 13694
rect 10558 13682 10610 13694
rect 16270 13682 16322 13694
rect 22430 13746 22482 13758
rect 22430 13682 22482 13694
rect 22654 13746 22706 13758
rect 22654 13682 22706 13694
rect 23102 13746 23154 13758
rect 23102 13682 23154 13694
rect 24334 13746 24386 13758
rect 32398 13746 32450 13758
rect 26114 13694 26126 13746
rect 26178 13694 26190 13746
rect 27682 13694 27694 13746
rect 27746 13694 27758 13746
rect 32162 13694 32174 13746
rect 32226 13694 32238 13746
rect 24334 13682 24386 13694
rect 32398 13682 32450 13694
rect 32622 13746 32674 13758
rect 33742 13746 33794 13758
rect 32834 13694 32846 13746
rect 32898 13694 32910 13746
rect 32622 13682 32674 13694
rect 33742 13682 33794 13694
rect 43262 13746 43314 13758
rect 43262 13682 43314 13694
rect 47406 13746 47458 13758
rect 47406 13682 47458 13694
rect 14926 13634 14978 13646
rect 3938 13582 3950 13634
rect 4002 13582 4014 13634
rect 14926 13570 14978 13582
rect 15374 13634 15426 13646
rect 15374 13570 15426 13582
rect 15822 13634 15874 13646
rect 15822 13570 15874 13582
rect 19182 13634 19234 13646
rect 19182 13570 19234 13582
rect 19742 13634 19794 13646
rect 19742 13570 19794 13582
rect 24894 13634 24946 13646
rect 30046 13634 30098 13646
rect 26450 13582 26462 13634
rect 26514 13582 26526 13634
rect 24894 13570 24946 13582
rect 30046 13570 30098 13582
rect 32510 13634 32562 13646
rect 32510 13570 32562 13582
rect 34078 13634 34130 13646
rect 34078 13570 34130 13582
rect 38222 13634 38274 13646
rect 38222 13570 38274 13582
rect 41470 13634 41522 13646
rect 41470 13570 41522 13582
rect 45614 13634 45666 13646
rect 51986 13582 51998 13634
rect 52050 13582 52062 13634
rect 45614 13570 45666 13582
rect 14254 13522 14306 13534
rect 30942 13522 30994 13534
rect 4274 13470 4286 13522
rect 4338 13470 4350 13522
rect 27570 13470 27582 13522
rect 27634 13470 27646 13522
rect 29698 13470 29710 13522
rect 29762 13519 29774 13522
rect 29922 13519 29934 13522
rect 29762 13473 29934 13519
rect 29762 13470 29774 13473
rect 29922 13470 29934 13473
rect 29986 13470 29998 13522
rect 14254 13458 14306 13470
rect 30942 13458 30994 13470
rect 43598 13522 43650 13534
rect 43598 13458 43650 13470
rect 46958 13522 47010 13534
rect 46958 13458 47010 13470
rect 54798 13522 54850 13534
rect 54798 13458 54850 13470
rect 1344 13354 59024 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 59024 13354
rect 1344 13268 59024 13302
rect 10222 13186 10274 13198
rect 10222 13122 10274 13134
rect 19070 13186 19122 13198
rect 19070 13122 19122 13134
rect 26574 13186 26626 13198
rect 26574 13122 26626 13134
rect 30046 13186 30098 13198
rect 30046 13122 30098 13134
rect 52334 13186 52386 13198
rect 52334 13122 52386 13134
rect 52670 13186 52722 13198
rect 52670 13122 52722 13134
rect 10894 13074 10946 13086
rect 10894 13010 10946 13022
rect 11342 13074 11394 13086
rect 11342 13010 11394 13022
rect 12350 13074 12402 13086
rect 12350 13010 12402 13022
rect 13582 13074 13634 13086
rect 13582 13010 13634 13022
rect 14590 13074 14642 13086
rect 23662 13074 23714 13086
rect 19618 13022 19630 13074
rect 19682 13022 19694 13074
rect 14590 13010 14642 13022
rect 23662 13010 23714 13022
rect 25454 13074 25506 13086
rect 25454 13010 25506 13022
rect 26462 13074 26514 13086
rect 26462 13010 26514 13022
rect 28030 13074 28082 13086
rect 28030 13010 28082 13022
rect 31166 13074 31218 13086
rect 31166 13010 31218 13022
rect 31726 13074 31778 13086
rect 31726 13010 31778 13022
rect 32174 13074 32226 13086
rect 32174 13010 32226 13022
rect 32734 13074 32786 13086
rect 34974 13074 35026 13086
rect 33730 13022 33742 13074
rect 33794 13022 33806 13074
rect 32734 13010 32786 13022
rect 34974 13010 35026 13022
rect 37662 13074 37714 13086
rect 37662 13010 37714 13022
rect 38894 13074 38946 13086
rect 38894 13010 38946 13022
rect 41918 13074 41970 13086
rect 41918 13010 41970 13022
rect 43822 13074 43874 13086
rect 43822 13010 43874 13022
rect 45726 13074 45778 13086
rect 51214 13074 51266 13086
rect 46610 13022 46622 13074
rect 46674 13022 46686 13074
rect 49298 13022 49310 13074
rect 49362 13022 49374 13074
rect 45726 13010 45778 13022
rect 51214 13010 51266 13022
rect 52110 13074 52162 13086
rect 52110 13010 52162 13022
rect 3838 12962 3890 12974
rect 3838 12898 3890 12910
rect 5630 12962 5682 12974
rect 10446 12962 10498 12974
rect 6178 12910 6190 12962
rect 6242 12910 6254 12962
rect 5630 12898 5682 12910
rect 10446 12898 10498 12910
rect 11902 12962 11954 12974
rect 11902 12898 11954 12910
rect 12910 12962 12962 12974
rect 12910 12898 12962 12910
rect 15374 12962 15426 12974
rect 27470 12962 27522 12974
rect 16034 12910 16046 12962
rect 16098 12910 16110 12962
rect 20514 12910 20526 12962
rect 20578 12910 20590 12962
rect 22306 12910 22318 12962
rect 22370 12910 22382 12962
rect 15374 12898 15426 12910
rect 27470 12898 27522 12910
rect 29710 12962 29762 12974
rect 29710 12898 29762 12910
rect 29822 12962 29874 12974
rect 29822 12898 29874 12910
rect 31390 12962 31442 12974
rect 40126 12962 40178 12974
rect 33506 12910 33518 12962
rect 33570 12910 33582 12962
rect 37762 12910 37774 12962
rect 37826 12910 37838 12962
rect 31390 12898 31442 12910
rect 40126 12898 40178 12910
rect 40798 12962 40850 12974
rect 40798 12898 40850 12910
rect 41246 12962 41298 12974
rect 50990 12962 51042 12974
rect 43138 12910 43150 12962
rect 43202 12910 43214 12962
rect 43586 12910 43598 12962
rect 43650 12910 43662 12962
rect 46386 12910 46398 12962
rect 46450 12910 46462 12962
rect 47730 12910 47742 12962
rect 47794 12910 47806 12962
rect 49746 12910 49758 12962
rect 49810 12910 49822 12962
rect 41246 12898 41298 12910
rect 50990 12898 51042 12910
rect 56478 12962 56530 12974
rect 56478 12898 56530 12910
rect 3502 12850 3554 12862
rect 3502 12786 3554 12798
rect 4286 12850 4338 12862
rect 4286 12786 4338 12798
rect 4734 12850 4786 12862
rect 18286 12850 18338 12862
rect 24782 12850 24834 12862
rect 9874 12798 9886 12850
rect 9938 12798 9950 12850
rect 23202 12798 23214 12850
rect 23266 12798 23278 12850
rect 4734 12786 4786 12798
rect 18286 12786 18338 12798
rect 24782 12786 24834 12798
rect 26350 12850 26402 12862
rect 26350 12786 26402 12798
rect 30158 12850 30210 12862
rect 30158 12786 30210 12798
rect 30718 12850 30770 12862
rect 30718 12786 30770 12798
rect 30942 12850 30994 12862
rect 30942 12786 30994 12798
rect 34414 12850 34466 12862
rect 34414 12786 34466 12798
rect 37550 12850 37602 12862
rect 37550 12786 37602 12798
rect 39566 12850 39618 12862
rect 39566 12786 39618 12798
rect 41358 12850 41410 12862
rect 41358 12786 41410 12798
rect 48526 12850 48578 12862
rect 48526 12786 48578 12798
rect 50206 12850 50258 12862
rect 50206 12786 50258 12798
rect 50766 12850 50818 12862
rect 50766 12786 50818 12798
rect 51326 12850 51378 12862
rect 51326 12786 51378 12798
rect 3614 12738 3666 12750
rect 3614 12674 3666 12686
rect 4510 12738 4562 12750
rect 4510 12674 4562 12686
rect 4846 12738 4898 12750
rect 9326 12738 9378 12750
rect 8754 12686 8766 12738
rect 8818 12686 8830 12738
rect 4846 12674 4898 12686
rect 9326 12674 9378 12686
rect 14142 12738 14194 12750
rect 24334 12738 24386 12750
rect 21746 12686 21758 12738
rect 21810 12686 21822 12738
rect 14142 12674 14194 12686
rect 24334 12674 24386 12686
rect 27134 12738 27186 12750
rect 27134 12674 27186 12686
rect 28366 12738 28418 12750
rect 28366 12674 28418 12686
rect 28814 12738 28866 12750
rect 28814 12674 28866 12686
rect 37998 12738 38050 12750
rect 37998 12674 38050 12686
rect 38446 12738 38498 12750
rect 38446 12674 38498 12686
rect 39454 12738 39506 12750
rect 39454 12674 39506 12686
rect 40238 12738 40290 12750
rect 40238 12674 40290 12686
rect 40350 12738 40402 12750
rect 40350 12674 40402 12686
rect 41582 12738 41634 12750
rect 41582 12674 41634 12686
rect 56254 12738 56306 12750
rect 56254 12674 56306 12686
rect 56366 12738 56418 12750
rect 56366 12674 56418 12686
rect 1344 12570 59024 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 59024 12570
rect 1344 12484 59024 12518
rect 9662 12402 9714 12414
rect 6178 12350 6190 12402
rect 6242 12350 6254 12402
rect 9662 12338 9714 12350
rect 10110 12402 10162 12414
rect 10110 12338 10162 12350
rect 10670 12402 10722 12414
rect 10670 12338 10722 12350
rect 20190 12402 20242 12414
rect 20190 12338 20242 12350
rect 22654 12402 22706 12414
rect 22654 12338 22706 12350
rect 22766 12402 22818 12414
rect 22766 12338 22818 12350
rect 23326 12402 23378 12414
rect 23326 12338 23378 12350
rect 23550 12402 23602 12414
rect 23550 12338 23602 12350
rect 26014 12402 26066 12414
rect 26014 12338 26066 12350
rect 27246 12402 27298 12414
rect 27246 12338 27298 12350
rect 28030 12402 28082 12414
rect 28030 12338 28082 12350
rect 28702 12402 28754 12414
rect 28702 12338 28754 12350
rect 31950 12402 32002 12414
rect 31950 12338 32002 12350
rect 32398 12402 32450 12414
rect 32398 12338 32450 12350
rect 32958 12402 33010 12414
rect 32958 12338 33010 12350
rect 33518 12402 33570 12414
rect 33518 12338 33570 12350
rect 33966 12402 34018 12414
rect 33966 12338 34018 12350
rect 35422 12402 35474 12414
rect 35422 12338 35474 12350
rect 40462 12402 40514 12414
rect 40462 12338 40514 12350
rect 42030 12402 42082 12414
rect 42030 12338 42082 12350
rect 43038 12402 43090 12414
rect 43038 12338 43090 12350
rect 43486 12402 43538 12414
rect 43486 12338 43538 12350
rect 43934 12402 43986 12414
rect 43934 12338 43986 12350
rect 45950 12402 46002 12414
rect 45950 12338 46002 12350
rect 47630 12402 47682 12414
rect 47630 12338 47682 12350
rect 49646 12402 49698 12414
rect 49646 12338 49698 12350
rect 49758 12402 49810 12414
rect 56578 12350 56590 12402
rect 56642 12350 56654 12402
rect 49758 12338 49810 12350
rect 21422 12290 21474 12302
rect 15138 12238 15150 12290
rect 15202 12238 15214 12290
rect 21422 12226 21474 12238
rect 21758 12290 21810 12302
rect 21758 12226 21810 12238
rect 22878 12290 22930 12302
rect 22878 12226 22930 12238
rect 23662 12290 23714 12302
rect 23662 12226 23714 12238
rect 24334 12290 24386 12302
rect 24334 12226 24386 12238
rect 30494 12290 30546 12302
rect 30494 12226 30546 12238
rect 31054 12290 31106 12302
rect 31054 12226 31106 12238
rect 34974 12290 35026 12302
rect 34974 12226 35026 12238
rect 36878 12290 36930 12302
rect 36878 12226 36930 12238
rect 36990 12290 37042 12302
rect 36990 12226 37042 12238
rect 38894 12290 38946 12302
rect 38894 12226 38946 12238
rect 39454 12290 39506 12302
rect 39454 12226 39506 12238
rect 41806 12290 41858 12302
rect 41806 12226 41858 12238
rect 42590 12290 42642 12302
rect 42590 12226 42642 12238
rect 47182 12290 47234 12302
rect 47182 12226 47234 12238
rect 47406 12290 47458 12302
rect 47406 12226 47458 12238
rect 47742 12290 47794 12302
rect 47742 12226 47794 12238
rect 49534 12290 49586 12302
rect 49534 12226 49586 12238
rect 53902 12290 53954 12302
rect 57598 12290 57650 12302
rect 56018 12238 56030 12290
rect 56082 12238 56094 12290
rect 53902 12226 53954 12238
rect 57598 12226 57650 12238
rect 5406 12178 5458 12190
rect 9102 12178 9154 12190
rect 4162 12126 4174 12178
rect 4226 12126 4238 12178
rect 8418 12126 8430 12178
rect 8482 12126 8494 12178
rect 5406 12114 5458 12126
rect 9102 12114 9154 12126
rect 11230 12178 11282 12190
rect 28814 12178 28866 12190
rect 11666 12126 11678 12178
rect 11730 12126 11742 12178
rect 18722 12126 18734 12178
rect 18786 12126 18798 12178
rect 11230 12114 11282 12126
rect 28814 12114 28866 12126
rect 29598 12178 29650 12190
rect 36654 12178 36706 12190
rect 39230 12178 39282 12190
rect 30034 12126 30046 12178
rect 30098 12126 30110 12178
rect 31266 12126 31278 12178
rect 31330 12126 31342 12178
rect 34626 12126 34638 12178
rect 34690 12126 34702 12178
rect 37314 12126 37326 12178
rect 37378 12126 37390 12178
rect 29598 12114 29650 12126
rect 36654 12114 36706 12126
rect 39230 12114 39282 12126
rect 40238 12178 40290 12190
rect 40238 12114 40290 12126
rect 40686 12178 40738 12190
rect 40686 12114 40738 12126
rect 41582 12178 41634 12190
rect 57374 12178 57426 12190
rect 55570 12126 55582 12178
rect 55634 12126 55646 12178
rect 56466 12126 56478 12178
rect 56530 12126 56542 12178
rect 41582 12114 41634 12126
rect 57374 12114 57426 12126
rect 57710 12178 57762 12190
rect 57710 12114 57762 12126
rect 4622 12066 4674 12078
rect 24446 12066 24498 12078
rect 4274 12014 4286 12066
rect 4338 12014 4350 12066
rect 19170 12014 19182 12066
rect 19234 12014 19246 12066
rect 4622 12002 4674 12014
rect 24446 12002 24498 12014
rect 26462 12066 26514 12078
rect 26462 12002 26514 12014
rect 27582 12066 27634 12078
rect 37886 12066 37938 12078
rect 37426 12014 37438 12066
rect 37490 12014 37502 12066
rect 27582 12002 27634 12014
rect 37886 12002 37938 12014
rect 38334 12066 38386 12078
rect 38334 12002 38386 12014
rect 39006 12066 39058 12078
rect 39006 12002 39058 12014
rect 40574 12066 40626 12078
rect 40574 12002 40626 12014
rect 41694 12066 41746 12078
rect 41694 12002 41746 12014
rect 45166 12066 45218 12078
rect 45166 12002 45218 12014
rect 28926 11954 28978 11966
rect 34638 11954 34690 11966
rect 32274 11902 32286 11954
rect 32338 11951 32350 11954
rect 32834 11951 32846 11954
rect 32338 11905 32846 11951
rect 32338 11902 32350 11905
rect 32834 11902 32846 11905
rect 32898 11902 32910 11954
rect 33842 11902 33854 11954
rect 33906 11951 33918 11954
rect 34402 11951 34414 11954
rect 33906 11905 34414 11951
rect 33906 11902 33918 11905
rect 34402 11902 34414 11905
rect 34466 11902 34478 11954
rect 28926 11890 28978 11902
rect 34638 11890 34690 11902
rect 40014 11954 40066 11966
rect 40014 11890 40066 11902
rect 53678 11954 53730 11966
rect 53678 11890 53730 11902
rect 54014 11954 54066 11966
rect 54014 11890 54066 11902
rect 1344 11786 59024 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 59024 11786
rect 1344 11700 59024 11734
rect 24670 11618 24722 11630
rect 33518 11618 33570 11630
rect 10882 11566 10894 11618
rect 10946 11615 10958 11618
rect 11666 11615 11678 11618
rect 10946 11569 11678 11615
rect 10946 11566 10958 11569
rect 11666 11566 11678 11569
rect 11730 11566 11742 11618
rect 26562 11566 26574 11618
rect 26626 11566 26638 11618
rect 24670 11554 24722 11566
rect 33518 11554 33570 11566
rect 35310 11618 35362 11630
rect 35310 11554 35362 11566
rect 41246 11618 41298 11630
rect 42814 11618 42866 11630
rect 41458 11566 41470 11618
rect 41522 11615 41534 11618
rect 41794 11615 41806 11618
rect 41522 11569 41806 11615
rect 41522 11566 41534 11569
rect 41794 11566 41806 11569
rect 41858 11566 41870 11618
rect 41246 11554 41298 11566
rect 42814 11554 42866 11566
rect 5070 11506 5122 11518
rect 5070 11442 5122 11454
rect 8094 11506 8146 11518
rect 11118 11506 11170 11518
rect 10546 11454 10558 11506
rect 10610 11454 10622 11506
rect 8094 11442 8146 11454
rect 11118 11442 11170 11454
rect 11678 11506 11730 11518
rect 11678 11442 11730 11454
rect 19070 11506 19122 11518
rect 19070 11442 19122 11454
rect 19630 11506 19682 11518
rect 19630 11442 19682 11454
rect 21646 11506 21698 11518
rect 21646 11442 21698 11454
rect 22318 11506 22370 11518
rect 22318 11442 22370 11454
rect 23214 11506 23266 11518
rect 23214 11442 23266 11454
rect 28366 11506 28418 11518
rect 28366 11442 28418 11454
rect 30606 11506 30658 11518
rect 30606 11442 30658 11454
rect 32958 11506 33010 11518
rect 41134 11506 41186 11518
rect 38994 11454 39006 11506
rect 39058 11454 39070 11506
rect 32958 11442 33010 11454
rect 41134 11442 41186 11454
rect 41806 11506 41858 11518
rect 41806 11442 41858 11454
rect 42142 11506 42194 11518
rect 42142 11442 42194 11454
rect 45502 11506 45554 11518
rect 56478 11506 56530 11518
rect 51314 11454 51326 11506
rect 51378 11454 51390 11506
rect 45502 11442 45554 11454
rect 56478 11442 56530 11454
rect 5742 11394 5794 11406
rect 5742 11330 5794 11342
rect 6638 11394 6690 11406
rect 22094 11394 22146 11406
rect 8978 11342 8990 11394
rect 9042 11342 9054 11394
rect 10322 11342 10334 11394
rect 10386 11342 10398 11394
rect 15474 11342 15486 11394
rect 15538 11342 15550 11394
rect 16034 11342 16046 11394
rect 16098 11342 16110 11394
rect 6638 11330 6690 11342
rect 22094 11330 22146 11342
rect 22430 11394 22482 11406
rect 22430 11330 22482 11342
rect 25342 11394 25394 11406
rect 25342 11330 25394 11342
rect 27470 11394 27522 11406
rect 30494 11394 30546 11406
rect 34190 11394 34242 11406
rect 44606 11394 44658 11406
rect 30146 11342 30158 11394
rect 30210 11342 30222 11394
rect 33842 11342 33854 11394
rect 33906 11342 33918 11394
rect 38770 11342 38782 11394
rect 38834 11342 38846 11394
rect 40450 11342 40462 11394
rect 40514 11342 40526 11394
rect 44034 11342 44046 11394
rect 44098 11342 44110 11394
rect 27470 11330 27522 11342
rect 30494 11330 30546 11342
rect 34190 11330 34242 11342
rect 44606 11330 44658 11342
rect 45726 11394 45778 11406
rect 57038 11394 57090 11406
rect 50978 11342 50990 11394
rect 51042 11342 51054 11394
rect 54002 11342 54014 11394
rect 54066 11342 54078 11394
rect 54898 11342 54910 11394
rect 54962 11342 54974 11394
rect 55346 11342 55358 11394
rect 55410 11342 55422 11394
rect 45726 11330 45778 11342
rect 57038 11330 57090 11342
rect 6078 11282 6130 11294
rect 6078 11218 6130 11230
rect 6974 11282 7026 11294
rect 6974 11218 7026 11230
rect 8542 11282 8594 11294
rect 8542 11218 8594 11230
rect 9662 11282 9714 11294
rect 9662 11218 9714 11230
rect 18286 11282 18338 11294
rect 18286 11218 18338 11230
rect 22766 11282 22818 11294
rect 22766 11218 22818 11230
rect 25902 11282 25954 11294
rect 25902 11218 25954 11230
rect 26014 11282 26066 11294
rect 26014 11218 26066 11230
rect 26126 11282 26178 11294
rect 26126 11218 26178 11230
rect 27134 11282 27186 11294
rect 27134 11218 27186 11230
rect 32174 11282 32226 11294
rect 38110 11282 38162 11294
rect 43038 11282 43090 11294
rect 35634 11230 35646 11282
rect 35698 11230 35710 11282
rect 35858 11230 35870 11282
rect 35922 11230 35934 11282
rect 40114 11230 40126 11282
rect 40178 11230 40190 11282
rect 32174 11218 32226 11230
rect 38110 11218 38162 11230
rect 43038 11218 43090 11230
rect 44718 11282 44770 11294
rect 44718 11218 44770 11230
rect 47070 11282 47122 11294
rect 47070 11218 47122 11230
rect 51662 11282 51714 11294
rect 56590 11282 56642 11294
rect 54114 11230 54126 11282
rect 54178 11230 54190 11282
rect 54674 11230 54686 11282
rect 54738 11230 54750 11282
rect 51662 11218 51714 11230
rect 56590 11218 56642 11230
rect 14926 11170 14978 11182
rect 14926 11106 14978 11118
rect 24222 11170 24274 11182
rect 24222 11106 24274 11118
rect 24782 11170 24834 11182
rect 24782 11106 24834 11118
rect 25006 11170 25058 11182
rect 25006 11106 25058 11118
rect 27246 11170 27298 11182
rect 27246 11106 27298 11118
rect 27806 11170 27858 11182
rect 27806 11106 27858 11118
rect 28926 11170 28978 11182
rect 28926 11106 28978 11118
rect 31054 11170 31106 11182
rect 31054 11106 31106 11118
rect 33966 11170 34018 11182
rect 33966 11106 34018 11118
rect 34078 11170 34130 11182
rect 34078 11106 34130 11118
rect 34974 11170 35026 11182
rect 42926 11170 42978 11182
rect 46622 11170 46674 11182
rect 40338 11118 40350 11170
rect 40402 11118 40414 11170
rect 46050 11118 46062 11170
rect 46114 11118 46126 11170
rect 34974 11106 35026 11118
rect 42926 11106 42978 11118
rect 46622 11106 46674 11118
rect 46734 11170 46786 11182
rect 46734 11106 46786 11118
rect 46846 11170 46898 11182
rect 46846 11106 46898 11118
rect 56366 11170 56418 11182
rect 56366 11106 56418 11118
rect 1344 11002 59024 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 59024 11002
rect 1344 10916 59024 10950
rect 9102 10834 9154 10846
rect 17054 10834 17106 10846
rect 16482 10782 16494 10834
rect 16546 10782 16558 10834
rect 9102 10770 9154 10782
rect 17054 10770 17106 10782
rect 18062 10834 18114 10846
rect 18062 10770 18114 10782
rect 24446 10834 24498 10846
rect 24446 10770 24498 10782
rect 25566 10834 25618 10846
rect 25566 10770 25618 10782
rect 25678 10834 25730 10846
rect 25678 10770 25730 10782
rect 25902 10834 25954 10846
rect 25902 10770 25954 10782
rect 29262 10834 29314 10846
rect 29262 10770 29314 10782
rect 29710 10834 29762 10846
rect 29710 10770 29762 10782
rect 31502 10834 31554 10846
rect 31502 10770 31554 10782
rect 33630 10834 33682 10846
rect 33630 10770 33682 10782
rect 39342 10834 39394 10846
rect 39342 10770 39394 10782
rect 39790 10834 39842 10846
rect 39790 10770 39842 10782
rect 40686 10834 40738 10846
rect 40686 10770 40738 10782
rect 41582 10834 41634 10846
rect 41582 10770 41634 10782
rect 42366 10834 42418 10846
rect 42366 10770 42418 10782
rect 42702 10834 42754 10846
rect 42702 10770 42754 10782
rect 44158 10834 44210 10846
rect 44158 10770 44210 10782
rect 48750 10834 48802 10846
rect 48750 10770 48802 10782
rect 49758 10834 49810 10846
rect 49758 10770 49810 10782
rect 9998 10722 10050 10734
rect 9998 10658 10050 10670
rect 10334 10722 10386 10734
rect 10334 10658 10386 10670
rect 19630 10722 19682 10734
rect 19630 10658 19682 10670
rect 22094 10722 22146 10734
rect 22094 10658 22146 10670
rect 23774 10722 23826 10734
rect 23774 10658 23826 10670
rect 26126 10722 26178 10734
rect 26126 10658 26178 10670
rect 26798 10722 26850 10734
rect 26798 10658 26850 10670
rect 32622 10722 32674 10734
rect 32622 10658 32674 10670
rect 34302 10722 34354 10734
rect 34302 10658 34354 10670
rect 43710 10722 43762 10734
rect 43710 10658 43762 10670
rect 43934 10722 43986 10734
rect 43934 10658 43986 10670
rect 49534 10722 49586 10734
rect 49534 10658 49586 10670
rect 55806 10722 55858 10734
rect 55806 10658 55858 10670
rect 13582 10610 13634 10622
rect 17614 10610 17666 10622
rect 4834 10558 4846 10610
rect 4898 10558 4910 10610
rect 14018 10558 14030 10610
rect 14082 10558 14094 10610
rect 13582 10546 13634 10558
rect 17614 10546 17666 10558
rect 19966 10610 20018 10622
rect 19966 10546 20018 10558
rect 20526 10610 20578 10622
rect 23662 10610 23714 10622
rect 25006 10610 25058 10622
rect 21186 10558 21198 10610
rect 21250 10558 21262 10610
rect 22642 10558 22654 10610
rect 22706 10558 22718 10610
rect 24658 10558 24670 10610
rect 24722 10558 24734 10610
rect 20526 10546 20578 10558
rect 23662 10546 23714 10558
rect 25006 10546 25058 10558
rect 31390 10610 31442 10622
rect 31390 10546 31442 10558
rect 31614 10610 31666 10622
rect 31614 10546 31666 10558
rect 32062 10610 32114 10622
rect 32062 10546 32114 10558
rect 32510 10610 32562 10622
rect 32510 10546 32562 10558
rect 35086 10610 35138 10622
rect 36542 10610 36594 10622
rect 35298 10558 35310 10610
rect 35362 10558 35374 10610
rect 35086 10546 35138 10558
rect 36542 10546 36594 10558
rect 37550 10610 37602 10622
rect 37550 10546 37602 10558
rect 37774 10610 37826 10622
rect 37774 10546 37826 10558
rect 44270 10610 44322 10622
rect 44270 10546 44322 10558
rect 44718 10610 44770 10622
rect 47406 10610 47458 10622
rect 53118 10610 53170 10622
rect 54798 10610 54850 10622
rect 46610 10558 46622 10610
rect 46674 10558 46686 10610
rect 50978 10558 50990 10610
rect 51042 10558 51054 10610
rect 51314 10558 51326 10610
rect 51378 10558 51390 10610
rect 53330 10558 53342 10610
rect 53394 10558 53406 10610
rect 44718 10546 44770 10558
rect 47406 10546 47458 10558
rect 53118 10546 53170 10558
rect 54798 10546 54850 10558
rect 55694 10610 55746 10622
rect 55694 10546 55746 10558
rect 56030 10610 56082 10622
rect 56030 10546 56082 10558
rect 18510 10498 18562 10510
rect 24334 10498 24386 10510
rect 27470 10498 27522 10510
rect 5058 10446 5070 10498
rect 5122 10446 5134 10498
rect 21410 10446 21422 10498
rect 21474 10446 21486 10498
rect 22978 10446 22990 10498
rect 23042 10446 23054 10498
rect 26674 10446 26686 10498
rect 26738 10446 26750 10498
rect 18510 10434 18562 10446
rect 24334 10434 24386 10446
rect 27470 10434 27522 10446
rect 27918 10498 27970 10510
rect 27918 10434 27970 10446
rect 28478 10498 28530 10510
rect 28478 10434 28530 10446
rect 28814 10498 28866 10510
rect 28814 10434 28866 10446
rect 30158 10498 30210 10510
rect 30158 10434 30210 10446
rect 30718 10498 30770 10510
rect 30718 10434 30770 10446
rect 35982 10498 36034 10510
rect 35982 10434 36034 10446
rect 40238 10498 40290 10510
rect 40238 10434 40290 10446
rect 43150 10498 43202 10510
rect 43150 10434 43202 10446
rect 45166 10498 45218 10510
rect 45166 10434 45218 10446
rect 45614 10498 45666 10510
rect 51550 10498 51602 10510
rect 47058 10446 47070 10498
rect 47122 10446 47134 10498
rect 45614 10434 45666 10446
rect 51550 10434 51602 10446
rect 54014 10498 54066 10510
rect 54014 10434 54066 10446
rect 54574 10498 54626 10510
rect 54574 10434 54626 10446
rect 27022 10386 27074 10398
rect 5282 10334 5294 10386
rect 5346 10334 5358 10386
rect 27022 10322 27074 10334
rect 32622 10386 32674 10398
rect 32622 10322 32674 10334
rect 34078 10386 34130 10398
rect 34078 10322 34130 10334
rect 34414 10386 34466 10398
rect 49870 10386 49922 10398
rect 38098 10334 38110 10386
rect 38162 10334 38174 10386
rect 39218 10334 39230 10386
rect 39282 10383 39294 10386
rect 40226 10383 40238 10386
rect 39282 10337 40238 10383
rect 39282 10334 39294 10337
rect 40226 10334 40238 10337
rect 40290 10334 40302 10386
rect 34414 10322 34466 10334
rect 49870 10322 49922 10334
rect 55134 10386 55186 10398
rect 55134 10322 55186 10334
rect 1344 10218 59024 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 59024 10218
rect 1344 10132 59024 10166
rect 13022 10050 13074 10062
rect 13022 9986 13074 9998
rect 22990 10050 23042 10062
rect 26686 10050 26738 10062
rect 26338 9998 26350 10050
rect 26402 9998 26414 10050
rect 22990 9986 23042 9998
rect 26686 9986 26738 9998
rect 27358 10050 27410 10062
rect 27358 9986 27410 9998
rect 29710 10050 29762 10062
rect 29710 9986 29762 9998
rect 38894 10050 38946 10062
rect 38894 9986 38946 9998
rect 44270 10050 44322 10062
rect 44270 9986 44322 9998
rect 46286 10050 46338 10062
rect 46286 9986 46338 9998
rect 46622 10050 46674 10062
rect 46622 9986 46674 9998
rect 55470 10050 55522 10062
rect 55470 9986 55522 9998
rect 14030 9938 14082 9950
rect 8418 9886 8430 9938
rect 8482 9886 8494 9938
rect 14030 9874 14082 9886
rect 19294 9938 19346 9950
rect 23550 9938 23602 9950
rect 22754 9886 22766 9938
rect 22818 9886 22830 9938
rect 19294 9874 19346 9886
rect 23550 9874 23602 9886
rect 28590 9938 28642 9950
rect 28590 9874 28642 9886
rect 33518 9938 33570 9950
rect 48302 9938 48354 9950
rect 51662 9938 51714 9950
rect 57486 9938 57538 9950
rect 43250 9886 43262 9938
rect 43314 9886 43326 9938
rect 49410 9886 49422 9938
rect 49474 9886 49486 9938
rect 56802 9886 56814 9938
rect 56866 9886 56878 9938
rect 33518 9874 33570 9886
rect 48302 9874 48354 9886
rect 51662 9874 51714 9886
rect 57486 9874 57538 9886
rect 4846 9826 4898 9838
rect 4274 9774 4286 9826
rect 4338 9774 4350 9826
rect 4846 9762 4898 9774
rect 9550 9826 9602 9838
rect 15486 9826 15538 9838
rect 25790 9826 25842 9838
rect 9874 9774 9886 9826
rect 9938 9774 9950 9826
rect 15922 9774 15934 9826
rect 15986 9774 15998 9826
rect 22642 9774 22654 9826
rect 22706 9774 22718 9826
rect 9550 9762 9602 9774
rect 15486 9762 15538 9774
rect 25790 9762 25842 9774
rect 26910 9826 26962 9838
rect 26910 9762 26962 9774
rect 28030 9826 28082 9838
rect 28030 9762 28082 9774
rect 29598 9826 29650 9838
rect 34750 9826 34802 9838
rect 31490 9774 31502 9826
rect 31554 9774 31566 9826
rect 32162 9774 32174 9826
rect 32226 9774 32238 9826
rect 29598 9762 29650 9774
rect 34750 9762 34802 9774
rect 35086 9826 35138 9838
rect 35086 9762 35138 9774
rect 35310 9826 35362 9838
rect 35310 9762 35362 9774
rect 37886 9826 37938 9838
rect 37886 9762 37938 9774
rect 37998 9826 38050 9838
rect 40014 9826 40066 9838
rect 39218 9774 39230 9826
rect 39282 9774 39294 9826
rect 37998 9762 38050 9774
rect 40014 9762 40066 9774
rect 40462 9826 40514 9838
rect 40462 9762 40514 9774
rect 40910 9826 40962 9838
rect 40910 9762 40962 9774
rect 41134 9826 41186 9838
rect 47070 9826 47122 9838
rect 42018 9774 42030 9826
rect 42082 9774 42094 9826
rect 43026 9774 43038 9826
rect 43090 9774 43102 9826
rect 44594 9774 44606 9826
rect 44658 9774 44670 9826
rect 46610 9774 46622 9826
rect 46674 9774 46686 9826
rect 49186 9774 49198 9826
rect 49250 9774 49262 9826
rect 54338 9774 54350 9826
rect 54402 9774 54414 9826
rect 54562 9774 54574 9826
rect 54626 9774 54638 9826
rect 55234 9774 55246 9826
rect 55298 9774 55310 9826
rect 56914 9774 56926 9826
rect 56978 9774 56990 9826
rect 41134 9762 41186 9774
rect 47070 9762 47122 9774
rect 4958 9714 5010 9726
rect 4958 9650 5010 9662
rect 5742 9714 5794 9726
rect 5742 9650 5794 9662
rect 18958 9714 19010 9726
rect 18958 9650 19010 9662
rect 27694 9714 27746 9726
rect 27694 9650 27746 9662
rect 28478 9714 28530 9726
rect 34078 9714 34130 9726
rect 30930 9662 30942 9714
rect 30994 9662 31006 9714
rect 28478 9650 28530 9662
rect 34078 9650 34130 9662
rect 34974 9714 35026 9726
rect 34974 9650 35026 9662
rect 37550 9714 37602 9726
rect 37550 9650 37602 9662
rect 41694 9714 41746 9726
rect 41694 9650 41746 9662
rect 43710 9714 43762 9726
rect 43710 9650 43762 9662
rect 49870 9714 49922 9726
rect 49870 9650 49922 9662
rect 6078 9602 6130 9614
rect 6078 9538 6130 9550
rect 8878 9602 8930 9614
rect 13582 9602 13634 9614
rect 12450 9550 12462 9602
rect 12514 9550 12526 9602
rect 8878 9538 8930 9550
rect 13582 9538 13634 9550
rect 14814 9602 14866 9614
rect 25118 9602 25170 9614
rect 18386 9550 18398 9602
rect 18450 9550 18462 9602
rect 14814 9538 14866 9550
rect 25118 9538 25170 9550
rect 27470 9602 27522 9614
rect 27470 9538 27522 9550
rect 28702 9602 28754 9614
rect 28702 9538 28754 9550
rect 29710 9602 29762 9614
rect 37774 9602 37826 9614
rect 32722 9550 32734 9602
rect 32786 9550 32798 9602
rect 29710 9538 29762 9550
rect 37774 9538 37826 9550
rect 39006 9602 39058 9614
rect 39006 9538 39058 9550
rect 40798 9602 40850 9614
rect 40798 9538 40850 9550
rect 41806 9602 41858 9614
rect 41806 9538 41858 9550
rect 44382 9602 44434 9614
rect 44382 9538 44434 9550
rect 45390 9602 45442 9614
rect 45390 9538 45442 9550
rect 51550 9602 51602 9614
rect 51550 9538 51602 9550
rect 1344 9434 59024 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 59024 9434
rect 1344 9348 59024 9382
rect 4398 9266 4450 9278
rect 4398 9202 4450 9214
rect 4846 9266 4898 9278
rect 8990 9266 9042 9278
rect 8306 9214 8318 9266
rect 8370 9214 8382 9266
rect 4846 9202 4898 9214
rect 8990 9202 9042 9214
rect 13022 9266 13074 9278
rect 21310 9266 21362 9278
rect 14018 9214 14030 9266
rect 14082 9214 14094 9266
rect 13022 9202 13074 9214
rect 21310 9202 21362 9214
rect 21870 9266 21922 9278
rect 21870 9202 21922 9214
rect 22654 9266 22706 9278
rect 22654 9202 22706 9214
rect 23550 9266 23602 9278
rect 23550 9202 23602 9214
rect 25678 9266 25730 9278
rect 25678 9202 25730 9214
rect 26238 9266 26290 9278
rect 26238 9202 26290 9214
rect 26686 9266 26738 9278
rect 26686 9202 26738 9214
rect 27134 9266 27186 9278
rect 27134 9202 27186 9214
rect 31054 9266 31106 9278
rect 31054 9202 31106 9214
rect 31726 9266 31778 9278
rect 31726 9202 31778 9214
rect 33742 9266 33794 9278
rect 33742 9202 33794 9214
rect 34638 9266 34690 9278
rect 34638 9202 34690 9214
rect 34974 9266 35026 9278
rect 34974 9202 35026 9214
rect 35646 9266 35698 9278
rect 35646 9202 35698 9214
rect 36318 9266 36370 9278
rect 36318 9202 36370 9214
rect 42030 9266 42082 9278
rect 42030 9202 42082 9214
rect 42254 9266 42306 9278
rect 42254 9202 42306 9214
rect 43150 9266 43202 9278
rect 43150 9202 43202 9214
rect 45502 9266 45554 9278
rect 45502 9202 45554 9214
rect 54686 9266 54738 9278
rect 54686 9202 54738 9214
rect 57598 9266 57650 9278
rect 57598 9202 57650 9214
rect 10110 9154 10162 9166
rect 10110 9090 10162 9102
rect 11006 9154 11058 9166
rect 11006 9090 11058 9102
rect 22990 9154 23042 9166
rect 22990 9090 23042 9102
rect 31614 9154 31666 9166
rect 31614 9090 31666 9102
rect 32398 9154 32450 9166
rect 32398 9090 32450 9102
rect 32734 9154 32786 9166
rect 32734 9090 32786 9102
rect 36206 9154 36258 9166
rect 36206 9090 36258 9102
rect 39118 9154 39170 9166
rect 39118 9090 39170 9102
rect 41918 9154 41970 9166
rect 41918 9090 41970 9102
rect 42702 9154 42754 9166
rect 42702 9090 42754 9102
rect 43822 9154 43874 9166
rect 43822 9090 43874 9102
rect 44494 9154 44546 9166
rect 44494 9090 44546 9102
rect 44718 9154 44770 9166
rect 44718 9090 44770 9102
rect 44942 9154 44994 9166
rect 44942 9090 44994 9102
rect 45054 9154 45106 9166
rect 45054 9090 45106 9102
rect 46286 9154 46338 9166
rect 46286 9090 46338 9102
rect 46510 9154 46562 9166
rect 46510 9090 46562 9102
rect 47406 9154 47458 9166
rect 47406 9090 47458 9102
rect 47630 9154 47682 9166
rect 47630 9090 47682 9102
rect 49534 9154 49586 9166
rect 49534 9090 49586 9102
rect 49758 9154 49810 9166
rect 49758 9090 49810 9102
rect 50430 9154 50482 9166
rect 50430 9090 50482 9102
rect 51662 9154 51714 9166
rect 51662 9090 51714 9102
rect 53678 9154 53730 9166
rect 53678 9090 53730 9102
rect 54462 9154 54514 9166
rect 54462 9090 54514 9102
rect 54798 9154 54850 9166
rect 54798 9090 54850 9102
rect 57486 9154 57538 9166
rect 57698 9102 57710 9154
rect 57762 9102 57774 9154
rect 57486 9090 57538 9102
rect 4286 9042 4338 9054
rect 4286 8978 4338 8990
rect 5518 9042 5570 9054
rect 9774 9042 9826 9054
rect 5954 8990 5966 9042
rect 6018 8990 6030 9042
rect 5518 8978 5570 8990
rect 9774 8978 9826 8990
rect 10558 9042 10610 9054
rect 17054 9042 17106 9054
rect 16482 8990 16494 9042
rect 16546 8990 16558 9042
rect 10558 8978 10610 8990
rect 17054 8978 17106 8990
rect 21646 9042 21698 9054
rect 21646 8978 21698 8990
rect 21982 9042 22034 9054
rect 21982 8978 22034 8990
rect 22542 9042 22594 9054
rect 22542 8978 22594 8990
rect 22766 9042 22818 9054
rect 22766 8978 22818 8990
rect 27582 9042 27634 9054
rect 37886 9042 37938 9054
rect 40686 9042 40738 9054
rect 28130 8990 28142 9042
rect 28194 8990 28206 9042
rect 30034 8990 30046 9042
rect 30098 8990 30110 9042
rect 30258 8990 30270 9042
rect 30322 8990 30334 9042
rect 37426 8990 37438 9042
rect 37490 8990 37502 9042
rect 38770 8990 38782 9042
rect 38834 8990 38846 9042
rect 39218 8990 39230 9042
rect 39282 9039 39294 9042
rect 39554 9039 39566 9042
rect 39282 8993 39566 9039
rect 39282 8990 39294 8993
rect 39554 8990 39566 8993
rect 39618 8990 39630 9042
rect 40450 8990 40462 9042
rect 40514 8990 40526 9042
rect 27582 8978 27634 8990
rect 37886 8978 37938 8990
rect 40686 8978 40738 8990
rect 42926 9042 42978 9054
rect 42926 8978 42978 8990
rect 47182 9042 47234 9054
rect 47182 8978 47234 8990
rect 47742 9042 47794 9054
rect 47742 8978 47794 8990
rect 50654 9042 50706 9054
rect 50654 8978 50706 8990
rect 51550 9042 51602 9054
rect 51550 8978 51602 8990
rect 51886 9042 51938 9054
rect 51886 8978 51938 8990
rect 52782 9042 52834 9054
rect 54238 9042 54290 9054
rect 52994 8990 53006 9042
rect 53058 8990 53070 9042
rect 56018 8990 56030 9042
rect 56082 8990 56094 9042
rect 58034 8990 58046 9042
rect 58098 8990 58110 9042
rect 52782 8978 52834 8990
rect 54238 8978 54290 8990
rect 13358 8930 13410 8942
rect 13358 8866 13410 8878
rect 17614 8930 17666 8942
rect 17614 8866 17666 8878
rect 18062 8930 18114 8942
rect 18062 8866 18114 8878
rect 18622 8930 18674 8942
rect 18622 8866 18674 8878
rect 23998 8930 24050 8942
rect 23998 8866 24050 8878
rect 29150 8930 29202 8942
rect 31838 8930 31890 8942
rect 39006 8930 39058 8942
rect 29810 8878 29822 8930
rect 29874 8878 29886 8930
rect 37538 8878 37550 8930
rect 37602 8878 37614 8930
rect 29150 8866 29202 8878
rect 31838 8866 31890 8878
rect 39006 8866 39058 8878
rect 39790 8930 39842 8942
rect 39790 8866 39842 8878
rect 42814 8930 42866 8942
rect 56702 8930 56754 8942
rect 46610 8878 46622 8930
rect 46674 8878 46686 8930
rect 56242 8878 56254 8930
rect 56306 8878 56318 8930
rect 42814 8866 42866 8878
rect 56702 8866 56754 8878
rect 28142 8818 28194 8830
rect 28142 8754 28194 8766
rect 28478 8818 28530 8830
rect 28478 8754 28530 8766
rect 43934 8818 43986 8830
rect 43934 8754 43986 8766
rect 49870 8818 49922 8830
rect 49870 8754 49922 8766
rect 50990 8818 51042 8830
rect 50990 8754 51042 8766
rect 57934 8818 57986 8830
rect 57934 8754 57986 8766
rect 1344 8650 59024 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 59024 8650
rect 1344 8564 59024 8598
rect 29710 8482 29762 8494
rect 29710 8418 29762 8430
rect 39566 8482 39618 8494
rect 39566 8418 39618 8430
rect 55022 8482 55074 8494
rect 56914 8430 56926 8482
rect 56978 8430 56990 8482
rect 55022 8418 55074 8430
rect 6750 8370 6802 8382
rect 13022 8370 13074 8382
rect 8082 8318 8094 8370
rect 8146 8318 8158 8370
rect 6750 8306 6802 8318
rect 13022 8306 13074 8318
rect 19070 8370 19122 8382
rect 19070 8306 19122 8318
rect 22878 8370 22930 8382
rect 22878 8306 22930 8318
rect 25454 8370 25506 8382
rect 25454 8306 25506 8318
rect 32286 8370 32338 8382
rect 32286 8306 32338 8318
rect 33294 8370 33346 8382
rect 33294 8306 33346 8318
rect 34078 8370 34130 8382
rect 41582 8370 41634 8382
rect 35186 8318 35198 8370
rect 35250 8318 35262 8370
rect 38098 8318 38110 8370
rect 38162 8318 38174 8370
rect 34078 8306 34130 8318
rect 41582 8306 41634 8318
rect 43150 8370 43202 8382
rect 47058 8318 47070 8370
rect 47122 8318 47134 8370
rect 56578 8318 56590 8370
rect 56642 8318 56654 8370
rect 43150 8306 43202 8318
rect 9550 8258 9602 8270
rect 15038 8258 15090 8270
rect 18622 8258 18674 8270
rect 7746 8206 7758 8258
rect 7810 8206 7822 8258
rect 9874 8206 9886 8258
rect 9938 8206 9950 8258
rect 15362 8206 15374 8258
rect 15426 8206 15438 8258
rect 9550 8194 9602 8206
rect 15038 8194 15090 8206
rect 18622 8194 18674 8206
rect 22654 8258 22706 8270
rect 22654 8194 22706 8206
rect 23326 8258 23378 8270
rect 26014 8258 26066 8270
rect 24210 8206 24222 8258
rect 24274 8206 24286 8258
rect 24658 8206 24670 8258
rect 24722 8206 24734 8258
rect 23326 8194 23378 8206
rect 26014 8194 26066 8206
rect 26686 8258 26738 8270
rect 28254 8258 28306 8270
rect 27794 8206 27806 8258
rect 27858 8206 27870 8258
rect 26686 8194 26738 8206
rect 28254 8194 28306 8206
rect 29822 8258 29874 8270
rect 29822 8194 29874 8206
rect 31950 8258 32002 8270
rect 31950 8194 32002 8206
rect 32174 8258 32226 8270
rect 32174 8194 32226 8206
rect 32510 8258 32562 8270
rect 32510 8194 32562 8206
rect 34302 8258 34354 8270
rect 34302 8194 34354 8206
rect 35534 8258 35586 8270
rect 35534 8194 35586 8206
rect 35982 8258 36034 8270
rect 39118 8258 39170 8270
rect 40798 8258 40850 8270
rect 37874 8206 37886 8258
rect 37938 8206 37950 8258
rect 39330 8206 39342 8258
rect 39394 8206 39406 8258
rect 39666 8206 39678 8258
rect 39730 8206 39742 8258
rect 35982 8194 36034 8206
rect 39118 8194 39170 8206
rect 40798 8194 40850 8206
rect 42478 8258 42530 8270
rect 42478 8194 42530 8206
rect 42702 8258 42754 8270
rect 42702 8194 42754 8206
rect 42926 8258 42978 8270
rect 44606 8258 44658 8270
rect 52670 8258 52722 8270
rect 44146 8206 44158 8258
rect 44210 8206 44222 8258
rect 46946 8206 46958 8258
rect 47010 8206 47022 8258
rect 49074 8206 49086 8258
rect 49138 8206 49150 8258
rect 49522 8206 49534 8258
rect 49586 8206 49598 8258
rect 51090 8206 51102 8258
rect 51154 8206 51166 8258
rect 52098 8206 52110 8258
rect 52162 8206 52174 8258
rect 53442 8206 53454 8258
rect 53506 8206 53518 8258
rect 54226 8206 54238 8258
rect 54290 8206 54302 8258
rect 54674 8206 54686 8258
rect 54738 8206 54750 8258
rect 55906 8206 55918 8258
rect 55970 8206 55982 8258
rect 56690 8206 56702 8258
rect 56754 8206 56766 8258
rect 42926 8194 42978 8206
rect 44606 8194 44658 8206
rect 52670 8194 52722 8206
rect 8206 8146 8258 8158
rect 8206 8082 8258 8094
rect 21982 8146 22034 8158
rect 21982 8082 22034 8094
rect 23102 8146 23154 8158
rect 23102 8082 23154 8094
rect 23998 8146 24050 8158
rect 23998 8082 24050 8094
rect 26238 8146 26290 8158
rect 30606 8146 30658 8158
rect 27122 8094 27134 8146
rect 27186 8094 27198 8146
rect 28802 8094 28814 8146
rect 28866 8094 28878 8146
rect 26238 8082 26290 8094
rect 30606 8082 30658 8094
rect 35310 8146 35362 8158
rect 35310 8082 35362 8094
rect 38558 8146 38610 8158
rect 38558 8082 38610 8094
rect 44718 8146 44770 8158
rect 44718 8082 44770 8094
rect 47854 8146 47906 8158
rect 47854 8082 47906 8094
rect 49758 8146 49810 8158
rect 53678 8146 53730 8158
rect 50754 8094 50766 8146
rect 50818 8094 50830 8146
rect 49758 8082 49810 8094
rect 53678 8082 53730 8094
rect 55582 8146 55634 8158
rect 55582 8082 55634 8094
rect 7198 8034 7250 8046
rect 7198 7970 7250 7982
rect 7982 8034 8034 8046
rect 7982 7970 8034 7982
rect 8654 8034 8706 8046
rect 13582 8034 13634 8046
rect 12450 7982 12462 8034
rect 12514 7982 12526 8034
rect 8654 7970 8706 7982
rect 13582 7970 13634 7982
rect 14030 8034 14082 8046
rect 19518 8034 19570 8046
rect 17938 7982 17950 8034
rect 18002 7982 18014 8034
rect 14030 7970 14082 7982
rect 19518 7970 19570 7982
rect 20862 8034 20914 8046
rect 20862 7970 20914 7982
rect 21646 8034 21698 8046
rect 21646 7970 21698 7982
rect 26350 8034 26402 8046
rect 29710 8034 29762 8046
rect 27234 7982 27246 8034
rect 27298 7982 27310 8034
rect 26350 7970 26402 7982
rect 29710 7970 29762 7982
rect 30270 8034 30322 8046
rect 30270 7970 30322 7982
rect 30494 8034 30546 8046
rect 30494 7970 30546 7982
rect 31166 8034 31218 8046
rect 31166 7970 31218 7982
rect 32846 8034 32898 8046
rect 39902 8034 39954 8046
rect 34626 7982 34638 8034
rect 34690 7982 34702 8034
rect 32846 7970 32898 7982
rect 39902 7970 39954 7982
rect 40574 8034 40626 8046
rect 40574 7970 40626 7982
rect 40910 8034 40962 8046
rect 40910 7970 40962 7982
rect 41022 8034 41074 8046
rect 41022 7970 41074 7982
rect 42590 8034 42642 8046
rect 42590 7970 42642 7982
rect 45950 8034 46002 8046
rect 45950 7970 46002 7982
rect 57710 8034 57762 8046
rect 57710 7970 57762 7982
rect 1344 7866 59024 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 59024 7866
rect 1344 7780 59024 7814
rect 13358 7698 13410 7710
rect 12786 7646 12798 7698
rect 12850 7646 12862 7698
rect 13358 7634 13410 7646
rect 18734 7698 18786 7710
rect 18734 7634 18786 7646
rect 19182 7698 19234 7710
rect 22878 7698 22930 7710
rect 22082 7646 22094 7698
rect 22146 7646 22158 7698
rect 19182 7634 19234 7646
rect 22878 7634 22930 7646
rect 27470 7698 27522 7710
rect 27470 7634 27522 7646
rect 33630 7698 33682 7710
rect 41582 7698 41634 7710
rect 39554 7646 39566 7698
rect 39618 7646 39630 7698
rect 33630 7634 33682 7646
rect 41582 7634 41634 7646
rect 42030 7698 42082 7710
rect 42030 7634 42082 7646
rect 44494 7698 44546 7710
rect 44494 7634 44546 7646
rect 53230 7698 53282 7710
rect 53230 7634 53282 7646
rect 53454 7698 53506 7710
rect 53454 7634 53506 7646
rect 54462 7698 54514 7710
rect 54462 7634 54514 7646
rect 54686 7698 54738 7710
rect 55906 7646 55918 7698
rect 55970 7646 55982 7698
rect 54686 7634 54738 7646
rect 6190 7586 6242 7598
rect 6190 7522 6242 7534
rect 8990 7586 9042 7598
rect 22990 7586 23042 7598
rect 20850 7534 20862 7586
rect 20914 7534 20926 7586
rect 22194 7534 22206 7586
rect 22258 7534 22270 7586
rect 8990 7522 9042 7534
rect 22990 7522 23042 7534
rect 23438 7586 23490 7598
rect 23438 7522 23490 7534
rect 24670 7586 24722 7598
rect 24670 7522 24722 7534
rect 24894 7586 24946 7598
rect 24894 7522 24946 7534
rect 25678 7586 25730 7598
rect 25678 7522 25730 7534
rect 25790 7586 25842 7598
rect 25790 7522 25842 7534
rect 27358 7586 27410 7598
rect 27358 7522 27410 7534
rect 27582 7586 27634 7598
rect 27582 7522 27634 7534
rect 28254 7586 28306 7598
rect 28254 7522 28306 7534
rect 34750 7586 34802 7598
rect 34750 7522 34802 7534
rect 34974 7586 35026 7598
rect 34974 7522 35026 7534
rect 37326 7586 37378 7598
rect 37326 7522 37378 7534
rect 45390 7586 45442 7598
rect 45390 7522 45442 7534
rect 46958 7586 47010 7598
rect 53118 7586 53170 7598
rect 50642 7534 50654 7586
rect 50706 7534 50718 7586
rect 46958 7522 47010 7534
rect 53118 7522 53170 7534
rect 54350 7586 54402 7598
rect 54350 7522 54402 7534
rect 5854 7474 5906 7486
rect 9662 7474 9714 7486
rect 24222 7474 24274 7486
rect 8306 7422 8318 7474
rect 8370 7422 8382 7474
rect 10210 7422 10222 7474
rect 10274 7422 10286 7474
rect 21074 7422 21086 7474
rect 21138 7422 21150 7474
rect 23202 7422 23214 7474
rect 23266 7422 23278 7474
rect 5854 7410 5906 7422
rect 9662 7410 9714 7422
rect 24222 7410 24274 7422
rect 24446 7474 24498 7486
rect 28814 7474 28866 7486
rect 26002 7422 26014 7474
rect 26066 7422 26078 7474
rect 24446 7410 24498 7422
rect 28814 7410 28866 7422
rect 29822 7474 29874 7486
rect 32622 7474 32674 7486
rect 39902 7474 39954 7486
rect 31602 7422 31614 7474
rect 31666 7422 31678 7474
rect 37650 7422 37662 7474
rect 37714 7422 37726 7474
rect 29822 7410 29874 7422
rect 32622 7410 32674 7422
rect 39902 7410 39954 7422
rect 40126 7474 40178 7486
rect 46062 7474 46114 7486
rect 55358 7474 55410 7486
rect 43138 7422 43150 7474
rect 43202 7422 43214 7474
rect 46498 7422 46510 7474
rect 46562 7422 46574 7474
rect 49970 7422 49982 7474
rect 50034 7422 50046 7474
rect 50866 7422 50878 7474
rect 50930 7422 50942 7474
rect 40126 7410 40178 7422
rect 46062 7410 46114 7422
rect 55358 7410 55410 7422
rect 55582 7474 55634 7486
rect 55582 7410 55634 7422
rect 5182 7362 5234 7374
rect 13694 7362 13746 7374
rect 8082 7310 8094 7362
rect 8146 7310 8158 7362
rect 5182 7298 5234 7310
rect 13694 7298 13746 7310
rect 19630 7362 19682 7374
rect 19630 7298 19682 7310
rect 26798 7362 26850 7374
rect 26798 7298 26850 7310
rect 30270 7362 30322 7374
rect 32174 7362 32226 7374
rect 31266 7310 31278 7362
rect 31330 7310 31342 7362
rect 30270 7298 30322 7310
rect 32174 7298 32226 7310
rect 42478 7362 42530 7374
rect 43934 7362 43986 7374
rect 53790 7362 53842 7374
rect 42914 7310 42926 7362
rect 42978 7310 42990 7362
rect 50978 7310 50990 7362
rect 51042 7310 51054 7362
rect 42478 7298 42530 7310
rect 43934 7298 43986 7310
rect 53790 7298 53842 7310
rect 29934 7250 29986 7262
rect 29934 7186 29986 7198
rect 30158 7250 30210 7262
rect 30158 7186 30210 7198
rect 34638 7250 34690 7262
rect 34638 7186 34690 7198
rect 37662 7250 37714 7262
rect 37662 7186 37714 7198
rect 1344 7082 59024 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 59024 7082
rect 1344 6996 59024 7030
rect 18734 6914 18786 6926
rect 18734 6850 18786 6862
rect 31838 6914 31890 6926
rect 31838 6850 31890 6862
rect 13582 6802 13634 6814
rect 28030 6802 28082 6814
rect 27010 6750 27022 6802
rect 27074 6750 27086 6802
rect 13582 6738 13634 6750
rect 28030 6738 28082 6750
rect 30718 6802 30770 6814
rect 30718 6738 30770 6750
rect 32846 6802 32898 6814
rect 43822 6802 43874 6814
rect 34626 6750 34638 6802
rect 34690 6750 34702 6802
rect 32846 6738 32898 6750
rect 43822 6738 43874 6750
rect 7646 6690 7698 6702
rect 6738 6638 6750 6690
rect 6802 6638 6814 6690
rect 7646 6626 7698 6638
rect 8542 6690 8594 6702
rect 8542 6626 8594 6638
rect 8878 6690 8930 6702
rect 8878 6626 8930 6638
rect 9550 6690 9602 6702
rect 15038 6690 15090 6702
rect 20638 6690 20690 6702
rect 9986 6638 9998 6690
rect 10050 6638 10062 6690
rect 15698 6638 15710 6690
rect 15762 6638 15774 6690
rect 19618 6638 19630 6690
rect 19682 6638 19694 6690
rect 9550 6626 9602 6638
rect 15038 6626 15090 6638
rect 20638 6626 20690 6638
rect 22542 6690 22594 6702
rect 22542 6626 22594 6638
rect 24670 6690 24722 6702
rect 24670 6626 24722 6638
rect 25790 6690 25842 6702
rect 26686 6690 26738 6702
rect 26450 6638 26462 6690
rect 26514 6638 26526 6690
rect 25790 6626 25842 6638
rect 26686 6626 26738 6638
rect 28590 6690 28642 6702
rect 28590 6626 28642 6638
rect 31614 6690 31666 6702
rect 35982 6690 36034 6702
rect 32162 6638 32174 6690
rect 32226 6638 32238 6690
rect 34850 6638 34862 6690
rect 34914 6638 34926 6690
rect 31614 6626 31666 6638
rect 35982 6626 36034 6638
rect 4734 6578 4786 6590
rect 4734 6514 4786 6526
rect 4846 6578 4898 6590
rect 4846 6514 4898 6526
rect 20302 6578 20354 6590
rect 20302 6514 20354 6526
rect 21982 6578 22034 6590
rect 21982 6514 22034 6526
rect 23998 6578 24050 6590
rect 23998 6514 24050 6526
rect 24222 6578 24274 6590
rect 24222 6514 24274 6526
rect 27582 6578 27634 6590
rect 27582 6514 27634 6526
rect 28702 6578 28754 6590
rect 28702 6514 28754 6526
rect 35534 6578 35586 6590
rect 35534 6514 35586 6526
rect 5070 6466 5122 6478
rect 5070 6402 5122 6414
rect 5630 6466 5682 6478
rect 5630 6402 5682 6414
rect 6526 6466 6578 6478
rect 6526 6402 6578 6414
rect 7982 6466 8034 6478
rect 13022 6466 13074 6478
rect 12450 6414 12462 6466
rect 12514 6414 12526 6466
rect 7982 6402 8034 6414
rect 13022 6402 13074 6414
rect 14030 6466 14082 6478
rect 14030 6402 14082 6414
rect 14478 6466 14530 6478
rect 19406 6466 19458 6478
rect 17938 6414 17950 6466
rect 18002 6414 18014 6466
rect 14478 6402 14530 6414
rect 19406 6402 19458 6414
rect 21646 6466 21698 6478
rect 21646 6402 21698 6414
rect 22990 6466 23042 6478
rect 22990 6402 23042 6414
rect 23438 6466 23490 6478
rect 23438 6402 23490 6414
rect 24446 6466 24498 6478
rect 24446 6402 24498 6414
rect 25454 6466 25506 6478
rect 25454 6402 25506 6414
rect 29822 6466 29874 6478
rect 29822 6402 29874 6414
rect 30270 6466 30322 6478
rect 30270 6402 30322 6414
rect 32734 6466 32786 6478
rect 32734 6402 32786 6414
rect 32958 6466 33010 6478
rect 32958 6402 33010 6414
rect 33182 6466 33234 6478
rect 33182 6402 33234 6414
rect 33742 6466 33794 6478
rect 33742 6402 33794 6414
rect 45390 6466 45442 6478
rect 45390 6402 45442 6414
rect 55022 6466 55074 6478
rect 55022 6402 55074 6414
rect 55470 6466 55522 6478
rect 55470 6402 55522 6414
rect 1344 6298 59024 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 59024 6298
rect 1344 6212 59024 6246
rect 9102 6130 9154 6142
rect 14366 6130 14418 6142
rect 8306 6078 8318 6130
rect 8370 6078 8382 6130
rect 13234 6078 13246 6130
rect 13298 6078 13310 6130
rect 9102 6066 9154 6078
rect 14366 6066 14418 6078
rect 15150 6130 15202 6142
rect 23326 6130 23378 6142
rect 20514 6078 20526 6130
rect 20578 6078 20590 6130
rect 15150 6066 15202 6078
rect 23326 6066 23378 6078
rect 23550 6130 23602 6142
rect 23550 6066 23602 6078
rect 24446 6130 24498 6142
rect 24446 6066 24498 6078
rect 26014 6130 26066 6142
rect 26014 6066 26066 6078
rect 27022 6130 27074 6142
rect 27022 6066 27074 6078
rect 28590 6130 28642 6142
rect 28590 6066 28642 6078
rect 30606 6130 30658 6142
rect 30606 6066 30658 6078
rect 30830 6130 30882 6142
rect 30830 6066 30882 6078
rect 44494 6130 44546 6142
rect 44494 6066 44546 6078
rect 45278 6130 45330 6142
rect 47954 6078 47966 6130
rect 48018 6078 48030 6130
rect 45278 6066 45330 6078
rect 21982 6018 22034 6030
rect 21982 5954 22034 5966
rect 23102 6018 23154 6030
rect 23102 5954 23154 5966
rect 26462 6018 26514 6030
rect 26462 5954 26514 5966
rect 29038 6018 29090 6030
rect 33630 6018 33682 6030
rect 29362 5966 29374 6018
rect 29426 5966 29438 6018
rect 29038 5954 29090 5966
rect 33630 5954 33682 5966
rect 35534 6018 35586 6030
rect 35534 5954 35586 5966
rect 41582 6018 41634 6030
rect 41582 5954 41634 5966
rect 45502 6018 45554 6030
rect 45502 5954 45554 5966
rect 46286 6018 46338 6030
rect 47058 5966 47070 6018
rect 47122 5966 47134 6018
rect 46286 5954 46338 5966
rect 5630 5906 5682 5918
rect 10110 5906 10162 5918
rect 15710 5906 15762 5918
rect 6066 5854 6078 5906
rect 6130 5854 6142 5906
rect 10770 5854 10782 5906
rect 10834 5854 10846 5906
rect 5630 5842 5682 5854
rect 10110 5842 10162 5854
rect 15710 5842 15762 5854
rect 16158 5906 16210 5918
rect 16158 5842 16210 5854
rect 16718 5906 16770 5918
rect 16718 5842 16770 5854
rect 17614 5906 17666 5918
rect 23662 5906 23714 5918
rect 18274 5854 18286 5906
rect 18338 5854 18350 5906
rect 22194 5854 22206 5906
rect 22258 5854 22270 5906
rect 17614 5842 17666 5854
rect 23662 5842 23714 5854
rect 23998 5906 24050 5918
rect 23998 5842 24050 5854
rect 24558 5906 24610 5918
rect 24558 5842 24610 5854
rect 24670 5906 24722 5918
rect 30942 5906 30994 5918
rect 32398 5906 32450 5918
rect 27906 5854 27918 5906
rect 27970 5854 27982 5906
rect 32050 5854 32062 5906
rect 32114 5854 32126 5906
rect 24670 5842 24722 5854
rect 30942 5842 30994 5854
rect 32398 5842 32450 5854
rect 32510 5906 32562 5918
rect 34862 5906 34914 5918
rect 33842 5854 33854 5906
rect 33906 5854 33918 5906
rect 32510 5842 32562 5854
rect 34862 5842 34914 5854
rect 35086 5906 35138 5918
rect 35086 5842 35138 5854
rect 35310 5906 35362 5918
rect 35310 5842 35362 5854
rect 35758 5906 35810 5918
rect 35758 5842 35810 5854
rect 36542 5906 36594 5918
rect 39454 5906 39506 5918
rect 36978 5854 36990 5906
rect 37042 5854 37054 5906
rect 36542 5842 36594 5854
rect 39454 5842 39506 5854
rect 39678 5906 39730 5918
rect 44606 5906 44658 5918
rect 43810 5854 43822 5906
rect 43874 5854 43886 5906
rect 44370 5854 44382 5906
rect 44434 5854 44446 5906
rect 39678 5842 39730 5854
rect 44606 5842 44658 5854
rect 45166 5906 45218 5918
rect 45166 5842 45218 5854
rect 46174 5906 46226 5918
rect 46946 5854 46958 5906
rect 47010 5854 47022 5906
rect 47842 5854 47854 5906
rect 47906 5854 47918 5906
rect 46174 5842 46226 5854
rect 9662 5794 9714 5806
rect 9662 5730 9714 5742
rect 27694 5794 27746 5806
rect 27694 5730 27746 5742
rect 30270 5794 30322 5806
rect 37438 5794 37490 5806
rect 35634 5742 35646 5794
rect 35698 5742 35710 5794
rect 30270 5730 30322 5742
rect 37438 5730 37490 5742
rect 39230 5794 39282 5806
rect 39230 5730 39282 5742
rect 43262 5794 43314 5806
rect 43262 5730 43314 5742
rect 13806 5682 13858 5694
rect 13806 5618 13858 5630
rect 21310 5682 21362 5694
rect 21310 5618 21362 5630
rect 27582 5682 27634 5694
rect 27582 5618 27634 5630
rect 40126 5682 40178 5694
rect 40126 5618 40178 5630
rect 41806 5682 41858 5694
rect 41806 5618 41858 5630
rect 42142 5682 42194 5694
rect 42142 5618 42194 5630
rect 44158 5682 44210 5694
rect 44158 5618 44210 5630
rect 46286 5682 46338 5694
rect 46286 5618 46338 5630
rect 1344 5514 59024 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 59024 5514
rect 1344 5428 59024 5462
rect 41470 5346 41522 5358
rect 5842 5294 5854 5346
rect 5906 5294 5918 5346
rect 26898 5294 26910 5346
rect 26962 5294 26974 5346
rect 41470 5282 41522 5294
rect 45502 5346 45554 5358
rect 45502 5282 45554 5294
rect 49646 5346 49698 5358
rect 49646 5282 49698 5294
rect 13582 5234 13634 5246
rect 5954 5182 5966 5234
rect 6018 5182 6030 5234
rect 9650 5182 9662 5234
rect 9714 5182 9726 5234
rect 13582 5170 13634 5182
rect 14254 5234 14306 5246
rect 14254 5170 14306 5182
rect 14926 5234 14978 5246
rect 14926 5170 14978 5182
rect 19854 5234 19906 5246
rect 19854 5170 19906 5182
rect 24782 5234 24834 5246
rect 26350 5234 26402 5246
rect 25218 5182 25230 5234
rect 25282 5182 25294 5234
rect 24782 5170 24834 5182
rect 26350 5170 26402 5182
rect 28366 5234 28418 5246
rect 28366 5170 28418 5182
rect 34190 5234 34242 5246
rect 42926 5234 42978 5246
rect 48750 5234 48802 5246
rect 34738 5182 34750 5234
rect 34802 5182 34814 5234
rect 45826 5182 45838 5234
rect 45890 5182 45902 5234
rect 47282 5182 47294 5234
rect 47346 5182 47358 5234
rect 34190 5170 34242 5182
rect 42926 5170 42978 5182
rect 48750 5170 48802 5182
rect 49198 5234 49250 5246
rect 49198 5170 49250 5182
rect 15374 5122 15426 5134
rect 19070 5122 19122 5134
rect 6626 5070 6638 5122
rect 6690 5070 6702 5122
rect 8306 5070 8318 5122
rect 8370 5070 8382 5122
rect 16034 5070 16046 5122
rect 16098 5070 16110 5122
rect 15374 5058 15426 5070
rect 19070 5058 19122 5070
rect 20302 5122 20354 5134
rect 20302 5058 20354 5070
rect 20862 5122 20914 5134
rect 27470 5122 27522 5134
rect 23090 5070 23102 5122
rect 23154 5070 23166 5122
rect 25442 5070 25454 5122
rect 25506 5070 25518 5122
rect 20862 5058 20914 5070
rect 27470 5058 27522 5070
rect 28142 5122 28194 5134
rect 28142 5058 28194 5070
rect 28478 5122 28530 5134
rect 35646 5122 35698 5134
rect 29698 5070 29710 5122
rect 29762 5070 29774 5122
rect 31938 5070 31950 5122
rect 32002 5070 32014 5122
rect 34962 5070 34974 5122
rect 35026 5070 35038 5122
rect 28478 5058 28530 5070
rect 35646 5058 35698 5070
rect 36430 5122 36482 5134
rect 36430 5058 36482 5070
rect 37662 5122 37714 5134
rect 38558 5122 38610 5134
rect 38098 5070 38110 5122
rect 38162 5070 38174 5122
rect 37662 5058 37714 5070
rect 38558 5058 38610 5070
rect 39230 5122 39282 5134
rect 39230 5058 39282 5070
rect 39678 5122 39730 5134
rect 39678 5058 39730 5070
rect 39902 5122 39954 5134
rect 41358 5122 41410 5134
rect 41010 5070 41022 5122
rect 41074 5070 41086 5122
rect 39902 5058 39954 5070
rect 41358 5058 41410 5070
rect 41694 5122 41746 5134
rect 41694 5058 41746 5070
rect 41806 5122 41858 5134
rect 41806 5058 41858 5070
rect 43038 5122 43090 5134
rect 44606 5122 44658 5134
rect 48974 5122 49026 5134
rect 44034 5070 44046 5122
rect 44098 5070 44110 5122
rect 47730 5070 47742 5122
rect 47794 5070 47806 5122
rect 43038 5058 43090 5070
rect 44606 5058 44658 5070
rect 48974 5058 49026 5070
rect 27358 5010 27410 5022
rect 21858 4958 21870 5010
rect 21922 4958 21934 5010
rect 23202 4958 23214 5010
rect 23266 4958 23278 5010
rect 27358 4946 27410 4958
rect 27582 5010 27634 5022
rect 27582 4946 27634 4958
rect 28814 5010 28866 5022
rect 28814 4946 28866 4958
rect 30382 5010 30434 5022
rect 36654 5010 36706 5022
rect 33506 4958 33518 5010
rect 33570 4958 33582 5010
rect 30382 4946 30434 4958
rect 36654 4946 36706 4958
rect 41918 5010 41970 5022
rect 41918 4946 41970 4958
rect 42478 5010 42530 5022
rect 42478 4946 42530 4958
rect 42702 5010 42754 5022
rect 42702 4946 42754 4958
rect 44718 5010 44770 5022
rect 44718 4946 44770 4958
rect 48190 5010 48242 5022
rect 48190 4946 48242 4958
rect 36542 4898 36594 4910
rect 18274 4846 18286 4898
rect 18338 4846 18350 4898
rect 21970 4846 21982 4898
rect 22034 4846 22046 4898
rect 31826 4846 31838 4898
rect 31890 4846 31902 4898
rect 36542 4834 36594 4846
rect 39790 4898 39842 4910
rect 39790 4834 39842 4846
rect 45726 4898 45778 4910
rect 45726 4834 45778 4846
rect 1344 4730 59024 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 59024 4730
rect 1344 4644 59024 4678
rect 23214 4562 23266 4574
rect 8418 4510 8430 4562
rect 8482 4510 8494 4562
rect 20738 4510 20750 4562
rect 20802 4510 20814 4562
rect 23214 4498 23266 4510
rect 23438 4562 23490 4574
rect 23438 4498 23490 4510
rect 24110 4562 24162 4574
rect 24110 4498 24162 4510
rect 24558 4562 24610 4574
rect 24558 4498 24610 4510
rect 25006 4562 25058 4574
rect 25006 4498 25058 4510
rect 25790 4562 25842 4574
rect 25790 4498 25842 4510
rect 30382 4562 30434 4574
rect 30382 4498 30434 4510
rect 32846 4562 32898 4574
rect 32846 4498 32898 4510
rect 40686 4562 40738 4574
rect 40686 4498 40738 4510
rect 40910 4562 40962 4574
rect 40910 4498 40962 4510
rect 43150 4562 43202 4574
rect 43150 4498 43202 4510
rect 45726 4562 45778 4574
rect 45726 4498 45778 4510
rect 45950 4562 46002 4574
rect 45950 4498 46002 4510
rect 21758 4450 21810 4462
rect 15026 4398 15038 4450
rect 15090 4398 15102 4450
rect 21758 4386 21810 4398
rect 23550 4450 23602 4462
rect 23550 4386 23602 4398
rect 26014 4450 26066 4462
rect 26014 4386 26066 4398
rect 26238 4450 26290 4462
rect 26238 4386 26290 4398
rect 28030 4450 28082 4462
rect 32398 4450 32450 4462
rect 28578 4398 28590 4450
rect 28642 4447 28654 4450
rect 28914 4447 28926 4450
rect 28642 4401 28926 4447
rect 28642 4398 28654 4401
rect 28914 4398 28926 4401
rect 28978 4398 28990 4450
rect 28030 4386 28082 4398
rect 32398 4386 32450 4398
rect 33630 4450 33682 4462
rect 33630 4386 33682 4398
rect 35198 4450 35250 4462
rect 35198 4386 35250 4398
rect 40574 4450 40626 4462
rect 40574 4386 40626 4398
rect 44046 4450 44098 4462
rect 44046 4386 44098 4398
rect 45614 4450 45666 4462
rect 45614 4386 45666 4398
rect 48638 4450 48690 4462
rect 48638 4386 48690 4398
rect 5630 4338 5682 4350
rect 9102 4338 9154 4350
rect 6066 4286 6078 4338
rect 6130 4286 6142 4338
rect 5630 4274 5682 4286
rect 9102 4274 9154 4286
rect 9774 4338 9826 4350
rect 17614 4338 17666 4350
rect 21310 4338 21362 4350
rect 25566 4338 25618 4350
rect 13010 4286 13022 4338
rect 13074 4286 13086 4338
rect 18162 4286 18174 4338
rect 18226 4286 18238 4338
rect 22194 4286 22206 4338
rect 22258 4286 22270 4338
rect 9774 4274 9826 4286
rect 17614 4274 17666 4286
rect 21310 4274 21362 4286
rect 25566 4274 25618 4286
rect 27246 4338 27298 4350
rect 27246 4274 27298 4286
rect 28366 4338 28418 4350
rect 28366 4274 28418 4286
rect 28478 4338 28530 4350
rect 36094 4338 36146 4350
rect 29250 4286 29262 4338
rect 29314 4286 29326 4338
rect 31490 4286 31502 4338
rect 31554 4286 31566 4338
rect 33842 4286 33854 4338
rect 33906 4286 33918 4338
rect 35522 4286 35534 4338
rect 35586 4286 35598 4338
rect 28478 4274 28530 4286
rect 36094 4274 36146 4286
rect 37214 4338 37266 4350
rect 37214 4274 37266 4286
rect 37438 4338 37490 4350
rect 48302 4338 48354 4350
rect 42018 4286 42030 4338
rect 42082 4286 42094 4338
rect 44482 4286 44494 4338
rect 44546 4286 44558 4338
rect 48066 4286 48078 4338
rect 48130 4286 48142 4338
rect 37438 4274 37490 4286
rect 48302 4274 48354 4286
rect 48526 4338 48578 4350
rect 48526 4274 48578 4286
rect 27470 4226 27522 4238
rect 10210 4174 10222 4226
rect 10274 4174 10286 4226
rect 22642 4174 22654 4226
rect 22706 4174 22718 4226
rect 26898 4174 26910 4226
rect 26962 4174 26974 4226
rect 27470 4162 27522 4174
rect 28142 4226 28194 4238
rect 34414 4226 34466 4238
rect 36206 4226 36258 4238
rect 29586 4174 29598 4226
rect 29650 4174 29662 4226
rect 31826 4174 31838 4226
rect 31890 4174 31902 4226
rect 35410 4174 35422 4226
rect 35474 4174 35486 4226
rect 28142 4162 28194 4174
rect 34414 4162 34466 4174
rect 36206 4162 36258 4174
rect 36990 4226 37042 4238
rect 36990 4162 37042 4174
rect 38782 4226 38834 4238
rect 42590 4226 42642 4238
rect 41906 4174 41918 4226
rect 41970 4174 41982 4226
rect 44818 4174 44830 4226
rect 44882 4174 44894 4226
rect 38782 4162 38834 4174
rect 42590 4162 42642 4174
rect 37886 4114 37938 4126
rect 37886 4050 37938 4062
rect 39006 4114 39058 4126
rect 39330 4062 39342 4114
rect 39394 4062 39406 4114
rect 39006 4050 39058 4062
rect 1344 3946 59024 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 59024 3946
rect 1344 3860 59024 3894
rect 25442 3726 25454 3778
rect 25506 3775 25518 3778
rect 25890 3775 25902 3778
rect 25506 3729 25902 3775
rect 25506 3726 25518 3729
rect 25890 3726 25902 3729
rect 25954 3726 25966 3778
rect 27682 3726 27694 3778
rect 27746 3775 27758 3778
rect 28466 3775 28478 3778
rect 27746 3729 28478 3775
rect 27746 3726 27758 3729
rect 28466 3726 28478 3729
rect 28530 3726 28542 3778
rect 6750 3666 6802 3678
rect 6750 3602 6802 3614
rect 7310 3666 7362 3678
rect 7310 3602 7362 3614
rect 7646 3666 7698 3678
rect 7646 3602 7698 3614
rect 9662 3666 9714 3678
rect 9662 3602 9714 3614
rect 10110 3666 10162 3678
rect 16382 3666 16434 3678
rect 15026 3614 15038 3666
rect 15090 3614 15102 3666
rect 10110 3602 10162 3614
rect 16382 3602 16434 3614
rect 16830 3666 16882 3678
rect 16830 3602 16882 3614
rect 18174 3666 18226 3678
rect 22094 3666 22146 3678
rect 19618 3614 19630 3666
rect 19682 3614 19694 3666
rect 18174 3602 18226 3614
rect 22094 3602 22146 3614
rect 22878 3666 22930 3678
rect 22878 3602 22930 3614
rect 23326 3666 23378 3678
rect 23326 3602 23378 3614
rect 23774 3666 23826 3678
rect 23774 3602 23826 3614
rect 24222 3666 24274 3678
rect 24222 3602 24274 3614
rect 24670 3666 24722 3678
rect 24670 3602 24722 3614
rect 25454 3666 25506 3678
rect 25454 3602 25506 3614
rect 25902 3666 25954 3678
rect 25902 3602 25954 3614
rect 26350 3666 26402 3678
rect 26350 3602 26402 3614
rect 26798 3666 26850 3678
rect 26798 3602 26850 3614
rect 27694 3666 27746 3678
rect 27694 3602 27746 3614
rect 28590 3666 28642 3678
rect 28590 3602 28642 3614
rect 29710 3666 29762 3678
rect 29710 3602 29762 3614
rect 32286 3666 32338 3678
rect 32286 3602 32338 3614
rect 33070 3666 33122 3678
rect 33070 3602 33122 3614
rect 34078 3666 34130 3678
rect 34078 3602 34130 3614
rect 34526 3666 34578 3678
rect 34526 3602 34578 3614
rect 35422 3666 35474 3678
rect 35422 3602 35474 3614
rect 35758 3666 35810 3678
rect 35758 3602 35810 3614
rect 36206 3666 36258 3678
rect 47518 3666 47570 3678
rect 39442 3614 39454 3666
rect 39506 3614 39518 3666
rect 36206 3602 36258 3614
rect 47518 3602 47570 3614
rect 5070 3554 5122 3566
rect 5070 3490 5122 3502
rect 5854 3554 5906 3566
rect 17726 3554 17778 3566
rect 21310 3554 21362 3566
rect 6290 3502 6302 3554
rect 6354 3502 6366 3554
rect 18610 3502 18622 3554
rect 18674 3502 18686 3554
rect 5854 3490 5906 3502
rect 17726 3490 17778 3502
rect 21310 3490 21362 3502
rect 21646 3554 21698 3566
rect 21646 3490 21698 3502
rect 28142 3554 28194 3566
rect 28142 3490 28194 3502
rect 29262 3554 29314 3566
rect 32174 3554 32226 3566
rect 31602 3502 31614 3554
rect 31666 3502 31678 3554
rect 29262 3490 29314 3502
rect 32174 3490 32226 3502
rect 37102 3554 37154 3566
rect 37102 3490 37154 3502
rect 37326 3554 37378 3566
rect 37326 3490 37378 3502
rect 41022 3554 41074 3566
rect 41022 3490 41074 3502
rect 42142 3554 42194 3566
rect 42142 3490 42194 3502
rect 12910 3442 12962 3454
rect 21534 3442 21586 3454
rect 13682 3390 13694 3442
rect 13746 3390 13758 3442
rect 12910 3378 12962 3390
rect 21534 3378 21586 3390
rect 27246 3442 27298 3454
rect 27246 3378 27298 3390
rect 30382 3442 30434 3454
rect 30382 3378 30434 3390
rect 34974 3442 35026 3454
rect 34974 3378 35026 3390
rect 37550 3442 37602 3454
rect 37550 3378 37602 3390
rect 38558 3442 38610 3454
rect 38558 3378 38610 3390
rect 40350 3442 40402 3454
rect 40350 3378 40402 3390
rect 41134 3442 41186 3454
rect 41134 3378 41186 3390
rect 41358 3442 41410 3454
rect 41358 3378 41410 3390
rect 41806 3442 41858 3454
rect 41806 3378 41858 3390
rect 41918 3442 41970 3454
rect 41918 3378 41970 3390
rect 48750 3442 48802 3454
rect 48750 3378 48802 3390
rect 55694 3442 55746 3454
rect 55694 3378 55746 3390
rect 56590 3442 56642 3454
rect 56590 3378 56642 3390
rect 37214 3330 37266 3342
rect 30706 3278 30718 3330
rect 30770 3278 30782 3330
rect 37214 3266 37266 3278
rect 39006 3330 39058 3342
rect 39006 3266 39058 3278
rect 48078 3330 48130 3342
rect 55346 3278 55358 3330
rect 55410 3278 55422 3330
rect 48078 3266 48130 3278
rect 1344 3162 59024 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 59024 3162
rect 1344 3076 59024 3110
rect 47394 2942 47406 2994
rect 47458 2991 47470 2994
rect 48066 2991 48078 2994
rect 47458 2945 48078 2991
rect 47458 2942 47470 2945
rect 48066 2942 48078 2945
rect 48130 2942 48142 2994
<< via1 >>
rect 4478 60342 4530 60394
rect 4582 60342 4634 60394
rect 4686 60342 4738 60394
rect 35198 60342 35250 60394
rect 35302 60342 35354 60394
rect 35406 60342 35458 60394
rect 21982 60174 22034 60226
rect 22542 60174 22594 60226
rect 22878 60174 22930 60226
rect 10446 60062 10498 60114
rect 31054 60062 31106 60114
rect 51102 60062 51154 60114
rect 4622 59950 4674 60002
rect 9774 59950 9826 60002
rect 11342 59950 11394 60002
rect 14590 59950 14642 60002
rect 23326 59950 23378 60002
rect 23550 59950 23602 60002
rect 30382 59950 30434 60002
rect 33966 59950 34018 60002
rect 50430 59950 50482 60002
rect 5070 59838 5122 59890
rect 6302 59838 6354 59890
rect 14702 59838 14754 59890
rect 15038 59838 15090 59890
rect 22766 59838 22818 59890
rect 22990 59838 23042 59890
rect 26910 59838 26962 59890
rect 33630 59838 33682 59890
rect 43710 59838 43762 59890
rect 3726 59726 3778 59778
rect 4174 59726 4226 59778
rect 5854 59726 5906 59778
rect 6750 59726 6802 59778
rect 7198 59726 7250 59778
rect 7646 59726 7698 59778
rect 8094 59726 8146 59778
rect 8542 59726 8594 59778
rect 8990 59726 9042 59778
rect 12350 59726 12402 59778
rect 12910 59726 12962 59778
rect 13582 59726 13634 59778
rect 14030 59726 14082 59778
rect 14926 59726 14978 59778
rect 15710 59726 15762 59778
rect 16158 59726 16210 59778
rect 16606 59726 16658 59778
rect 17614 59726 17666 59778
rect 18062 59726 18114 59778
rect 18734 59726 18786 59778
rect 19182 59726 19234 59778
rect 19742 59726 19794 59778
rect 20190 59726 20242 59778
rect 20638 59726 20690 59778
rect 21422 59726 21474 59778
rect 21870 59726 21922 59778
rect 22318 59726 22370 59778
rect 24222 59726 24274 59778
rect 24558 59726 24610 59778
rect 25230 59726 25282 59778
rect 27022 59726 27074 59778
rect 29822 59726 29874 59778
rect 33182 59726 33234 59778
rect 33742 59726 33794 59778
rect 34750 59726 34802 59778
rect 35534 59726 35586 59778
rect 42926 59726 42978 59778
rect 43822 59726 43874 59778
rect 44942 59726 44994 59778
rect 49870 59726 49922 59778
rect 19838 59558 19890 59610
rect 19942 59558 19994 59610
rect 20046 59558 20098 59610
rect 50558 59558 50610 59610
rect 50662 59558 50714 59610
rect 50766 59558 50818 59610
rect 4622 59390 4674 59442
rect 8990 59390 9042 59442
rect 10110 59390 10162 59442
rect 11006 59390 11058 59442
rect 12798 59390 12850 59442
rect 15934 59390 15986 59442
rect 17950 59390 18002 59442
rect 24894 59390 24946 59442
rect 25678 59390 25730 59442
rect 27918 59390 27970 59442
rect 34190 59390 34242 59442
rect 36990 59390 37042 59442
rect 5070 59278 5122 59330
rect 6414 59278 6466 59330
rect 8654 59278 8706 59330
rect 10670 59278 10722 59330
rect 19518 59278 19570 59330
rect 20078 59278 20130 59330
rect 29934 59278 29986 59330
rect 30158 59278 30210 59330
rect 30718 59278 30770 59330
rect 32622 59278 32674 59330
rect 34414 59278 34466 59330
rect 36430 59278 36482 59330
rect 38222 59278 38274 59330
rect 42030 59278 42082 59330
rect 42254 59278 42306 59330
rect 45502 59278 45554 59330
rect 14366 59166 14418 59218
rect 14590 59166 14642 59218
rect 14702 59166 14754 59218
rect 19070 59166 19122 59218
rect 20302 59166 20354 59218
rect 20526 59166 20578 59218
rect 21758 59166 21810 59218
rect 23886 59166 23938 59218
rect 24110 59166 24162 59218
rect 24334 59166 24386 59218
rect 26686 59166 26738 59218
rect 28030 59166 28082 59218
rect 28142 59166 28194 59218
rect 29822 59166 29874 59218
rect 30830 59166 30882 59218
rect 32510 59166 32562 59218
rect 32846 59166 32898 59218
rect 33966 59166 34018 59218
rect 35198 59166 35250 59218
rect 36318 59166 36370 59218
rect 36654 59166 36706 59218
rect 38110 59166 38162 59218
rect 38446 59166 38498 59218
rect 40574 59166 40626 59218
rect 41470 59166 41522 59218
rect 42702 59166 42754 59218
rect 43038 59166 43090 59218
rect 43486 59166 43538 59218
rect 43710 59166 43762 59218
rect 44270 59166 44322 59218
rect 44494 59166 44546 59218
rect 44942 59166 44994 59218
rect 45390 59166 45442 59218
rect 2718 59054 2770 59106
rect 3278 59054 3330 59106
rect 3614 59054 3666 59106
rect 4174 59054 4226 59106
rect 5406 59054 5458 59106
rect 5966 59054 6018 59106
rect 6862 59054 6914 59106
rect 7310 59054 7362 59106
rect 7758 59054 7810 59106
rect 8094 59054 8146 59106
rect 9662 59054 9714 59106
rect 11902 59054 11954 59106
rect 12350 59054 12402 59106
rect 13246 59054 13298 59106
rect 13694 59054 13746 59106
rect 16046 59054 16098 59106
rect 16606 59054 16658 59106
rect 17054 59054 17106 59106
rect 18622 59054 18674 59106
rect 20190 59054 20242 59106
rect 22094 59054 22146 59106
rect 26798 59054 26850 59106
rect 27246 59054 27298 59106
rect 28366 59054 28418 59106
rect 29374 59054 29426 59106
rect 31278 59054 31330 59106
rect 39454 59054 39506 59106
rect 42478 59054 42530 59106
rect 43262 59054 43314 59106
rect 44382 59054 44434 59106
rect 45950 59054 46002 59106
rect 15150 58942 15202 58994
rect 15710 58942 15762 58994
rect 22430 58942 22482 58994
rect 23550 58942 23602 58994
rect 28590 58942 28642 58994
rect 30718 58942 30770 58994
rect 34078 58942 34130 58994
rect 35086 58942 35138 58994
rect 35422 58942 35474 58994
rect 35534 58942 35586 58994
rect 38894 58942 38946 58994
rect 39230 58942 39282 58994
rect 40014 58942 40066 58994
rect 40350 58942 40402 58994
rect 4478 58774 4530 58826
rect 4582 58774 4634 58826
rect 4686 58774 4738 58826
rect 35198 58774 35250 58826
rect 35302 58774 35354 58826
rect 35406 58774 35458 58826
rect 11230 58606 11282 58658
rect 11902 58606 11954 58658
rect 30158 58606 30210 58658
rect 37662 58606 37714 58658
rect 40574 58606 40626 58658
rect 44382 58606 44434 58658
rect 12126 58494 12178 58546
rect 16606 58494 16658 58546
rect 18174 58494 18226 58546
rect 19070 58494 19122 58546
rect 22094 58494 22146 58546
rect 24558 58494 24610 58546
rect 27358 58494 27410 58546
rect 28702 58494 28754 58546
rect 29934 58494 29986 58546
rect 32958 58494 33010 58546
rect 36430 58494 36482 58546
rect 36766 58494 36818 58546
rect 41246 58494 41298 58546
rect 42814 58494 42866 58546
rect 46398 58494 46450 58546
rect 47182 58494 47234 58546
rect 50654 58494 50706 58546
rect 51214 58494 51266 58546
rect 13022 58382 13074 58434
rect 13806 58382 13858 58434
rect 14030 58382 14082 58434
rect 15150 58382 15202 58434
rect 16270 58382 16322 58434
rect 17502 58382 17554 58434
rect 18062 58382 18114 58434
rect 19182 58382 19234 58434
rect 22318 58382 22370 58434
rect 23774 58382 23826 58434
rect 24782 58382 24834 58434
rect 25454 58382 25506 58434
rect 25902 58382 25954 58434
rect 26910 58382 26962 58434
rect 30494 58382 30546 58434
rect 31502 58382 31554 58434
rect 32062 58382 32114 58434
rect 33182 58382 33234 58434
rect 33518 58382 33570 58434
rect 34414 58382 34466 58434
rect 34750 58382 34802 58434
rect 34974 58382 35026 58434
rect 36094 58382 36146 58434
rect 37550 58382 37602 58434
rect 38670 58382 38722 58434
rect 39118 58382 39170 58434
rect 39454 58382 39506 58434
rect 40014 58382 40066 58434
rect 40574 58382 40626 58434
rect 42030 58382 42082 58434
rect 42366 58382 42418 58434
rect 43486 58382 43538 58434
rect 44158 58382 44210 58434
rect 44606 58382 44658 58434
rect 46622 58382 46674 58434
rect 47518 58382 47570 58434
rect 50094 58382 50146 58434
rect 50430 58382 50482 58434
rect 7310 58270 7362 58322
rect 9102 58270 9154 58322
rect 9886 58270 9938 58322
rect 12686 58270 12738 58322
rect 14702 58270 14754 58322
rect 15486 58270 15538 58322
rect 19854 58270 19906 58322
rect 22878 58270 22930 58322
rect 23438 58270 23490 58322
rect 24446 58270 24498 58322
rect 26350 58270 26402 58322
rect 27134 58270 27186 58322
rect 27470 58270 27522 58322
rect 28814 58270 28866 58322
rect 32286 58270 32338 58322
rect 37662 58270 37714 58322
rect 40238 58270 40290 58322
rect 43150 58270 43202 58322
rect 51550 58270 51602 58322
rect 1934 58158 1986 58210
rect 2494 58158 2546 58210
rect 2942 58158 2994 58210
rect 3390 58158 3442 58210
rect 3950 58158 4002 58210
rect 4510 58158 4562 58210
rect 4958 58158 5010 58210
rect 5966 58158 6018 58210
rect 6302 58158 6354 58210
rect 6750 58158 6802 58210
rect 7758 58158 7810 58210
rect 8206 58158 8258 58210
rect 8654 58158 8706 58210
rect 9438 58158 9490 58210
rect 10446 58158 10498 58210
rect 10782 58158 10834 58210
rect 11342 58158 11394 58210
rect 11678 58158 11730 58210
rect 12798 58158 12850 58210
rect 15374 58158 15426 58210
rect 16494 58158 16546 58210
rect 20526 58158 20578 58210
rect 20974 58158 21026 58210
rect 23550 58158 23602 58210
rect 28590 58158 28642 58210
rect 31166 58158 31218 58210
rect 34862 58158 34914 58210
rect 38782 58158 38834 58210
rect 38894 58158 38946 58210
rect 40126 58158 40178 58210
rect 44270 58158 44322 58210
rect 45390 58158 45442 58210
rect 46062 58158 46114 58210
rect 47294 58158 47346 58210
rect 51326 58158 51378 58210
rect 19838 57990 19890 58042
rect 19942 57990 19994 58042
rect 20046 57990 20098 58042
rect 50558 57990 50610 58042
rect 50662 57990 50714 58042
rect 50766 57990 50818 58042
rect 3166 57822 3218 57874
rect 4062 57822 4114 57874
rect 8990 57822 9042 57874
rect 16382 57822 16434 57874
rect 19294 57822 19346 57874
rect 20414 57822 20466 57874
rect 27918 57822 27970 57874
rect 28142 57822 28194 57874
rect 29486 57822 29538 57874
rect 29822 57822 29874 57874
rect 33742 57822 33794 57874
rect 33966 57822 34018 57874
rect 35646 57822 35698 57874
rect 36430 57822 36482 57874
rect 38110 57822 38162 57874
rect 39678 57822 39730 57874
rect 40462 57822 40514 57874
rect 42142 57822 42194 57874
rect 43262 57822 43314 57874
rect 43486 57822 43538 57874
rect 44158 57822 44210 57874
rect 44494 57822 44546 57874
rect 44606 57822 44658 57874
rect 46734 57822 46786 57874
rect 14366 57710 14418 57762
rect 23102 57710 23154 57762
rect 27806 57710 27858 57762
rect 28590 57710 28642 57762
rect 29710 57710 29762 57762
rect 31278 57710 31330 57762
rect 33630 57710 33682 57762
rect 34526 57710 34578 57762
rect 36318 57710 36370 57762
rect 36990 57710 37042 57762
rect 40350 57710 40402 57762
rect 51214 57710 51266 57762
rect 9998 57598 10050 57650
rect 10446 57598 10498 57650
rect 13806 57598 13858 57650
rect 14254 57598 14306 57650
rect 18958 57598 19010 57650
rect 19854 57598 19906 57650
rect 20078 57598 20130 57650
rect 21982 57598 22034 57650
rect 23438 57598 23490 57650
rect 23662 57598 23714 57650
rect 28702 57598 28754 57650
rect 29150 57598 29202 57650
rect 30606 57598 30658 57650
rect 31166 57598 31218 57650
rect 32062 57598 32114 57650
rect 32398 57598 32450 57650
rect 32734 57598 32786 57650
rect 34750 57598 34802 57650
rect 35086 57598 35138 57650
rect 38222 57598 38274 57650
rect 38446 57598 38498 57650
rect 38670 57598 38722 57650
rect 39230 57598 39282 57650
rect 39454 57598 39506 57650
rect 39790 57598 39842 57650
rect 41806 57598 41858 57650
rect 42814 57598 42866 57650
rect 44382 57598 44434 57650
rect 46286 57598 46338 57650
rect 46510 57598 46562 57650
rect 46958 57598 47010 57650
rect 47518 57598 47570 57650
rect 47742 57598 47794 57650
rect 48078 57598 48130 57650
rect 50206 57598 50258 57650
rect 51886 57598 51938 57650
rect 52110 57598 52162 57650
rect 52334 57598 52386 57650
rect 2158 57486 2210 57538
rect 2830 57486 2882 57538
rect 3726 57486 3778 57538
rect 4622 57486 4674 57538
rect 5070 57486 5122 57538
rect 5518 57486 5570 57538
rect 5854 57486 5906 57538
rect 6414 57486 6466 57538
rect 6862 57486 6914 57538
rect 7198 57486 7250 57538
rect 7646 57486 7698 57538
rect 8094 57486 8146 57538
rect 8542 57486 8594 57538
rect 10894 57486 10946 57538
rect 11230 57486 11282 57538
rect 12014 57486 12066 57538
rect 12350 57486 12402 57538
rect 12798 57486 12850 57538
rect 14926 57486 14978 57538
rect 15374 57486 15426 57538
rect 16270 57486 16322 57538
rect 17614 57486 17666 57538
rect 18174 57486 18226 57538
rect 18734 57486 18786 57538
rect 20974 57486 21026 57538
rect 21422 57486 21474 57538
rect 23214 57486 23266 57538
rect 24110 57486 24162 57538
rect 24558 57486 24610 57538
rect 25566 57486 25618 57538
rect 26014 57486 26066 57538
rect 32510 57486 32562 57538
rect 34974 57486 35026 57538
rect 37438 57486 37490 57538
rect 38334 57486 38386 57538
rect 41582 57486 41634 57538
rect 43374 57486 43426 57538
rect 45054 57486 45106 57538
rect 45502 57486 45554 57538
rect 47854 57486 47906 57538
rect 50318 57486 50370 57538
rect 50542 57486 50594 57538
rect 51998 57486 52050 57538
rect 53118 57486 53170 57538
rect 53566 57486 53618 57538
rect 54014 57486 54066 57538
rect 6750 57374 6802 57426
rect 7870 57374 7922 57426
rect 8094 57374 8146 57426
rect 8542 57374 8594 57426
rect 16606 57374 16658 57426
rect 22206 57374 22258 57426
rect 22542 57374 22594 57426
rect 36542 57374 36594 57426
rect 51326 57374 51378 57426
rect 53118 57374 53170 57426
rect 53902 57374 53954 57426
rect 4478 57206 4530 57258
rect 4582 57206 4634 57258
rect 4686 57206 4738 57258
rect 35198 57206 35250 57258
rect 35302 57206 35354 57258
rect 35406 57206 35458 57258
rect 6974 57038 7026 57090
rect 11118 57038 11170 57090
rect 17726 57038 17778 57090
rect 22766 57038 22818 57090
rect 23550 57038 23602 57090
rect 23998 57038 24050 57090
rect 34638 57038 34690 57090
rect 35646 57038 35698 57090
rect 35870 57038 35922 57090
rect 43486 57038 43538 57090
rect 43822 57038 43874 57090
rect 47070 57038 47122 57090
rect 1934 56926 1986 56978
rect 2382 56926 2434 56978
rect 6974 56926 7026 56978
rect 8206 56926 8258 56978
rect 8766 56926 8818 56978
rect 13582 56926 13634 56978
rect 16718 56926 16770 56978
rect 19070 56926 19122 56978
rect 20190 56926 20242 56978
rect 25790 56926 25842 56978
rect 26126 56926 26178 56978
rect 26574 56926 26626 56978
rect 28702 56926 28754 56978
rect 29598 56926 29650 56978
rect 34750 56926 34802 56978
rect 42590 56926 42642 56978
rect 43262 56926 43314 56978
rect 46286 56926 46338 56978
rect 51998 56926 52050 56978
rect 53790 56926 53842 56978
rect 11118 56814 11170 56866
rect 12350 56814 12402 56866
rect 14142 56814 14194 56866
rect 16046 56814 16098 56866
rect 16494 56814 16546 56866
rect 17502 56814 17554 56866
rect 17838 56814 17890 56866
rect 22206 56814 22258 56866
rect 23326 56814 23378 56866
rect 23774 56814 23826 56866
rect 24558 56814 24610 56866
rect 25006 56814 25058 56866
rect 25118 56814 25170 56866
rect 28814 56814 28866 56866
rect 30046 56814 30098 56866
rect 30494 56814 30546 56866
rect 31054 56814 31106 56866
rect 31726 56814 31778 56866
rect 36094 56814 36146 56866
rect 36318 56814 36370 56866
rect 36542 56814 36594 56866
rect 38670 56814 38722 56866
rect 38782 56814 38834 56866
rect 39342 56814 39394 56866
rect 39454 56814 39506 56866
rect 40014 56814 40066 56866
rect 40686 56814 40738 56866
rect 46398 56814 46450 56866
rect 48190 56814 48242 56866
rect 48302 56814 48354 56866
rect 49982 56814 50034 56866
rect 50094 56814 50146 56866
rect 50654 56814 50706 56866
rect 51214 56814 51266 56866
rect 51662 56814 51714 56866
rect 52222 56814 52274 56866
rect 53342 56814 53394 56866
rect 54126 56814 54178 56866
rect 54686 56814 54738 56866
rect 17278 56702 17330 56754
rect 18958 56702 19010 56754
rect 19182 56702 19234 56754
rect 22094 56702 22146 56754
rect 22318 56702 22370 56754
rect 24110 56702 24162 56754
rect 28590 56702 28642 56754
rect 31502 56702 31554 56754
rect 32174 56702 32226 56754
rect 36430 56702 36482 56754
rect 38558 56702 38610 56754
rect 48414 56702 48466 56754
rect 52334 56702 52386 56754
rect 2830 56590 2882 56642
rect 3502 56590 3554 56642
rect 3950 56590 4002 56642
rect 4286 56590 4338 56642
rect 4846 56590 4898 56642
rect 6078 56590 6130 56642
rect 6414 56590 6466 56642
rect 7422 56590 7474 56642
rect 7870 56590 7922 56642
rect 9214 56590 9266 56642
rect 9774 56590 9826 56642
rect 10222 56590 10274 56642
rect 10670 56590 10722 56642
rect 11566 56590 11618 56642
rect 11902 56590 11954 56642
rect 12686 56590 12738 56642
rect 12910 56590 12962 56642
rect 13022 56590 13074 56642
rect 14590 56590 14642 56642
rect 15038 56590 15090 56642
rect 18062 56590 18114 56642
rect 19854 56590 19906 56642
rect 20750 56590 20802 56642
rect 25230 56590 25282 56642
rect 27022 56590 27074 56642
rect 31390 56590 31442 56642
rect 32622 56590 32674 56642
rect 37662 56590 37714 56642
rect 39006 56590 39058 56642
rect 40126 56590 40178 56642
rect 40238 56590 40290 56642
rect 41022 56590 41074 56642
rect 47742 56590 47794 56642
rect 50206 56590 50258 56642
rect 55246 56590 55298 56642
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 2718 56254 2770 56306
rect 5406 56254 5458 56306
rect 5854 56254 5906 56306
rect 6862 56254 6914 56306
rect 7646 56254 7698 56306
rect 8542 56254 8594 56306
rect 11118 56254 11170 56306
rect 14366 56254 14418 56306
rect 15262 56254 15314 56306
rect 16494 56254 16546 56306
rect 16942 56254 16994 56306
rect 18622 56254 18674 56306
rect 20974 56254 21026 56306
rect 22542 56254 22594 56306
rect 23662 56254 23714 56306
rect 26462 56254 26514 56306
rect 27806 56254 27858 56306
rect 30158 56254 30210 56306
rect 30718 56254 30770 56306
rect 35534 56254 35586 56306
rect 38222 56254 38274 56306
rect 40014 56254 40066 56306
rect 42814 56254 42866 56306
rect 43934 56254 43986 56306
rect 44158 56254 44210 56306
rect 51102 56254 51154 56306
rect 54014 56254 54066 56306
rect 9998 56142 10050 56194
rect 12798 56142 12850 56194
rect 13470 56142 13522 56194
rect 13694 56142 13746 56194
rect 19294 56142 19346 56194
rect 46510 56142 46562 56194
rect 51214 56142 51266 56194
rect 52334 56142 52386 56194
rect 1934 56030 1986 56082
rect 8094 56030 8146 56082
rect 11006 56030 11058 56082
rect 11342 56030 11394 56082
rect 12126 56030 12178 56082
rect 14254 56030 14306 56082
rect 21422 56030 21474 56082
rect 21982 56030 22034 56082
rect 22318 56030 22370 56082
rect 22430 56030 22482 56082
rect 22654 56030 22706 56082
rect 23886 56030 23938 56082
rect 24334 56030 24386 56082
rect 26238 56030 26290 56082
rect 26574 56030 26626 56082
rect 26798 56030 26850 56082
rect 39118 56030 39170 56082
rect 39342 56030 39394 56082
rect 44606 56030 44658 56082
rect 46734 56030 46786 56082
rect 50206 56030 50258 56082
rect 51774 56030 51826 56082
rect 51998 56030 52050 56082
rect 52222 56030 52274 56082
rect 2382 55918 2434 55970
rect 3166 55918 3218 55970
rect 3614 55918 3666 55970
rect 4062 55918 4114 55970
rect 4622 55918 4674 55970
rect 5070 55918 5122 55970
rect 6302 55918 6354 55970
rect 7310 55918 7362 55970
rect 8990 55918 9042 55970
rect 10446 55918 10498 55970
rect 11902 55918 11954 55970
rect 14030 55918 14082 55970
rect 14926 55918 14978 55970
rect 16046 55918 16098 55970
rect 17614 55918 17666 55970
rect 18174 55918 18226 55970
rect 19182 55918 19234 55970
rect 20190 55918 20242 55970
rect 23774 55918 23826 55970
rect 24670 55918 24722 55970
rect 25566 55918 25618 55970
rect 27358 55918 27410 55970
rect 28254 55918 28306 55970
rect 31278 55918 31330 55970
rect 31838 55918 31890 55970
rect 35086 55918 35138 55970
rect 38558 55918 38610 55970
rect 40350 55918 40402 55970
rect 43374 55918 43426 55970
rect 44046 55918 44098 55970
rect 44382 55918 44434 55970
rect 44830 55918 44882 55970
rect 48302 55918 48354 55970
rect 49534 55918 49586 55970
rect 50318 55918 50370 55970
rect 52894 55918 52946 55970
rect 53902 55918 53954 55970
rect 54462 55918 54514 55970
rect 5966 55806 6018 55858
rect 7870 55806 7922 55858
rect 19518 55806 19570 55858
rect 20078 55806 20130 55858
rect 31390 55806 31442 55858
rect 39566 55806 39618 55858
rect 47070 55806 47122 55858
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 6750 55470 6802 55522
rect 6974 55470 7026 55522
rect 7646 55470 7698 55522
rect 8206 55470 8258 55522
rect 8878 55470 8930 55522
rect 10670 55470 10722 55522
rect 11678 55470 11730 55522
rect 14142 55470 14194 55522
rect 14478 55470 14530 55522
rect 14926 55470 14978 55522
rect 22990 55470 23042 55522
rect 37550 55470 37602 55522
rect 38782 55470 38834 55522
rect 43262 55470 43314 55522
rect 3614 55358 3666 55410
rect 5854 55358 5906 55410
rect 6750 55358 6802 55410
rect 7646 55358 7698 55410
rect 8542 55358 8594 55410
rect 12126 55358 12178 55410
rect 12910 55358 12962 55410
rect 13806 55358 13858 55410
rect 15150 55358 15202 55410
rect 16606 55358 16658 55410
rect 18958 55358 19010 55410
rect 20638 55358 20690 55410
rect 23326 55358 23378 55410
rect 25566 55358 25618 55410
rect 28030 55358 28082 55410
rect 32286 55358 32338 55410
rect 35982 55358 36034 55410
rect 41358 55358 41410 55410
rect 42590 55358 42642 55410
rect 46510 55358 46562 55410
rect 47854 55358 47906 55410
rect 53678 55358 53730 55410
rect 12462 55246 12514 55298
rect 18734 55246 18786 55298
rect 19742 55246 19794 55298
rect 19966 55246 20018 55298
rect 24670 55246 24722 55298
rect 26014 55246 26066 55298
rect 26462 55246 26514 55298
rect 27134 55246 27186 55298
rect 27582 55246 27634 55298
rect 32174 55246 32226 55298
rect 33406 55246 33458 55298
rect 33742 55246 33794 55298
rect 34302 55246 34354 55298
rect 35646 55246 35698 55298
rect 37886 55246 37938 55298
rect 38110 55246 38162 55298
rect 39454 55246 39506 55298
rect 39678 55246 39730 55298
rect 40462 55246 40514 55298
rect 40686 55246 40738 55298
rect 42478 55246 42530 55298
rect 46958 55246 47010 55298
rect 47294 55246 47346 55298
rect 47518 55246 47570 55298
rect 47742 55246 47794 55298
rect 1822 55134 1874 55186
rect 9998 55134 10050 55186
rect 16718 55134 16770 55186
rect 16942 55134 16994 55186
rect 19070 55134 19122 55186
rect 28478 55134 28530 55186
rect 29934 55134 29986 55186
rect 32510 55134 32562 55186
rect 32734 55134 32786 55186
rect 36318 55134 36370 55186
rect 38670 55134 38722 55186
rect 39790 55134 39842 55186
rect 47966 55134 48018 55186
rect 48414 55134 48466 55186
rect 53790 55134 53842 55186
rect 54014 55134 54066 55186
rect 2158 55022 2210 55074
rect 2606 55022 2658 55074
rect 3054 55022 3106 55074
rect 3950 55022 4002 55074
rect 4398 55022 4450 55074
rect 4846 55022 4898 55074
rect 6414 55022 6466 55074
rect 7198 55022 7250 55074
rect 8094 55022 8146 55074
rect 8990 55022 9042 55074
rect 9550 55022 9602 55074
rect 10446 55022 10498 55074
rect 10894 55022 10946 55074
rect 11342 55022 11394 55074
rect 13918 55022 13970 55074
rect 14590 55022 14642 55074
rect 15710 55022 15762 55074
rect 16158 55022 16210 55074
rect 17390 55022 17442 55074
rect 17838 55022 17890 55074
rect 21758 55022 21810 55074
rect 22206 55022 22258 55074
rect 23214 55022 23266 55074
rect 23774 55022 23826 55074
rect 24222 55022 24274 55074
rect 29822 55022 29874 55074
rect 38782 55022 38834 55074
rect 49086 55022 49138 55074
rect 54462 55022 54514 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 2270 54686 2322 54738
rect 2718 54686 2770 54738
rect 7646 54686 7698 54738
rect 8542 54686 8594 54738
rect 8990 54686 9042 54738
rect 10558 54686 10610 54738
rect 11454 54686 11506 54738
rect 12014 54686 12066 54738
rect 13022 54686 13074 54738
rect 16830 54686 16882 54738
rect 21870 54686 21922 54738
rect 22766 54686 22818 54738
rect 23998 54686 24050 54738
rect 24446 54686 24498 54738
rect 26686 54686 26738 54738
rect 35422 54686 35474 54738
rect 35534 54686 35586 54738
rect 41806 54686 41858 54738
rect 46398 54686 46450 54738
rect 47406 54686 47458 54738
rect 48302 54686 48354 54738
rect 48414 54686 48466 54738
rect 51438 54686 51490 54738
rect 52222 54686 52274 54738
rect 53454 54686 53506 54738
rect 1822 54574 1874 54626
rect 13246 54574 13298 54626
rect 14030 54574 14082 54626
rect 14142 54574 14194 54626
rect 15038 54574 15090 54626
rect 16606 54574 16658 54626
rect 19070 54574 19122 54626
rect 27134 54574 27186 54626
rect 32846 54574 32898 54626
rect 39454 54574 39506 54626
rect 41918 54574 41970 54626
rect 42926 54574 42978 54626
rect 46174 54574 46226 54626
rect 47294 54574 47346 54626
rect 48526 54574 48578 54626
rect 50542 54574 50594 54626
rect 52446 54574 52498 54626
rect 54350 54574 54402 54626
rect 4398 54462 4450 54514
rect 4958 54462 5010 54514
rect 13806 54462 13858 54514
rect 15598 54462 15650 54514
rect 19518 54462 19570 54514
rect 19966 54462 20018 54514
rect 27246 54462 27298 54514
rect 27470 54462 27522 54514
rect 28142 54462 28194 54514
rect 28590 54462 28642 54514
rect 29038 54462 29090 54514
rect 30158 54462 30210 54514
rect 32398 54462 32450 54514
rect 35758 54462 35810 54514
rect 35982 54462 36034 54514
rect 36542 54462 36594 54514
rect 41582 54462 41634 54514
rect 46062 54462 46114 54514
rect 48078 54462 48130 54514
rect 48750 54462 48802 54514
rect 49870 54462 49922 54514
rect 51214 54462 51266 54514
rect 51438 54462 51490 54514
rect 51774 54462 51826 54514
rect 52558 54462 52610 54514
rect 53006 54462 53058 54514
rect 53678 54462 53730 54514
rect 54238 54462 54290 54514
rect 3166 54350 3218 54402
rect 3502 54350 3554 54402
rect 3950 54350 4002 54402
rect 5294 54350 5346 54402
rect 5742 54350 5794 54402
rect 6414 54350 6466 54402
rect 6750 54350 6802 54402
rect 7310 54350 7362 54402
rect 8206 54350 8258 54402
rect 9662 54350 9714 54402
rect 10222 54350 10274 54402
rect 11118 54350 11170 54402
rect 12350 54350 12402 54402
rect 12910 54350 12962 54402
rect 17614 54350 17666 54402
rect 18062 54350 18114 54402
rect 18622 54350 18674 54402
rect 20638 54350 20690 54402
rect 21086 54350 21138 54402
rect 22318 54350 22370 54402
rect 23326 54350 23378 54402
rect 25006 54350 25058 54402
rect 25678 54350 25730 54402
rect 26126 54350 26178 54402
rect 29934 54350 29986 54402
rect 30830 54350 30882 54402
rect 32510 54350 32562 54402
rect 33742 54350 33794 54402
rect 35646 54350 35698 54402
rect 36430 54350 36482 54402
rect 39342 54350 39394 54402
rect 43038 54350 43090 54402
rect 50094 54350 50146 54402
rect 53566 54350 53618 54402
rect 2158 54238 2210 54290
rect 2494 54238 2546 54290
rect 10894 54238 10946 54290
rect 12350 54238 12402 54290
rect 33630 54238 33682 54290
rect 36206 54238 36258 54290
rect 39678 54238 39730 54290
rect 43150 54238 43202 54290
rect 47518 54238 47570 54290
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 5854 53902 5906 53954
rect 6302 53902 6354 53954
rect 14030 53902 14082 53954
rect 15822 53902 15874 53954
rect 15934 53902 15986 53954
rect 16382 53902 16434 53954
rect 16606 53902 16658 53954
rect 19070 53902 19122 53954
rect 28702 53902 28754 53954
rect 32510 53902 32562 53954
rect 40350 53902 40402 53954
rect 3278 53790 3330 53842
rect 3726 53790 3778 53842
rect 7086 53790 7138 53842
rect 8766 53790 8818 53842
rect 9662 53790 9714 53842
rect 11902 53790 11954 53842
rect 12238 53790 12290 53842
rect 13694 53790 13746 53842
rect 18510 53790 18562 53842
rect 20414 53790 20466 53842
rect 20526 53790 20578 53842
rect 29710 53790 29762 53842
rect 32734 53790 32786 53842
rect 35982 53790 36034 53842
rect 39678 53790 39730 53842
rect 42702 53790 42754 53842
rect 44718 53790 44770 53842
rect 45950 53790 46002 53842
rect 48190 53790 48242 53842
rect 52222 53790 52274 53842
rect 2382 53678 2434 53730
rect 4174 53678 4226 53730
rect 4958 53678 5010 53730
rect 6526 53678 6578 53730
rect 7534 53678 7586 53730
rect 9214 53678 9266 53730
rect 10110 53678 10162 53730
rect 12574 53678 12626 53730
rect 14590 53678 14642 53730
rect 14926 53678 14978 53730
rect 15934 53678 15986 53730
rect 19406 53678 19458 53730
rect 19630 53678 19682 53730
rect 19742 53678 19794 53730
rect 22430 53678 22482 53730
rect 23662 53678 23714 53730
rect 23998 53678 24050 53730
rect 24222 53678 24274 53730
rect 26238 53678 26290 53730
rect 27246 53678 27298 53730
rect 27582 53678 27634 53730
rect 29598 53678 29650 53730
rect 29822 53678 29874 53730
rect 30158 53678 30210 53730
rect 35422 53678 35474 53730
rect 35758 53678 35810 53730
rect 36430 53678 36482 53730
rect 39566 53678 39618 53730
rect 41694 53678 41746 53730
rect 44046 53678 44098 53730
rect 46174 53678 46226 53730
rect 46846 53678 46898 53730
rect 48526 53678 48578 53730
rect 49422 53678 49474 53730
rect 51326 53678 51378 53730
rect 51774 53678 51826 53730
rect 53454 53678 53506 53730
rect 53566 53678 53618 53730
rect 53902 53678 53954 53730
rect 2046 53566 2098 53618
rect 14702 53566 14754 53618
rect 22990 53566 23042 53618
rect 27358 53566 27410 53618
rect 28814 53566 28866 53618
rect 32734 53566 32786 53618
rect 33406 53566 33458 53618
rect 33518 53566 33570 53618
rect 35086 53566 35138 53618
rect 36206 53566 36258 53618
rect 43038 53566 43090 53618
rect 48190 53566 48242 53618
rect 49086 53566 49138 53618
rect 2830 53454 2882 53506
rect 5630 53454 5682 53506
rect 6078 53454 6130 53506
rect 7982 53454 8034 53506
rect 8318 53454 8370 53506
rect 10894 53454 10946 53506
rect 11342 53454 11394 53506
rect 13806 53454 13858 53506
rect 15374 53454 15426 53506
rect 17166 53454 17218 53506
rect 17614 53454 17666 53506
rect 18062 53454 18114 53506
rect 19518 53454 19570 53506
rect 20638 53454 20690 53506
rect 21982 53454 22034 53506
rect 22654 53454 22706 53506
rect 22766 53454 22818 53506
rect 22878 53454 22930 53506
rect 23886 53454 23938 53506
rect 24110 53454 24162 53506
rect 24894 53454 24946 53506
rect 25342 53454 25394 53506
rect 25678 53454 25730 53506
rect 26798 53454 26850 53506
rect 28030 53454 28082 53506
rect 35198 53454 35250 53506
rect 41806 53454 41858 53506
rect 42030 53454 42082 53506
rect 47294 53454 47346 53506
rect 47966 53454 48018 53506
rect 49198 53454 49250 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 3054 53118 3106 53170
rect 4510 53118 4562 53170
rect 5070 53118 5122 53170
rect 5854 53118 5906 53170
rect 6302 53118 6354 53170
rect 6750 53118 6802 53170
rect 7198 53118 7250 53170
rect 8990 53118 9042 53170
rect 9886 53118 9938 53170
rect 10334 53118 10386 53170
rect 11790 53118 11842 53170
rect 12686 53118 12738 53170
rect 20526 53118 20578 53170
rect 21534 53118 21586 53170
rect 22430 53118 22482 53170
rect 26910 53118 26962 53170
rect 33966 53118 34018 53170
rect 39566 53118 39618 53170
rect 42814 53118 42866 53170
rect 5406 53006 5458 53058
rect 18286 53006 18338 53058
rect 19854 53006 19906 53058
rect 20414 53006 20466 53058
rect 20638 53006 20690 53058
rect 21982 53006 22034 53058
rect 23774 53006 23826 53058
rect 24670 53006 24722 53058
rect 24894 53006 24946 53058
rect 29038 53006 29090 53058
rect 30270 53006 30322 53058
rect 33742 53006 33794 53058
rect 38334 53006 38386 53058
rect 43262 53006 43314 53058
rect 50654 53006 50706 53058
rect 2270 52894 2322 52946
rect 14814 52894 14866 52946
rect 22206 52894 22258 52946
rect 22542 52894 22594 52946
rect 23326 52894 23378 52946
rect 23550 52894 23602 52946
rect 23998 52894 24050 52946
rect 26462 52894 26514 52946
rect 26798 52894 26850 52946
rect 27022 52894 27074 52946
rect 29710 52894 29762 52946
rect 30046 52894 30098 52946
rect 33630 52894 33682 52946
rect 36542 52894 36594 52946
rect 37550 52894 37602 52946
rect 39342 52894 39394 52946
rect 39566 52894 39618 52946
rect 39790 52894 39842 52946
rect 42590 52894 42642 52946
rect 43038 52894 43090 52946
rect 49870 52894 49922 52946
rect 53230 52894 53282 52946
rect 53566 52894 53618 52946
rect 1822 52782 1874 52834
rect 2718 52782 2770 52834
rect 3502 52782 3554 52834
rect 4174 52782 4226 52834
rect 7646 52782 7698 52834
rect 8094 52782 8146 52834
rect 8542 52782 8594 52834
rect 10894 52782 10946 52834
rect 11342 52782 11394 52834
rect 12238 52782 12290 52834
rect 13134 52782 13186 52834
rect 13918 52782 13970 52834
rect 14366 52782 14418 52834
rect 15374 52782 15426 52834
rect 16046 52782 16098 52834
rect 16494 52782 16546 52834
rect 16942 52782 16994 52834
rect 18958 52782 19010 52834
rect 19518 52782 19570 52834
rect 22430 52782 22482 52834
rect 23886 52782 23938 52834
rect 24558 52782 24610 52834
rect 25678 52782 25730 52834
rect 27470 52782 27522 52834
rect 27918 52782 27970 52834
rect 28366 52782 28418 52834
rect 30158 52782 30210 52834
rect 36654 52782 36706 52834
rect 40350 52782 40402 52834
rect 47742 52782 47794 52834
rect 50094 52782 50146 52834
rect 53118 52782 53170 52834
rect 5966 52670 6018 52722
rect 8430 52670 8482 52722
rect 11790 52670 11842 52722
rect 12126 52670 12178 52722
rect 13918 52670 13970 52722
rect 14478 52670 14530 52722
rect 18062 52670 18114 52722
rect 18398 52670 18450 52722
rect 18734 52670 18786 52722
rect 19966 52670 20018 52722
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 2494 52334 2546 52386
rect 2718 52334 2770 52386
rect 25006 52334 25058 52386
rect 40574 52334 40626 52386
rect 1822 52222 1874 52274
rect 2270 52222 2322 52274
rect 3054 52222 3106 52274
rect 4286 52222 4338 52274
rect 6078 52222 6130 52274
rect 6526 52222 6578 52274
rect 6974 52222 7026 52274
rect 8094 52222 8146 52274
rect 8542 52222 8594 52274
rect 9438 52222 9490 52274
rect 13806 52222 13858 52274
rect 14254 52222 14306 52274
rect 17166 52222 17218 52274
rect 18398 52222 18450 52274
rect 19406 52222 19458 52274
rect 19966 52222 20018 52274
rect 20526 52222 20578 52274
rect 22094 52222 22146 52274
rect 22766 52222 22818 52274
rect 24334 52222 24386 52274
rect 26350 52222 26402 52274
rect 30606 52222 30658 52274
rect 33070 52222 33122 52274
rect 35086 52222 35138 52274
rect 39902 52222 39954 52274
rect 46062 52222 46114 52274
rect 53454 52222 53506 52274
rect 4846 52110 4898 52162
rect 9102 52110 9154 52162
rect 10558 52110 10610 52162
rect 11118 52110 11170 52162
rect 11678 52110 11730 52162
rect 12462 52110 12514 52162
rect 13022 52110 13074 52162
rect 15150 52110 15202 52162
rect 15710 52110 15762 52162
rect 16046 52110 16098 52162
rect 18286 52110 18338 52162
rect 20862 52110 20914 52162
rect 21534 52110 21586 52162
rect 22542 52110 22594 52162
rect 22990 52110 23042 52162
rect 23214 52110 23266 52162
rect 23774 52110 23826 52162
rect 24222 52110 24274 52162
rect 24670 52110 24722 52162
rect 24894 52110 24946 52162
rect 28926 52110 28978 52162
rect 29710 52110 29762 52162
rect 30158 52110 30210 52162
rect 31166 52110 31218 52162
rect 34638 52110 34690 52162
rect 39790 52110 39842 52162
rect 41134 52110 41186 52162
rect 46174 52110 46226 52162
rect 46622 52110 46674 52162
rect 52782 52110 52834 52162
rect 53566 52110 53618 52162
rect 53902 52110 53954 52162
rect 10446 51998 10498 52050
rect 10894 51998 10946 52050
rect 14814 51998 14866 52050
rect 14926 51998 14978 52050
rect 26910 51998 26962 52050
rect 27134 51998 27186 52050
rect 27358 51998 27410 52050
rect 27470 51998 27522 52050
rect 33294 51998 33346 52050
rect 45950 51998 46002 52050
rect 52446 51998 52498 52050
rect 2606 51886 2658 51938
rect 3950 51886 4002 51938
rect 5630 51886 5682 51938
rect 7646 51886 7698 51938
rect 23102 51886 23154 51938
rect 24446 51886 24498 51938
rect 25118 51886 25170 51938
rect 25230 51886 25282 51938
rect 26014 51886 26066 51938
rect 27918 51886 27970 51938
rect 28478 51886 28530 51938
rect 32174 51886 32226 51938
rect 52558 51886 52610 51938
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 2270 51550 2322 51602
rect 3166 51550 3218 51602
rect 4846 51550 4898 51602
rect 5294 51550 5346 51602
rect 5742 51550 5794 51602
rect 12462 51550 12514 51602
rect 15710 51550 15762 51602
rect 15822 51550 15874 51602
rect 17838 51550 17890 51602
rect 18846 51550 18898 51602
rect 21198 51550 21250 51602
rect 22094 51550 22146 51602
rect 23550 51550 23602 51602
rect 29150 51550 29202 51602
rect 33854 51550 33906 51602
rect 36654 51550 36706 51602
rect 37550 51550 37602 51602
rect 42142 51550 42194 51602
rect 55134 51550 55186 51602
rect 8878 51438 8930 51490
rect 13022 51438 13074 51490
rect 19406 51438 19458 51490
rect 22990 51438 23042 51490
rect 25902 51438 25954 51490
rect 28254 51438 28306 51490
rect 29374 51438 29426 51490
rect 39454 51438 39506 51490
rect 42254 51438 42306 51490
rect 45950 51438 46002 51490
rect 47854 51438 47906 51490
rect 52334 51438 52386 51490
rect 3614 51326 3666 51378
rect 6190 51326 6242 51378
rect 6638 51326 6690 51378
rect 6862 51326 6914 51378
rect 7534 51326 7586 51378
rect 7758 51326 7810 51378
rect 7982 51326 8034 51378
rect 8654 51326 8706 51378
rect 8990 51326 9042 51378
rect 10446 51326 10498 51378
rect 10670 51326 10722 51378
rect 10894 51326 10946 51378
rect 11118 51326 11170 51378
rect 11342 51326 11394 51378
rect 14254 51326 14306 51378
rect 15598 51326 15650 51378
rect 15934 51326 15986 51378
rect 18286 51326 18338 51378
rect 18622 51326 18674 51378
rect 20078 51326 20130 51378
rect 23214 51326 23266 51378
rect 24334 51326 24386 51378
rect 24558 51326 24610 51378
rect 25006 51326 25058 51378
rect 26126 51326 26178 51378
rect 27806 51326 27858 51378
rect 29486 51326 29538 51378
rect 30270 51326 30322 51378
rect 32398 51326 32450 51378
rect 32622 51326 32674 51378
rect 33742 51326 33794 51378
rect 33966 51326 34018 51378
rect 34078 51326 34130 51378
rect 36206 51326 36258 51378
rect 36542 51326 36594 51378
rect 36878 51326 36930 51378
rect 37326 51326 37378 51378
rect 39006 51326 39058 51378
rect 39342 51326 39394 51378
rect 43150 51326 43202 51378
rect 44046 51326 44098 51378
rect 44942 51326 44994 51378
rect 47182 51326 47234 51378
rect 51886 51326 51938 51378
rect 1934 51214 1986 51266
rect 2718 51214 2770 51266
rect 4062 51214 4114 51266
rect 6750 51214 6802 51266
rect 7870 51214 7922 51266
rect 13918 51214 13970 51266
rect 16942 51214 16994 51266
rect 18958 51214 19010 51266
rect 19742 51214 19794 51266
rect 21646 51214 21698 51266
rect 24446 51214 24498 51266
rect 27470 51214 27522 51266
rect 28702 51214 28754 51266
rect 30718 51214 30770 51266
rect 31054 51214 31106 51266
rect 32734 51214 32786 51266
rect 34638 51214 34690 51266
rect 39902 51214 39954 51266
rect 43262 51214 43314 51266
rect 45838 51214 45890 51266
rect 51550 51214 51602 51266
rect 55694 51214 55746 51266
rect 56254 51214 56306 51266
rect 58046 51214 58098 51266
rect 58382 51214 58434 51266
rect 1710 51102 1762 51154
rect 2718 51102 2770 51154
rect 11566 51102 11618 51154
rect 12126 51102 12178 51154
rect 12798 51102 12850 51154
rect 16270 51102 16322 51154
rect 21198 51102 21250 51154
rect 22206 51102 22258 51154
rect 26462 51102 26514 51154
rect 34414 51102 34466 51154
rect 37662 51102 37714 51154
rect 42030 51102 42082 51154
rect 45054 51102 45106 51154
rect 55470 51102 55522 51154
rect 57710 51102 57762 51154
rect 58382 51102 58434 51154
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 6302 50766 6354 50818
rect 12126 50766 12178 50818
rect 16382 50766 16434 50818
rect 16718 50766 16770 50818
rect 21870 50766 21922 50818
rect 23662 50766 23714 50818
rect 31278 50766 31330 50818
rect 32062 50766 32114 50818
rect 32510 50766 32562 50818
rect 33406 50766 33458 50818
rect 39342 50766 39394 50818
rect 39678 50766 39730 50818
rect 41918 50766 41970 50818
rect 42926 50766 42978 50818
rect 46286 50766 46338 50818
rect 51550 50766 51602 50818
rect 55918 50766 55970 50818
rect 58158 50766 58210 50818
rect 2606 50654 2658 50706
rect 2942 50654 2994 50706
rect 4510 50654 4562 50706
rect 6862 50654 6914 50706
rect 7758 50654 7810 50706
rect 12238 50654 12290 50706
rect 12910 50654 12962 50706
rect 13918 50654 13970 50706
rect 18174 50654 18226 50706
rect 19182 50654 19234 50706
rect 19966 50654 20018 50706
rect 21870 50654 21922 50706
rect 22318 50654 22370 50706
rect 23662 50654 23714 50706
rect 27022 50654 27074 50706
rect 27358 50654 27410 50706
rect 27918 50654 27970 50706
rect 30158 50654 30210 50706
rect 30606 50654 30658 50706
rect 32510 50654 32562 50706
rect 36430 50654 36482 50706
rect 37662 50654 37714 50706
rect 38558 50654 38610 50706
rect 40238 50654 40290 50706
rect 41806 50654 41858 50706
rect 43150 50654 43202 50706
rect 46062 50654 46114 50706
rect 48526 50654 48578 50706
rect 50654 50654 50706 50706
rect 2158 50542 2210 50594
rect 4062 50542 4114 50594
rect 6638 50542 6690 50594
rect 6974 50542 7026 50594
rect 9102 50542 9154 50594
rect 9886 50542 9938 50594
rect 10894 50542 10946 50594
rect 14030 50542 14082 50594
rect 14142 50542 14194 50594
rect 14478 50542 14530 50594
rect 14702 50542 14754 50594
rect 15150 50542 15202 50594
rect 20302 50542 20354 50594
rect 23326 50542 23378 50594
rect 24558 50542 24610 50594
rect 24894 50542 24946 50594
rect 26910 50542 26962 50594
rect 29934 50542 29986 50594
rect 31390 50542 31442 50594
rect 33406 50542 33458 50594
rect 36318 50542 36370 50594
rect 36766 50542 36818 50594
rect 37886 50542 37938 50594
rect 39118 50542 39170 50594
rect 40574 50542 40626 50594
rect 41022 50542 41074 50594
rect 41582 50542 41634 50594
rect 43374 50542 43426 50594
rect 46734 50542 46786 50594
rect 47070 50542 47122 50594
rect 49982 50542 50034 50594
rect 54238 50542 54290 50594
rect 54462 50542 54514 50594
rect 56142 50542 56194 50594
rect 56366 50542 56418 50594
rect 56814 50542 56866 50594
rect 57262 50542 57314 50594
rect 57486 50542 57538 50594
rect 5070 50430 5122 50482
rect 7646 50430 7698 50482
rect 7870 50430 7922 50482
rect 8766 50430 8818 50482
rect 9774 50430 9826 50482
rect 12350 50430 12402 50482
rect 13806 50430 13858 50482
rect 15598 50430 15650 50482
rect 15822 50430 15874 50482
rect 16494 50430 16546 50482
rect 20862 50430 20914 50482
rect 25118 50430 25170 50482
rect 25790 50430 25842 50482
rect 28030 50430 28082 50482
rect 28254 50430 28306 50482
rect 28814 50430 28866 50482
rect 31278 50430 31330 50482
rect 32062 50430 32114 50482
rect 33070 50430 33122 50482
rect 35198 50430 35250 50482
rect 40350 50430 40402 50482
rect 48974 50430 49026 50482
rect 51774 50430 51826 50482
rect 54126 50430 54178 50482
rect 58046 50430 58098 50482
rect 3502 50318 3554 50370
rect 5742 50318 5794 50370
rect 6750 50318 6802 50370
rect 11006 50318 11058 50370
rect 11342 50318 11394 50370
rect 15486 50318 15538 50370
rect 17614 50318 17666 50370
rect 18734 50318 18786 50370
rect 22766 50318 22818 50370
rect 25006 50318 25058 50370
rect 33854 50318 33906 50370
rect 34302 50318 34354 50370
rect 34750 50318 34802 50370
rect 46062 50318 46114 50370
rect 46958 50318 47010 50370
rect 51214 50318 51266 50370
rect 53566 50318 53618 50370
rect 56254 50318 56306 50370
rect 57150 50318 57202 50370
rect 58158 50318 58210 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 3390 49982 3442 50034
rect 4958 49982 5010 50034
rect 5630 49982 5682 50034
rect 8318 49982 8370 50034
rect 10222 49982 10274 50034
rect 10558 49982 10610 50034
rect 11454 49982 11506 50034
rect 11678 49982 11730 50034
rect 12686 49982 12738 50034
rect 14254 49982 14306 50034
rect 15710 49982 15762 50034
rect 17838 49982 17890 50034
rect 18062 49982 18114 50034
rect 19294 49982 19346 50034
rect 25678 49982 25730 50034
rect 26686 49982 26738 50034
rect 29598 49982 29650 50034
rect 30382 49982 30434 50034
rect 30494 49982 30546 50034
rect 31950 49982 32002 50034
rect 32622 49982 32674 50034
rect 36094 49982 36146 50034
rect 39790 49982 39842 50034
rect 43262 49982 43314 50034
rect 45950 49982 46002 50034
rect 52558 49982 52610 50034
rect 53118 49982 53170 50034
rect 57598 49982 57650 50034
rect 57822 49982 57874 50034
rect 4734 49870 4786 49922
rect 7982 49870 8034 49922
rect 12462 49870 12514 49922
rect 17726 49870 17778 49922
rect 19854 49870 19906 49922
rect 29486 49870 29538 49922
rect 31726 49870 31778 49922
rect 39678 49870 39730 49922
rect 39902 49870 39954 49922
rect 40350 49870 40402 49922
rect 58382 49870 58434 49922
rect 58494 49870 58546 49922
rect 2382 49758 2434 49810
rect 3950 49758 4002 49810
rect 6974 49758 7026 49810
rect 8318 49758 8370 49810
rect 8542 49758 8594 49810
rect 10110 49758 10162 49810
rect 10334 49758 10386 49810
rect 11790 49758 11842 49810
rect 12350 49758 12402 49810
rect 13134 49758 13186 49810
rect 13358 49758 13410 49810
rect 13806 49758 13858 49810
rect 18510 49758 18562 49810
rect 20526 49758 20578 49810
rect 20750 49758 20802 49810
rect 23550 49758 23602 49810
rect 27246 49758 27298 49810
rect 27918 49758 27970 49810
rect 29710 49758 29762 49810
rect 30270 49758 30322 49810
rect 30942 49758 30994 49810
rect 31614 49758 31666 49810
rect 32398 49758 32450 49810
rect 33966 49758 34018 49810
rect 34526 49758 34578 49810
rect 42030 49758 42082 49810
rect 45726 49758 45778 49810
rect 46062 49758 46114 49810
rect 48190 49758 48242 49810
rect 49534 49758 49586 49810
rect 52222 49758 52274 49810
rect 52334 49758 52386 49810
rect 55470 49758 55522 49810
rect 55694 49758 55746 49810
rect 57486 49758 57538 49810
rect 58158 49758 58210 49810
rect 2046 49646 2098 49698
rect 2942 49646 2994 49698
rect 6078 49646 6130 49698
rect 7310 49646 7362 49698
rect 8990 49646 9042 49698
rect 13246 49646 13298 49698
rect 14814 49646 14866 49698
rect 15822 49646 15874 49698
rect 16494 49646 16546 49698
rect 16942 49646 16994 49698
rect 22542 49646 22594 49698
rect 23774 49646 23826 49698
rect 24782 49646 24834 49698
rect 26126 49646 26178 49698
rect 27022 49646 27074 49698
rect 28366 49646 28418 49698
rect 28814 49646 28866 49698
rect 34638 49646 34690 49698
rect 35534 49646 35586 49698
rect 35758 49646 35810 49698
rect 36542 49646 36594 49698
rect 37102 49646 37154 49698
rect 37550 49646 37602 49698
rect 41918 49646 41970 49698
rect 42590 49646 42642 49698
rect 43822 49646 43874 49698
rect 49758 49646 49810 49698
rect 50878 49646 50930 49698
rect 51438 49646 51490 49698
rect 52446 49646 52498 49698
rect 53790 49646 53842 49698
rect 55918 49646 55970 49698
rect 56702 49646 56754 49698
rect 2046 49534 2098 49586
rect 3166 49534 3218 49586
rect 5070 49534 5122 49586
rect 10894 49534 10946 49586
rect 11006 49534 11058 49586
rect 14590 49534 14642 49586
rect 15486 49534 15538 49586
rect 25566 49534 25618 49586
rect 26126 49534 26178 49586
rect 32734 49534 32786 49586
rect 43598 49534 43650 49586
rect 48414 49534 48466 49586
rect 48750 49534 48802 49586
rect 50094 49534 50146 49586
rect 51886 49534 51938 49586
rect 56366 49534 56418 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 1934 49198 1986 49250
rect 2606 49198 2658 49250
rect 3054 49198 3106 49250
rect 5742 49198 5794 49250
rect 13918 49198 13970 49250
rect 14478 49198 14530 49250
rect 22878 49198 22930 49250
rect 30718 49198 30770 49250
rect 42142 49198 42194 49250
rect 44606 49198 44658 49250
rect 47182 49198 47234 49250
rect 52670 49198 52722 49250
rect 55470 49198 55522 49250
rect 1934 49086 1986 49138
rect 3838 49086 3890 49138
rect 4958 49086 5010 49138
rect 7310 49086 7362 49138
rect 9214 49086 9266 49138
rect 11454 49086 11506 49138
rect 12350 49086 12402 49138
rect 13918 49086 13970 49138
rect 14366 49086 14418 49138
rect 16942 49086 16994 49138
rect 17390 49086 17442 49138
rect 18398 49086 18450 49138
rect 20862 49086 20914 49138
rect 22654 49086 22706 49138
rect 24894 49086 24946 49138
rect 26350 49086 26402 49138
rect 27918 49086 27970 49138
rect 28366 49086 28418 49138
rect 28814 49086 28866 49138
rect 30494 49086 30546 49138
rect 35758 49086 35810 49138
rect 36542 49086 36594 49138
rect 38334 49086 38386 49138
rect 46734 49086 46786 49138
rect 49534 49086 49586 49138
rect 51774 49086 51826 49138
rect 54126 49086 54178 49138
rect 56478 49086 56530 49138
rect 57038 49086 57090 49138
rect 9886 48974 9938 49026
rect 9998 48974 10050 49026
rect 10334 48974 10386 49026
rect 12126 48974 12178 49026
rect 12798 48974 12850 49026
rect 14926 48974 14978 49026
rect 15262 48974 15314 49026
rect 15598 48974 15650 49026
rect 18062 48974 18114 49026
rect 19630 48974 19682 49026
rect 20078 48974 20130 49026
rect 21982 48974 22034 49026
rect 23102 48974 23154 49026
rect 23774 48974 23826 49026
rect 24222 48974 24274 49026
rect 24782 48974 24834 49026
rect 25006 48974 25058 49026
rect 25230 48974 25282 49026
rect 30718 48974 30770 49026
rect 32622 48974 32674 49026
rect 32958 48974 33010 49026
rect 34414 48974 34466 49026
rect 34862 48974 34914 49026
rect 36094 48974 36146 49026
rect 44718 48974 44770 49026
rect 46398 48974 46450 49026
rect 48974 48974 49026 49026
rect 49422 48974 49474 49026
rect 49646 48974 49698 49026
rect 51662 48974 51714 49026
rect 51998 48974 52050 49026
rect 52558 48974 52610 49026
rect 53678 48974 53730 49026
rect 56702 48974 56754 49026
rect 57598 48974 57650 49026
rect 57822 48974 57874 49026
rect 58270 48974 58322 49026
rect 6974 48862 7026 48914
rect 18174 48862 18226 48914
rect 21646 48862 21698 48914
rect 21758 48862 21810 48914
rect 25454 48862 25506 48914
rect 39566 48862 39618 48914
rect 41806 48862 41858 48914
rect 43262 48862 43314 48914
rect 43374 48862 43426 48914
rect 52334 48862 52386 48914
rect 53342 48862 53394 48914
rect 53566 48862 53618 48914
rect 55358 48862 55410 48914
rect 2382 48750 2434 48802
rect 2830 48750 2882 48802
rect 3278 48750 3330 48802
rect 4622 48750 4674 48802
rect 5854 48750 5906 48802
rect 5966 48750 6018 48802
rect 7198 48750 7250 48802
rect 7422 48750 7474 48802
rect 7870 48750 7922 48802
rect 8430 48750 8482 48802
rect 8878 48750 8930 48802
rect 10110 48750 10162 48802
rect 11006 48750 11058 48802
rect 12574 48750 12626 48802
rect 12686 48750 12738 48802
rect 15038 48750 15090 48802
rect 16046 48750 16098 48802
rect 16494 48750 16546 48802
rect 18398 48750 18450 48802
rect 18510 48750 18562 48802
rect 26014 48750 26066 48802
rect 26798 48750 26850 48802
rect 27582 48750 27634 48802
rect 37550 48750 37602 48802
rect 37886 48750 37938 48802
rect 39230 48750 39282 48802
rect 39454 48750 39506 48802
rect 42030 48750 42082 48802
rect 43598 48750 43650 48802
rect 44606 48750 44658 48802
rect 51102 48750 51154 48802
rect 55470 48750 55522 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 2046 48414 2098 48466
rect 2830 48414 2882 48466
rect 3390 48414 3442 48466
rect 8766 48414 8818 48466
rect 9774 48414 9826 48466
rect 11790 48414 11842 48466
rect 12238 48414 12290 48466
rect 14590 48414 14642 48466
rect 15710 48414 15762 48466
rect 16942 48414 16994 48466
rect 19294 48414 19346 48466
rect 21086 48414 21138 48466
rect 22654 48414 22706 48466
rect 23438 48414 23490 48466
rect 25790 48414 25842 48466
rect 49534 48414 49586 48466
rect 52558 48414 52610 48466
rect 53118 48414 53170 48466
rect 5406 48302 5458 48354
rect 15486 48302 15538 48354
rect 16158 48302 16210 48354
rect 20862 48302 20914 48354
rect 21534 48302 21586 48354
rect 23326 48302 23378 48354
rect 26574 48302 26626 48354
rect 33630 48302 33682 48354
rect 40462 48302 40514 48354
rect 43822 48302 43874 48354
rect 46622 48302 46674 48354
rect 52670 48302 52722 48354
rect 57486 48302 57538 48354
rect 5182 48190 5234 48242
rect 6750 48190 6802 48242
rect 7534 48190 7586 48242
rect 8430 48190 8482 48242
rect 9774 48190 9826 48242
rect 10110 48190 10162 48242
rect 10222 48190 10274 48242
rect 10558 48190 10610 48242
rect 11342 48190 11394 48242
rect 12798 48190 12850 48242
rect 12910 48190 12962 48242
rect 13134 48190 13186 48242
rect 13358 48190 13410 48242
rect 14142 48190 14194 48242
rect 14366 48190 14418 48242
rect 14814 48190 14866 48242
rect 15934 48190 15986 48242
rect 17950 48190 18002 48242
rect 20190 48190 20242 48242
rect 20750 48190 20802 48242
rect 21758 48190 21810 48242
rect 23550 48190 23602 48242
rect 23998 48190 24050 48242
rect 28254 48190 28306 48242
rect 30046 48190 30098 48242
rect 30830 48190 30882 48242
rect 31166 48190 31218 48242
rect 33854 48190 33906 48242
rect 34078 48190 34130 48242
rect 35982 48190 36034 48242
rect 36430 48190 36482 48242
rect 37886 48190 37938 48242
rect 38110 48190 38162 48242
rect 39566 48190 39618 48242
rect 43150 48190 43202 48242
rect 46174 48190 46226 48242
rect 46510 48190 46562 48242
rect 51662 48190 51714 48242
rect 51998 48190 52050 48242
rect 52446 48190 52498 48242
rect 54798 48190 54850 48242
rect 55358 48190 55410 48242
rect 57598 48190 57650 48242
rect 57934 48190 57986 48242
rect 2382 48078 2434 48130
rect 3950 48078 4002 48130
rect 14478 48078 14530 48130
rect 16270 48078 16322 48130
rect 17838 48078 17890 48130
rect 23774 48078 23826 48130
rect 24446 48078 24498 48130
rect 24894 48078 24946 48130
rect 28142 48078 28194 48130
rect 29934 48078 29986 48130
rect 35646 48078 35698 48130
rect 36990 48078 37042 48130
rect 38782 48078 38834 48130
rect 39678 48078 39730 48130
rect 43374 48078 43426 48130
rect 49646 48078 49698 48130
rect 50206 48078 50258 48130
rect 50654 48078 50706 48130
rect 51214 48078 51266 48130
rect 55694 48078 55746 48130
rect 56702 48078 56754 48130
rect 18398 47966 18450 48018
rect 27918 47966 27970 48018
rect 50878 47966 50930 48018
rect 52222 47966 52274 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 3838 47630 3890 47682
rect 9326 47630 9378 47682
rect 9774 47630 9826 47682
rect 12014 47630 12066 47682
rect 12910 47630 12962 47682
rect 26126 47630 26178 47682
rect 26574 47630 26626 47682
rect 26798 47630 26850 47682
rect 34526 47630 34578 47682
rect 36206 47630 36258 47682
rect 52222 47630 52274 47682
rect 2830 47518 2882 47570
rect 3502 47518 3554 47570
rect 7310 47518 7362 47570
rect 7534 47518 7586 47570
rect 8654 47518 8706 47570
rect 11454 47518 11506 47570
rect 12014 47518 12066 47570
rect 13022 47518 13074 47570
rect 15150 47518 15202 47570
rect 17614 47518 17666 47570
rect 18062 47518 18114 47570
rect 20078 47518 20130 47570
rect 21982 47518 22034 47570
rect 22878 47518 22930 47570
rect 26126 47518 26178 47570
rect 26574 47518 26626 47570
rect 27246 47518 27298 47570
rect 28366 47518 28418 47570
rect 28814 47518 28866 47570
rect 31278 47518 31330 47570
rect 32958 47518 33010 47570
rect 38558 47518 38610 47570
rect 40798 47518 40850 47570
rect 42478 47518 42530 47570
rect 45614 47518 45666 47570
rect 46734 47518 46786 47570
rect 55358 47518 55410 47570
rect 56366 47518 56418 47570
rect 2606 47406 2658 47458
rect 4174 47406 4226 47458
rect 6078 47406 6130 47458
rect 7086 47406 7138 47458
rect 7646 47406 7698 47458
rect 9438 47406 9490 47458
rect 9998 47406 10050 47458
rect 10670 47406 10722 47458
rect 15710 47406 15762 47458
rect 15934 47406 15986 47458
rect 16270 47406 16322 47458
rect 17278 47406 17330 47458
rect 18174 47406 18226 47458
rect 19854 47406 19906 47458
rect 20638 47406 20690 47458
rect 23326 47406 23378 47458
rect 27134 47406 27186 47458
rect 27358 47406 27410 47458
rect 31726 47406 31778 47458
rect 33182 47406 33234 47458
rect 34078 47406 34130 47458
rect 34526 47406 34578 47458
rect 36206 47406 36258 47458
rect 37438 47406 37490 47458
rect 38446 47406 38498 47458
rect 39118 47406 39170 47458
rect 41022 47406 41074 47458
rect 41582 47406 41634 47458
rect 41806 47406 41858 47458
rect 44046 47406 44098 47458
rect 44606 47406 44658 47458
rect 45390 47406 45442 47458
rect 46062 47406 46114 47458
rect 51662 47406 51714 47458
rect 51886 47406 51938 47458
rect 54574 47406 54626 47458
rect 55246 47406 55298 47458
rect 56814 47406 56866 47458
rect 3390 47294 3442 47346
rect 3614 47294 3666 47346
rect 9214 47294 9266 47346
rect 10894 47294 10946 47346
rect 11006 47294 11058 47346
rect 11118 47294 11170 47346
rect 18510 47294 18562 47346
rect 19294 47294 19346 47346
rect 20190 47294 20242 47346
rect 24558 47294 24610 47346
rect 27582 47294 27634 47346
rect 36542 47294 36594 47346
rect 39454 47294 39506 47346
rect 40350 47294 40402 47346
rect 40574 47294 40626 47346
rect 44718 47294 44770 47346
rect 45838 47294 45890 47346
rect 46622 47294 46674 47346
rect 46846 47294 46898 47346
rect 48190 47294 48242 47346
rect 56254 47294 56306 47346
rect 56590 47294 56642 47346
rect 1822 47182 1874 47234
rect 2270 47182 2322 47234
rect 4958 47182 5010 47234
rect 12462 47182 12514 47234
rect 13694 47182 13746 47234
rect 14478 47182 14530 47234
rect 15822 47182 15874 47234
rect 20078 47182 20130 47234
rect 21646 47182 21698 47234
rect 22430 47182 22482 47234
rect 23774 47182 23826 47234
rect 24334 47182 24386 47234
rect 24446 47182 24498 47234
rect 24782 47182 24834 47234
rect 25678 47182 25730 47234
rect 29710 47182 29762 47234
rect 37998 47182 38050 47234
rect 38670 47182 38722 47234
rect 48302 47182 48354 47234
rect 48526 47182 48578 47234
rect 48862 47182 48914 47234
rect 51102 47182 51154 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 2382 46846 2434 46898
rect 3166 46846 3218 46898
rect 4846 46846 4898 46898
rect 6078 46846 6130 46898
rect 6862 46846 6914 46898
rect 8766 46846 8818 46898
rect 10670 46846 10722 46898
rect 11454 46846 11506 46898
rect 12910 46846 12962 46898
rect 14142 46846 14194 46898
rect 16942 46846 16994 46898
rect 22990 46846 23042 46898
rect 32622 46846 32674 46898
rect 33630 46846 33682 46898
rect 36654 46846 36706 46898
rect 38110 46846 38162 46898
rect 38446 46846 38498 46898
rect 45614 46846 45666 46898
rect 49646 46846 49698 46898
rect 49982 46846 50034 46898
rect 3390 46734 3442 46786
rect 3502 46734 3554 46786
rect 4734 46734 4786 46786
rect 4958 46734 5010 46786
rect 6638 46734 6690 46786
rect 7646 46734 7698 46786
rect 8990 46734 9042 46786
rect 10334 46734 10386 46786
rect 10558 46734 10610 46786
rect 14254 46734 14306 46786
rect 14366 46734 14418 46786
rect 18510 46734 18562 46786
rect 21198 46734 21250 46786
rect 23774 46734 23826 46786
rect 36206 46734 36258 46786
rect 36878 46734 36930 46786
rect 37886 46734 37938 46786
rect 40014 46734 40066 46786
rect 45502 46734 45554 46786
rect 53230 46734 53282 46786
rect 55694 46734 55746 46786
rect 57486 46734 57538 46786
rect 2830 46622 2882 46674
rect 6974 46622 7026 46674
rect 7198 46622 7250 46674
rect 10782 46622 10834 46674
rect 11790 46622 11842 46674
rect 12350 46622 12402 46674
rect 12798 46622 12850 46674
rect 13022 46622 13074 46674
rect 13918 46622 13970 46674
rect 15262 46622 15314 46674
rect 16606 46622 16658 46674
rect 17838 46622 17890 46674
rect 19854 46622 19906 46674
rect 21310 46622 21362 46674
rect 23550 46622 23602 46674
rect 23998 46622 24050 46674
rect 24222 46622 24274 46674
rect 26238 46622 26290 46674
rect 28254 46622 28306 46674
rect 29934 46622 29986 46674
rect 30158 46622 30210 46674
rect 30606 46622 30658 46674
rect 30830 46622 30882 46674
rect 34190 46622 34242 46674
rect 35758 46622 35810 46674
rect 36990 46622 37042 46674
rect 37774 46622 37826 46674
rect 39566 46622 39618 46674
rect 47854 46622 47906 46674
rect 48750 46622 48802 46674
rect 49534 46622 49586 46674
rect 49758 46622 49810 46674
rect 55246 46622 55298 46674
rect 55470 46622 55522 46674
rect 55918 46622 55970 46674
rect 58158 46622 58210 46674
rect 1934 46510 1986 46562
rect 4174 46510 4226 46562
rect 5630 46510 5682 46562
rect 8094 46510 8146 46562
rect 8878 46510 8930 46562
rect 9774 46510 9826 46562
rect 14702 46510 14754 46562
rect 15822 46510 15874 46562
rect 16382 46510 16434 46562
rect 20414 46510 20466 46562
rect 22542 46510 22594 46562
rect 23886 46510 23938 46562
rect 25006 46510 25058 46562
rect 27806 46510 27858 46562
rect 35870 46510 35922 46562
rect 39230 46510 39282 46562
rect 42590 46510 42642 46562
rect 47070 46510 47122 46562
rect 47966 46510 48018 46562
rect 53118 46510 53170 46562
rect 54014 46510 54066 46562
rect 56478 46510 56530 46562
rect 57822 46510 57874 46562
rect 11454 46398 11506 46450
rect 11566 46398 11618 46450
rect 25678 46398 25730 46450
rect 26014 46398 26066 46450
rect 29374 46398 29426 46450
rect 33966 46398 34018 46450
rect 53454 46398 53506 46450
rect 56030 46398 56082 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 3614 46062 3666 46114
rect 30942 46062 30994 46114
rect 31726 46062 31778 46114
rect 38558 46062 38610 46114
rect 39342 46062 39394 46114
rect 39678 46062 39730 46114
rect 43150 46062 43202 46114
rect 46734 46062 46786 46114
rect 55582 46062 55634 46114
rect 57486 46062 57538 46114
rect 57822 46062 57874 46114
rect 1934 45950 1986 46002
rect 6750 45950 6802 46002
rect 9774 45950 9826 46002
rect 12126 45950 12178 46002
rect 12686 45950 12738 46002
rect 15262 45950 15314 46002
rect 22878 45950 22930 46002
rect 26910 45950 26962 46002
rect 29598 45950 29650 46002
rect 31166 45950 31218 46002
rect 31614 45950 31666 46002
rect 33406 45950 33458 46002
rect 34190 45950 34242 46002
rect 35646 45950 35698 46002
rect 37998 45950 38050 46002
rect 41246 45950 41298 46002
rect 44718 45950 44770 46002
rect 45614 45950 45666 46002
rect 48750 45950 48802 46002
rect 54462 45950 54514 46002
rect 56142 45950 56194 46002
rect 56590 45950 56642 46002
rect 2830 45838 2882 45890
rect 3278 45838 3330 45890
rect 6526 45838 6578 45890
rect 6638 45838 6690 45890
rect 7534 45838 7586 45890
rect 7982 45838 8034 45890
rect 8766 45838 8818 45890
rect 9102 45838 9154 45890
rect 10334 45838 10386 45890
rect 14702 45838 14754 45890
rect 15374 45838 15426 45890
rect 17390 45838 17442 45890
rect 18174 45838 18226 45890
rect 18510 45838 18562 45890
rect 20526 45838 20578 45890
rect 22654 45838 22706 45890
rect 23326 45838 23378 45890
rect 24334 45838 24386 45890
rect 25454 45838 25506 45890
rect 30718 45838 30770 45890
rect 33518 45838 33570 45890
rect 34302 45838 34354 45890
rect 34750 45838 34802 45890
rect 36206 45838 36258 45890
rect 37774 45838 37826 45890
rect 41694 45838 41746 45890
rect 42142 45838 42194 45890
rect 42814 45838 42866 45890
rect 45726 45838 45778 45890
rect 45950 45838 46002 45890
rect 48974 45838 49026 45890
rect 51326 45838 51378 45890
rect 51550 45838 51602 45890
rect 53790 45838 53842 45890
rect 54238 45838 54290 45890
rect 55918 45838 55970 45890
rect 58046 45838 58098 45890
rect 2494 45726 2546 45778
rect 4398 45726 4450 45778
rect 4510 45726 4562 45778
rect 7086 45726 7138 45778
rect 8206 45726 8258 45778
rect 10894 45726 10946 45778
rect 13918 45726 13970 45778
rect 14030 45726 14082 45778
rect 16046 45726 16098 45778
rect 20190 45726 20242 45778
rect 24222 45726 24274 45778
rect 24782 45726 24834 45778
rect 25566 45726 25618 45778
rect 25790 45726 25842 45778
rect 26798 45726 26850 45778
rect 27134 45726 27186 45778
rect 27358 45726 27410 45778
rect 29710 45726 29762 45778
rect 29934 45726 29986 45778
rect 30606 45726 30658 45778
rect 33070 45726 33122 45778
rect 34078 45726 34130 45778
rect 35758 45726 35810 45778
rect 40238 45726 40290 45778
rect 43038 45726 43090 45778
rect 45502 45726 45554 45778
rect 46622 45726 46674 45778
rect 49646 45726 49698 45778
rect 4734 45614 4786 45666
rect 5854 45614 5906 45666
rect 6862 45614 6914 45666
rect 7758 45614 7810 45666
rect 8878 45614 8930 45666
rect 14254 45614 14306 45666
rect 19854 45614 19906 45666
rect 21534 45614 21586 45666
rect 22094 45614 22146 45666
rect 23102 45614 23154 45666
rect 23214 45614 23266 45666
rect 24558 45614 24610 45666
rect 24670 45614 24722 45666
rect 25342 45614 25394 45666
rect 28030 45614 28082 45666
rect 28366 45614 28418 45666
rect 28926 45614 28978 45666
rect 30382 45614 30434 45666
rect 32174 45614 32226 45666
rect 33294 45614 33346 45666
rect 35534 45614 35586 45666
rect 36654 45614 36706 45666
rect 39566 45614 39618 45666
rect 40574 45614 40626 45666
rect 44158 45614 44210 45666
rect 46734 45614 46786 45666
rect 51886 45614 51938 45666
rect 54910 45614 54962 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 3054 45278 3106 45330
rect 4398 45278 4450 45330
rect 5182 45278 5234 45330
rect 5406 45278 5458 45330
rect 7198 45278 7250 45330
rect 10782 45278 10834 45330
rect 15598 45278 15650 45330
rect 16942 45278 16994 45330
rect 18286 45278 18338 45330
rect 23998 45278 24050 45330
rect 24110 45278 24162 45330
rect 25006 45278 25058 45330
rect 29486 45278 29538 45330
rect 30270 45278 30322 45330
rect 30494 45278 30546 45330
rect 30606 45278 30658 45330
rect 31726 45278 31778 45330
rect 34638 45278 34690 45330
rect 34750 45278 34802 45330
rect 37102 45278 37154 45330
rect 38446 45278 38498 45330
rect 38782 45278 38834 45330
rect 41470 45278 41522 45330
rect 42814 45278 42866 45330
rect 44494 45278 44546 45330
rect 45054 45278 45106 45330
rect 45166 45278 45218 45330
rect 53566 45278 53618 45330
rect 57934 45278 57986 45330
rect 2158 45166 2210 45218
rect 4174 45166 4226 45218
rect 11342 45166 11394 45218
rect 12798 45166 12850 45218
rect 14814 45166 14866 45218
rect 17838 45166 17890 45218
rect 20974 45166 21026 45218
rect 21646 45166 21698 45218
rect 27246 45166 27298 45218
rect 27582 45166 27634 45218
rect 29374 45166 29426 45218
rect 30830 45166 30882 45218
rect 31614 45166 31666 45218
rect 36654 45166 36706 45218
rect 38222 45166 38274 45218
rect 39790 45166 39842 45218
rect 43598 45166 43650 45218
rect 44158 45166 44210 45218
rect 44270 45166 44322 45218
rect 47518 45166 47570 45218
rect 52894 45166 52946 45218
rect 54014 45166 54066 45218
rect 56366 45166 56418 45218
rect 57598 45166 57650 45218
rect 2494 45054 2546 45106
rect 5070 45054 5122 45106
rect 6638 45054 6690 45106
rect 6862 45054 6914 45106
rect 7198 45054 7250 45106
rect 7646 45054 7698 45106
rect 8094 45054 8146 45106
rect 10782 45054 10834 45106
rect 11678 45054 11730 45106
rect 12574 45054 12626 45106
rect 14478 45054 14530 45106
rect 18062 45054 18114 45106
rect 20190 45054 20242 45106
rect 20862 45054 20914 45106
rect 21758 45054 21810 45106
rect 23774 45054 23826 45106
rect 24222 45054 24274 45106
rect 24334 45054 24386 45106
rect 25678 45054 25730 45106
rect 26910 45054 26962 45106
rect 27694 45054 27746 45106
rect 27806 45054 27858 45106
rect 28590 45054 28642 45106
rect 28814 45054 28866 45106
rect 29262 45054 29314 45106
rect 30382 45054 30434 45106
rect 31390 45054 31442 45106
rect 32062 45054 32114 45106
rect 34526 45054 34578 45106
rect 34862 45054 34914 45106
rect 35086 45054 35138 45106
rect 35758 45054 35810 45106
rect 35982 45054 36034 45106
rect 38110 45054 38162 45106
rect 39678 45054 39730 45106
rect 40014 45054 40066 45106
rect 42254 45054 42306 45106
rect 42702 45054 42754 45106
rect 42926 45054 42978 45106
rect 47070 45054 47122 45106
rect 48750 45054 48802 45106
rect 49870 45054 49922 45106
rect 51998 45054 52050 45106
rect 53342 45054 53394 45106
rect 53790 45054 53842 45106
rect 57822 45054 57874 45106
rect 58046 45054 58098 45106
rect 58494 45054 58546 45106
rect 2382 44942 2434 44994
rect 3614 44942 3666 44994
rect 4510 44942 4562 44994
rect 6078 44942 6130 44994
rect 8654 44942 8706 44994
rect 9662 44942 9714 44994
rect 10222 44942 10274 44994
rect 16158 44942 16210 44994
rect 16494 44942 16546 44994
rect 18846 44942 18898 44994
rect 19294 44942 19346 44994
rect 21534 44942 21586 44994
rect 22766 44942 22818 44994
rect 23214 44942 23266 44994
rect 29038 44942 29090 44994
rect 32510 44942 32562 44994
rect 32958 44942 33010 44994
rect 33630 44942 33682 44994
rect 37550 44942 37602 44994
rect 40350 44942 40402 44994
rect 45726 44942 45778 44994
rect 46622 44942 46674 44994
rect 48526 44942 48578 44994
rect 49646 44942 49698 44994
rect 50542 44942 50594 44994
rect 52110 44942 52162 44994
rect 56254 44942 56306 44994
rect 7086 44830 7138 44882
rect 25678 44830 25730 44882
rect 26014 44830 26066 44882
rect 27022 44830 27074 44882
rect 45278 44830 45330 44882
rect 48190 44830 48242 44882
rect 56590 44830 56642 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 6190 44494 6242 44546
rect 6862 44494 6914 44546
rect 24558 44494 24610 44546
rect 24670 44494 24722 44546
rect 24894 44494 24946 44546
rect 25006 44494 25058 44546
rect 27694 44494 27746 44546
rect 28142 44494 28194 44546
rect 28590 44494 28642 44546
rect 28814 44494 28866 44546
rect 30046 44494 30098 44546
rect 36094 44494 36146 44546
rect 56702 44494 56754 44546
rect 3166 44382 3218 44434
rect 4398 44382 4450 44434
rect 10670 44382 10722 44434
rect 13806 44382 13858 44434
rect 14926 44382 14978 44434
rect 20862 44382 20914 44434
rect 25790 44382 25842 44434
rect 27918 44382 27970 44434
rect 30382 44382 30434 44434
rect 35982 44382 36034 44434
rect 37886 44382 37938 44434
rect 39902 44382 39954 44434
rect 40238 44382 40290 44434
rect 44270 44382 44322 44434
rect 45838 44382 45890 44434
rect 48302 44382 48354 44434
rect 49086 44382 49138 44434
rect 49758 44382 49810 44434
rect 51102 44382 51154 44434
rect 51998 44382 52050 44434
rect 56590 44382 56642 44434
rect 57710 44382 57762 44434
rect 2718 44270 2770 44322
rect 2942 44270 2994 44322
rect 4286 44270 4338 44322
rect 5966 44270 6018 44322
rect 6414 44270 6466 44322
rect 8430 44270 8482 44322
rect 10334 44270 10386 44322
rect 11230 44270 11282 44322
rect 11790 44270 11842 44322
rect 12014 44270 12066 44322
rect 14366 44270 14418 44322
rect 14814 44270 14866 44322
rect 15822 44270 15874 44322
rect 16046 44270 16098 44322
rect 17726 44270 17778 44322
rect 18174 44270 18226 44322
rect 18286 44270 18338 44322
rect 19070 44270 19122 44322
rect 21646 44270 21698 44322
rect 21870 44270 21922 44322
rect 22094 44270 22146 44322
rect 22206 44270 22258 44322
rect 26462 44270 26514 44322
rect 27022 44270 27074 44322
rect 27470 44270 27522 44322
rect 31502 44270 31554 44322
rect 31838 44270 31890 44322
rect 33406 44270 33458 44322
rect 34750 44270 34802 44322
rect 35310 44270 35362 44322
rect 38222 44270 38274 44322
rect 38782 44270 38834 44322
rect 41246 44270 41298 44322
rect 41582 44270 41634 44322
rect 42590 44270 42642 44322
rect 42814 44270 42866 44322
rect 44158 44270 44210 44322
rect 44382 44270 44434 44322
rect 46174 44270 46226 44322
rect 46622 44270 46674 44322
rect 48414 44270 48466 44322
rect 49870 44270 49922 44322
rect 50094 44270 50146 44322
rect 51326 44270 51378 44322
rect 56814 44270 56866 44322
rect 4062 44158 4114 44210
rect 4958 44158 5010 44210
rect 5742 44158 5794 44210
rect 8990 44158 9042 44210
rect 9214 44158 9266 44210
rect 10446 44158 10498 44210
rect 14926 44158 14978 44210
rect 19182 44158 19234 44210
rect 19518 44158 19570 44210
rect 20302 44158 20354 44210
rect 20414 44158 20466 44210
rect 20526 44158 20578 44210
rect 26350 44158 26402 44210
rect 29486 44158 29538 44210
rect 30158 44158 30210 44210
rect 39678 44158 39730 44210
rect 41358 44158 41410 44210
rect 43486 44158 43538 44210
rect 44718 44158 44770 44210
rect 49646 44158 49698 44210
rect 7422 44046 7474 44098
rect 7870 44046 7922 44098
rect 8542 44046 8594 44098
rect 11902 44046 11954 44098
rect 14590 44046 14642 44098
rect 16382 44046 16434 44098
rect 16830 44046 16882 44098
rect 17278 44046 17330 44098
rect 18398 44046 18450 44098
rect 19406 44046 19458 44098
rect 20078 44046 20130 44098
rect 22094 44046 22146 44098
rect 22990 44046 23042 44098
rect 23550 44046 23602 44098
rect 23886 44046 23938 44098
rect 26574 44046 26626 44098
rect 27582 44046 27634 44098
rect 28814 44046 28866 44098
rect 30830 44046 30882 44098
rect 42030 44046 42082 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 1934 43710 1986 43762
rect 5294 43710 5346 43762
rect 8206 43710 8258 43762
rect 9886 43710 9938 43762
rect 12574 43710 12626 43762
rect 14702 43710 14754 43762
rect 16830 43710 16882 43762
rect 17950 43710 18002 43762
rect 26014 43710 26066 43762
rect 26462 43710 26514 43762
rect 28030 43710 28082 43762
rect 28142 43710 28194 43762
rect 28254 43710 28306 43762
rect 30270 43710 30322 43762
rect 35422 43710 35474 43762
rect 38222 43710 38274 43762
rect 44494 43710 44546 43762
rect 45502 43710 45554 43762
rect 56590 43710 56642 43762
rect 5070 43598 5122 43650
rect 5406 43598 5458 43650
rect 9774 43598 9826 43650
rect 10446 43598 10498 43650
rect 11454 43598 11506 43650
rect 12238 43598 12290 43650
rect 12350 43598 12402 43650
rect 13470 43598 13522 43650
rect 16270 43598 16322 43650
rect 16606 43598 16658 43650
rect 18062 43598 18114 43650
rect 20862 43598 20914 43650
rect 23998 43598 24050 43650
rect 24558 43598 24610 43650
rect 28478 43598 28530 43650
rect 31054 43598 31106 43650
rect 34526 43598 34578 43650
rect 39678 43598 39730 43650
rect 40350 43598 40402 43650
rect 43934 43598 43986 43650
rect 56366 43598 56418 43650
rect 57486 43598 57538 43650
rect 3166 43486 3218 43538
rect 3726 43486 3778 43538
rect 5518 43486 5570 43538
rect 6750 43486 6802 43538
rect 7646 43486 7698 43538
rect 10670 43486 10722 43538
rect 12014 43486 12066 43538
rect 12910 43486 12962 43538
rect 14366 43486 14418 43538
rect 14702 43486 14754 43538
rect 15038 43486 15090 43538
rect 16382 43486 16434 43538
rect 17726 43486 17778 43538
rect 18734 43486 18786 43538
rect 18958 43486 19010 43538
rect 20414 43486 20466 43538
rect 21646 43486 21698 43538
rect 27918 43486 27970 43538
rect 32846 43486 32898 43538
rect 34302 43486 34354 43538
rect 35086 43486 35138 43538
rect 35982 43486 36034 43538
rect 37326 43486 37378 43538
rect 40574 43486 40626 43538
rect 41582 43486 41634 43538
rect 42254 43486 42306 43538
rect 54126 43486 54178 43538
rect 55022 43486 55074 43538
rect 56030 43486 56082 43538
rect 56254 43486 56306 43538
rect 56478 43486 56530 43538
rect 57934 43486 57986 43538
rect 2494 43374 2546 43426
rect 4174 43374 4226 43426
rect 6302 43374 6354 43426
rect 7198 43374 7250 43426
rect 8542 43374 8594 43426
rect 8990 43374 9042 43426
rect 9998 43374 10050 43426
rect 13022 43374 13074 43426
rect 13918 43374 13970 43426
rect 15486 43374 15538 43426
rect 16494 43374 16546 43426
rect 18846 43374 18898 43426
rect 19182 43374 19234 43426
rect 19406 43374 19458 43426
rect 21086 43374 21138 43426
rect 21198 43374 21250 43426
rect 22766 43374 22818 43426
rect 23102 43374 23154 43426
rect 23662 43374 23714 43426
rect 25006 43374 25058 43426
rect 26798 43374 26850 43426
rect 27246 43374 27298 43426
rect 29262 43374 29314 43426
rect 29710 43374 29762 43426
rect 33518 43374 33570 43426
rect 36542 43374 36594 43426
rect 36878 43374 36930 43426
rect 37886 43374 37938 43426
rect 38670 43374 38722 43426
rect 39118 43374 39170 43426
rect 40798 43374 40850 43426
rect 42366 43374 42418 43426
rect 44046 43374 44098 43426
rect 44942 43374 44994 43426
rect 46062 43374 46114 43426
rect 46622 43374 46674 43426
rect 46958 43374 47010 43426
rect 47406 43374 47458 43426
rect 47854 43374 47906 43426
rect 48414 43374 48466 43426
rect 48862 43374 48914 43426
rect 54910 43374 54962 43426
rect 58382 43374 58434 43426
rect 4062 43262 4114 43314
rect 7198 43262 7250 43314
rect 8878 43262 8930 43314
rect 10222 43262 10274 43314
rect 19630 43262 19682 43314
rect 23662 43262 23714 43314
rect 25118 43262 25170 43314
rect 31278 43262 31330 43314
rect 31614 43262 31666 43314
rect 32510 43262 32562 43314
rect 32846 43262 32898 43314
rect 38782 43262 38834 43314
rect 39118 43262 39170 43314
rect 42814 43262 42866 43314
rect 43710 43262 43762 43314
rect 44270 43262 44322 43314
rect 45054 43262 45106 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 6638 42926 6690 42978
rect 12126 42926 12178 42978
rect 22094 42926 22146 42978
rect 27694 42926 27746 42978
rect 28254 42926 28306 42978
rect 29934 42926 29986 42978
rect 36206 42926 36258 42978
rect 45502 42926 45554 42978
rect 45838 42926 45890 42978
rect 48974 42926 49026 42978
rect 2158 42814 2210 42866
rect 2606 42814 2658 42866
rect 2942 42814 2994 42866
rect 3614 42814 3666 42866
rect 10334 42814 10386 42866
rect 14254 42814 14306 42866
rect 15150 42814 15202 42866
rect 15934 42814 15986 42866
rect 17838 42814 17890 42866
rect 18398 42814 18450 42866
rect 18734 42814 18786 42866
rect 25118 42814 25170 42866
rect 25902 42814 25954 42866
rect 26686 42814 26738 42866
rect 27918 42814 27970 42866
rect 35758 42814 35810 42866
rect 40462 42814 40514 42866
rect 47742 42814 47794 42866
rect 53902 42814 53954 42866
rect 55022 42814 55074 42866
rect 56702 42814 56754 42866
rect 4062 42702 4114 42754
rect 6078 42702 6130 42754
rect 6414 42702 6466 42754
rect 6862 42702 6914 42754
rect 8094 42702 8146 42754
rect 8542 42702 8594 42754
rect 8766 42702 8818 42754
rect 8990 42702 9042 42754
rect 9214 42702 9266 42754
rect 11790 42702 11842 42754
rect 13918 42702 13970 42754
rect 14366 42702 14418 42754
rect 15710 42702 15762 42754
rect 17054 42702 17106 42754
rect 17726 42702 17778 42754
rect 21982 42702 22034 42754
rect 22206 42702 22258 42754
rect 23662 42702 23714 42754
rect 23998 42702 24050 42754
rect 26126 42702 26178 42754
rect 26798 42702 26850 42754
rect 28814 42702 28866 42754
rect 31950 42702 32002 42754
rect 33070 42702 33122 42754
rect 33294 42702 33346 42754
rect 34414 42702 34466 42754
rect 35310 42702 35362 42754
rect 38110 42702 38162 42754
rect 38894 42702 38946 42754
rect 39118 42702 39170 42754
rect 46062 42702 46114 42754
rect 48750 42702 48802 42754
rect 53342 42702 53394 42754
rect 54014 42702 54066 42754
rect 55582 42702 55634 42754
rect 55918 42702 55970 42754
rect 7758 42590 7810 42642
rect 7870 42590 7922 42642
rect 9886 42590 9938 42642
rect 11118 42590 11170 42642
rect 11566 42590 11618 42642
rect 13694 42590 13746 42642
rect 14142 42590 14194 42642
rect 16046 42590 16098 42642
rect 16158 42590 16210 42642
rect 17278 42590 17330 42642
rect 17390 42590 17442 42642
rect 19966 42590 20018 42642
rect 21646 42590 21698 42642
rect 23102 42590 23154 42642
rect 25902 42590 25954 42642
rect 30046 42590 30098 42642
rect 37774 42590 37826 42642
rect 39790 42590 39842 42642
rect 40350 42590 40402 42642
rect 54910 42590 54962 42642
rect 56254 42590 56306 42642
rect 3502 42478 3554 42530
rect 3726 42478 3778 42530
rect 4622 42478 4674 42530
rect 5070 42478 5122 42530
rect 6526 42478 6578 42530
rect 8878 42478 8930 42530
rect 13022 42478 13074 42530
rect 15934 42478 15986 42530
rect 18622 42478 18674 42530
rect 19518 42478 19570 42530
rect 20414 42478 20466 42530
rect 20862 42478 20914 42530
rect 22430 42478 22482 42530
rect 26350 42478 26402 42530
rect 27470 42478 27522 42530
rect 28366 42478 28418 42530
rect 29934 42478 29986 42530
rect 30830 42478 30882 42530
rect 37886 42478 37938 42530
rect 40574 42478 40626 42530
rect 40798 42478 40850 42530
rect 41358 42478 41410 42530
rect 41806 42478 41858 42530
rect 42702 42478 42754 42530
rect 43374 42478 43426 42530
rect 44718 42478 44770 42530
rect 46510 42478 46562 42530
rect 47406 42478 47458 42530
rect 47630 42478 47682 42530
rect 47854 42478 47906 42530
rect 48302 42478 48354 42530
rect 49086 42478 49138 42530
rect 49310 42478 49362 42530
rect 49758 42478 49810 42530
rect 52222 42478 52274 42530
rect 53790 42478 53842 42530
rect 55134 42478 55186 42530
rect 56142 42478 56194 42530
rect 57150 42478 57202 42530
rect 57598 42478 57650 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 3726 42142 3778 42194
rect 10110 42142 10162 42194
rect 10670 42142 10722 42194
rect 13358 42142 13410 42194
rect 13470 42142 13522 42194
rect 13582 42142 13634 42194
rect 14926 42142 14978 42194
rect 17950 42142 18002 42194
rect 19518 42142 19570 42194
rect 19630 42142 19682 42194
rect 32846 42142 32898 42194
rect 37438 42142 37490 42194
rect 37550 42142 37602 42194
rect 37662 42142 37714 42194
rect 38446 42142 38498 42194
rect 44718 42142 44770 42194
rect 53342 42142 53394 42194
rect 2494 42030 2546 42082
rect 2718 42030 2770 42082
rect 3054 42030 3106 42082
rect 3614 42030 3666 42082
rect 6638 42030 6690 42082
rect 8766 42030 8818 42082
rect 21758 42030 21810 42082
rect 26574 42030 26626 42082
rect 29598 42030 29650 42082
rect 30830 42030 30882 42082
rect 31166 42030 31218 42082
rect 36542 42030 36594 42082
rect 37102 42030 37154 42082
rect 37326 42030 37378 42082
rect 38334 42030 38386 42082
rect 42366 42030 42418 42082
rect 48750 42030 48802 42082
rect 53902 42030 53954 42082
rect 57486 42030 57538 42082
rect 3950 41918 4002 41970
rect 4174 41918 4226 41970
rect 6526 41918 6578 41970
rect 7422 41918 7474 41970
rect 8542 41918 8594 41970
rect 9662 41918 9714 41970
rect 11230 41918 11282 41970
rect 12014 41918 12066 41970
rect 12910 41918 12962 41970
rect 14142 41918 14194 41970
rect 14590 41918 14642 41970
rect 14814 41918 14866 41970
rect 15038 41918 15090 41970
rect 15598 41918 15650 41970
rect 16494 41918 16546 41970
rect 19294 41918 19346 41970
rect 19742 41918 19794 41970
rect 19854 41918 19906 41970
rect 20862 41918 20914 41970
rect 21086 41918 21138 41970
rect 21870 41918 21922 41970
rect 21982 41918 22034 41970
rect 22430 41918 22482 41970
rect 22878 41918 22930 41970
rect 23662 41918 23714 41970
rect 24222 41918 24274 41970
rect 26686 41918 26738 41970
rect 28366 41918 28418 41970
rect 29038 41918 29090 41970
rect 30718 41918 30770 41970
rect 33854 41918 33906 41970
rect 34078 41918 34130 41970
rect 35870 41918 35922 41970
rect 38670 41918 38722 41970
rect 40126 41918 40178 41970
rect 43374 41918 43426 41970
rect 44606 41918 44658 41970
rect 44942 41918 44994 41970
rect 45726 41918 45778 41970
rect 46398 41918 46450 41970
rect 48302 41918 48354 41970
rect 48638 41918 48690 41970
rect 50094 41918 50146 41970
rect 51102 41918 51154 41970
rect 52670 41918 52722 41970
rect 56366 41918 56418 41970
rect 57598 41918 57650 41970
rect 57934 41918 57986 41970
rect 1710 41806 1762 41858
rect 2046 41806 2098 41858
rect 2942 41806 2994 41858
rect 4958 41806 5010 41858
rect 5518 41806 5570 41858
rect 5966 41806 6018 41858
rect 6974 41806 7026 41858
rect 7198 41806 7250 41858
rect 8878 41806 8930 41858
rect 12574 41806 12626 41858
rect 14366 41806 14418 41858
rect 16046 41806 16098 41858
rect 16942 41806 16994 41858
rect 17838 41806 17890 41858
rect 18846 41806 18898 41858
rect 24110 41806 24162 41858
rect 25902 41806 25954 41858
rect 27694 41806 27746 41858
rect 28926 41806 28978 41858
rect 31054 41806 31106 41858
rect 31726 41806 31778 41858
rect 32286 41806 32338 41858
rect 35646 41806 35698 41858
rect 39342 41806 39394 41858
rect 39790 41806 39842 41858
rect 41470 41806 41522 41858
rect 43150 41806 43202 41858
rect 43822 41806 43874 41858
rect 45278 41806 45330 41858
rect 49982 41806 50034 41858
rect 56254 41806 56306 41858
rect 2382 41694 2434 41746
rect 17726 41694 17778 41746
rect 20526 41694 20578 41746
rect 24558 41694 24610 41746
rect 32510 41694 32562 41746
rect 34526 41694 34578 41746
rect 42142 41694 42194 41746
rect 42478 41694 42530 41746
rect 43038 41694 43090 41746
rect 46622 41694 46674 41746
rect 46846 41694 46898 41746
rect 47294 41694 47346 41746
rect 51774 41694 51826 41746
rect 52446 41694 52498 41746
rect 53006 41694 53058 41746
rect 53230 41694 53282 41746
rect 54014 41694 54066 41746
rect 54238 41694 54290 41746
rect 54462 41694 54514 41746
rect 54574 41694 54626 41746
rect 55918 41694 55970 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 2270 41358 2322 41410
rect 2830 41358 2882 41410
rect 3054 41358 3106 41410
rect 3614 41358 3666 41410
rect 6974 41358 7026 41410
rect 8878 41358 8930 41410
rect 10558 41358 10610 41410
rect 11118 41358 11170 41410
rect 12014 41358 12066 41410
rect 12798 41358 12850 41410
rect 14814 41358 14866 41410
rect 17390 41358 17442 41410
rect 17614 41358 17666 41410
rect 24446 41358 24498 41410
rect 24670 41358 24722 41410
rect 27918 41358 27970 41410
rect 28030 41358 28082 41410
rect 28254 41358 28306 41410
rect 34190 41358 34242 41410
rect 34526 41358 34578 41410
rect 44494 41358 44546 41410
rect 48638 41358 48690 41410
rect 50206 41358 50258 41410
rect 53790 41358 53842 41410
rect 54350 41358 54402 41410
rect 54686 41358 54738 41410
rect 3838 41246 3890 41298
rect 7086 41246 7138 41298
rect 9886 41246 9938 41298
rect 11566 41246 11618 41298
rect 12462 41246 12514 41298
rect 15486 41246 15538 41298
rect 17390 41246 17442 41298
rect 17726 41246 17778 41298
rect 18622 41246 18674 41298
rect 19630 41246 19682 41298
rect 20190 41246 20242 41298
rect 20862 41246 20914 41298
rect 23214 41246 23266 41298
rect 23774 41246 23826 41298
rect 28814 41246 28866 41298
rect 30942 41246 30994 41298
rect 36542 41246 36594 41298
rect 39566 41246 39618 41298
rect 46958 41246 47010 41298
rect 53678 41246 53730 41298
rect 54910 41246 54962 41298
rect 55358 41246 55410 41298
rect 56590 41246 56642 41298
rect 57262 41246 57314 41298
rect 3278 41134 3330 41186
rect 4510 41134 4562 41186
rect 5630 41134 5682 41186
rect 8990 41134 9042 41186
rect 9550 41134 9602 41186
rect 10670 41134 10722 41186
rect 14142 41134 14194 41186
rect 19294 41134 19346 41186
rect 19406 41134 19458 41186
rect 24334 41134 24386 41186
rect 27246 41134 27298 41186
rect 29934 41134 29986 41186
rect 32286 41134 32338 41186
rect 33630 41134 33682 41186
rect 35982 41134 36034 41186
rect 36206 41134 36258 41186
rect 36430 41134 36482 41186
rect 37662 41134 37714 41186
rect 37886 41134 37938 41186
rect 39454 41134 39506 41186
rect 39678 41134 39730 41186
rect 40014 41134 40066 41186
rect 40462 41134 40514 41186
rect 43934 41134 43986 41186
rect 46174 41134 46226 41186
rect 48078 41134 48130 41186
rect 49198 41134 49250 41186
rect 49422 41134 49474 41186
rect 53902 41134 53954 41186
rect 54126 41134 54178 41186
rect 57150 41134 57202 41186
rect 57374 41134 57426 41186
rect 2606 41022 2658 41074
rect 6078 41022 6130 41074
rect 7422 41022 7474 41074
rect 9214 41022 9266 41074
rect 9774 41022 9826 41074
rect 12910 41022 12962 41074
rect 14254 41022 14306 41074
rect 14366 41022 14418 41074
rect 16942 41022 16994 41074
rect 19742 41022 19794 41074
rect 25230 41022 25282 41074
rect 26462 41022 26514 41074
rect 26798 41022 26850 41074
rect 30158 41022 30210 41074
rect 33518 41022 33570 41074
rect 38558 41022 38610 41074
rect 40798 41022 40850 41074
rect 43598 41022 43650 41074
rect 44382 41022 44434 41074
rect 47406 41022 47458 41074
rect 50094 41022 50146 41074
rect 2046 40910 2098 40962
rect 3950 40910 4002 40962
rect 5070 40910 5122 40962
rect 8318 40910 8370 40962
rect 11230 40910 11282 40962
rect 12014 40910 12066 40962
rect 15934 40910 15986 40962
rect 16382 40910 16434 40962
rect 18174 40910 18226 40962
rect 21534 40910 21586 40962
rect 22318 40910 22370 40962
rect 22766 40910 22818 40962
rect 27134 40910 27186 40962
rect 32846 40910 32898 40962
rect 35198 40910 35250 40962
rect 36654 40910 36706 40962
rect 40686 40910 40738 40962
rect 41246 40910 41298 40962
rect 41806 40910 41858 40962
rect 42142 40910 42194 40962
rect 42702 40910 42754 40962
rect 43150 40910 43202 40962
rect 43710 40910 43762 40962
rect 44494 40910 44546 40962
rect 45502 40910 45554 40962
rect 50206 40910 50258 40962
rect 50766 40910 50818 40962
rect 51214 40910 51266 40962
rect 51886 40910 51938 40962
rect 52670 40910 52722 40962
rect 53566 40910 53618 40962
rect 55806 40910 55858 40962
rect 57598 40910 57650 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 2942 40574 2994 40626
rect 4286 40574 4338 40626
rect 4734 40574 4786 40626
rect 5518 40574 5570 40626
rect 6414 40574 6466 40626
rect 6974 40574 7026 40626
rect 8878 40574 8930 40626
rect 11678 40574 11730 40626
rect 13694 40574 13746 40626
rect 13918 40574 13970 40626
rect 14478 40574 14530 40626
rect 15038 40574 15090 40626
rect 17726 40574 17778 40626
rect 18734 40574 18786 40626
rect 19182 40574 19234 40626
rect 19630 40574 19682 40626
rect 21310 40574 21362 40626
rect 21422 40574 21474 40626
rect 22206 40574 22258 40626
rect 25566 40574 25618 40626
rect 27806 40574 27858 40626
rect 28030 40574 28082 40626
rect 29038 40574 29090 40626
rect 30830 40574 30882 40626
rect 32286 40574 32338 40626
rect 35982 40574 36034 40626
rect 37774 40574 37826 40626
rect 42590 40574 42642 40626
rect 50990 40574 51042 40626
rect 54126 40574 54178 40626
rect 54462 40574 54514 40626
rect 57486 40574 57538 40626
rect 1822 40462 1874 40514
rect 5742 40462 5794 40514
rect 11230 40462 11282 40514
rect 11454 40462 11506 40514
rect 13022 40462 13074 40514
rect 15262 40462 15314 40514
rect 16382 40462 16434 40514
rect 16494 40462 16546 40514
rect 16942 40462 16994 40514
rect 22654 40462 22706 40514
rect 24894 40462 24946 40514
rect 27694 40462 27746 40514
rect 29598 40462 29650 40514
rect 31502 40462 31554 40514
rect 38446 40462 38498 40514
rect 43038 40462 43090 40514
rect 46846 40462 46898 40514
rect 48302 40462 48354 40514
rect 48526 40462 48578 40514
rect 50766 40462 50818 40514
rect 57710 40462 57762 40514
rect 58270 40462 58322 40514
rect 2270 40350 2322 40402
rect 5070 40350 5122 40402
rect 5854 40350 5906 40402
rect 7758 40350 7810 40402
rect 8318 40350 8370 40402
rect 8766 40350 8818 40402
rect 8990 40350 9042 40402
rect 10558 40350 10610 40402
rect 12014 40350 12066 40402
rect 12126 40350 12178 40402
rect 13582 40350 13634 40402
rect 14366 40350 14418 40402
rect 14702 40350 14754 40402
rect 15374 40350 15426 40402
rect 16606 40350 16658 40402
rect 18062 40350 18114 40402
rect 18510 40350 18562 40402
rect 20750 40350 20802 40402
rect 21198 40350 21250 40402
rect 23326 40350 23378 40402
rect 23662 40350 23714 40402
rect 26574 40350 26626 40402
rect 26798 40350 26850 40402
rect 27134 40350 27186 40402
rect 29822 40350 29874 40402
rect 32846 40350 32898 40402
rect 33518 40350 33570 40402
rect 34302 40350 34354 40402
rect 34526 40350 34578 40402
rect 34638 40350 34690 40402
rect 36430 40350 36482 40402
rect 37326 40350 37378 40402
rect 38894 40350 38946 40402
rect 39230 40350 39282 40402
rect 40014 40350 40066 40402
rect 42142 40350 42194 40402
rect 44270 40350 44322 40402
rect 45614 40350 45666 40402
rect 48190 40350 48242 40402
rect 49534 40350 49586 40402
rect 49982 40350 50034 40402
rect 50654 40350 50706 40402
rect 53566 40350 53618 40402
rect 57822 40350 57874 40402
rect 3502 40238 3554 40290
rect 9774 40238 9826 40290
rect 11118 40238 11170 40290
rect 12574 40238 12626 40290
rect 15934 40238 15986 40290
rect 7086 40126 7138 40178
rect 7310 40126 7362 40178
rect 7870 40126 7922 40178
rect 10222 40126 10274 40178
rect 10558 40126 10610 40178
rect 17502 40126 17554 40178
rect 18174 40238 18226 40290
rect 18622 40238 18674 40290
rect 20078 40238 20130 40290
rect 26126 40238 26178 40290
rect 28702 40238 28754 40290
rect 31390 40238 31442 40290
rect 31726 40238 31778 40290
rect 35646 40238 35698 40290
rect 36878 40238 36930 40290
rect 39902 40238 39954 40290
rect 43822 40238 43874 40290
rect 44606 40238 44658 40290
rect 45726 40238 45778 40290
rect 19518 40126 19570 40178
rect 19966 40126 20018 40178
rect 28702 40126 28754 40178
rect 29150 40126 29202 40178
rect 30158 40126 30210 40178
rect 35086 40126 35138 40178
rect 36206 40126 36258 40178
rect 36878 40126 36930 40178
rect 40238 40126 40290 40178
rect 46062 40126 46114 40178
rect 47070 40126 47122 40178
rect 47406 40126 47458 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 2718 39790 2770 39842
rect 3502 39790 3554 39842
rect 4734 39790 4786 39842
rect 9774 39790 9826 39842
rect 11566 39790 11618 39842
rect 34750 39790 34802 39842
rect 42814 39790 42866 39842
rect 2494 39678 2546 39730
rect 3614 39678 3666 39730
rect 4062 39678 4114 39730
rect 4958 39678 5010 39730
rect 5630 39678 5682 39730
rect 7758 39678 7810 39730
rect 8766 39678 8818 39730
rect 9214 39678 9266 39730
rect 10782 39678 10834 39730
rect 12910 39678 12962 39730
rect 15038 39678 15090 39730
rect 16158 39678 16210 39730
rect 18622 39678 18674 39730
rect 19966 39678 20018 39730
rect 22878 39678 22930 39730
rect 25118 39678 25170 39730
rect 25678 39678 25730 39730
rect 27246 39678 27298 39730
rect 28478 39678 28530 39730
rect 34414 39678 34466 39730
rect 38558 39678 38610 39730
rect 40462 39678 40514 39730
rect 41134 39678 41186 39730
rect 42030 39678 42082 39730
rect 42590 39678 42642 39730
rect 43150 39678 43202 39730
rect 43822 39678 43874 39730
rect 45502 39678 45554 39730
rect 50878 39678 50930 39730
rect 7646 39566 7698 39618
rect 7870 39566 7922 39618
rect 9886 39566 9938 39618
rect 10446 39566 10498 39618
rect 10670 39566 10722 39618
rect 11790 39566 11842 39618
rect 12014 39566 12066 39618
rect 14590 39566 14642 39618
rect 14926 39566 14978 39618
rect 15374 39566 15426 39618
rect 16718 39566 16770 39618
rect 16830 39566 16882 39618
rect 17614 39566 17666 39618
rect 18286 39566 18338 39618
rect 19406 39566 19458 39618
rect 20974 39566 21026 39618
rect 21758 39566 21810 39618
rect 22318 39566 22370 39618
rect 23550 39566 23602 39618
rect 23886 39566 23938 39618
rect 27022 39566 27074 39618
rect 29822 39566 29874 39618
rect 30494 39566 30546 39618
rect 31726 39566 31778 39618
rect 32174 39566 32226 39618
rect 35086 39566 35138 39618
rect 36094 39566 36146 39618
rect 36430 39566 36482 39618
rect 41582 39566 41634 39618
rect 44270 39566 44322 39618
rect 45726 39566 45778 39618
rect 47294 39566 47346 39618
rect 50318 39566 50370 39618
rect 51438 39566 51490 39618
rect 53902 39566 53954 39618
rect 57150 39566 57202 39618
rect 57374 39566 57426 39618
rect 57822 39566 57874 39618
rect 4622 39454 4674 39506
rect 6190 39454 6242 39506
rect 6302 39454 6354 39506
rect 7422 39454 7474 39506
rect 10110 39454 10162 39506
rect 11454 39454 11506 39506
rect 12462 39454 12514 39506
rect 17166 39454 17218 39506
rect 17390 39454 17442 39506
rect 18734 39454 18786 39506
rect 19854 39454 19906 39506
rect 21870 39454 21922 39506
rect 35870 39454 35922 39506
rect 44718 39454 44770 39506
rect 47070 39454 47122 39506
rect 49982 39454 50034 39506
rect 53566 39454 53618 39506
rect 54686 39454 54738 39506
rect 2046 39342 2098 39394
rect 3054 39342 3106 39394
rect 6526 39342 6578 39394
rect 8318 39342 8370 39394
rect 13582 39342 13634 39394
rect 14030 39342 14082 39394
rect 15150 39342 15202 39394
rect 17502 39342 17554 39394
rect 18510 39342 18562 39394
rect 18846 39342 18898 39394
rect 20078 39342 20130 39394
rect 22094 39342 22146 39394
rect 26126 39342 26178 39394
rect 35982 39342 36034 39394
rect 46062 39342 46114 39394
rect 46510 39342 46562 39394
rect 48638 39342 48690 39394
rect 50094 39342 50146 39394
rect 50766 39342 50818 39394
rect 50990 39342 51042 39394
rect 53678 39342 53730 39394
rect 54350 39342 54402 39394
rect 54574 39342 54626 39394
rect 56590 39342 56642 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 2382 39006 2434 39058
rect 3726 39006 3778 39058
rect 3838 39006 3890 39058
rect 8990 39006 9042 39058
rect 12462 39006 12514 39058
rect 13246 39006 13298 39058
rect 13694 39006 13746 39058
rect 14590 39006 14642 39058
rect 15486 39006 15538 39058
rect 15710 39006 15762 39058
rect 16046 39006 16098 39058
rect 16718 39006 16770 39058
rect 16830 39006 16882 39058
rect 22654 39006 22706 39058
rect 23102 39006 23154 39058
rect 28590 39006 28642 39058
rect 34078 39006 34130 39058
rect 36318 39006 36370 39058
rect 36654 39006 36706 39058
rect 37102 39006 37154 39058
rect 37550 39006 37602 39058
rect 42030 39006 42082 39058
rect 42590 39006 42642 39058
rect 42926 39006 42978 39058
rect 45502 39006 45554 39058
rect 46734 39006 46786 39058
rect 47182 39006 47234 39058
rect 56478 39006 56530 39058
rect 3614 38894 3666 38946
rect 4622 38894 4674 38946
rect 4846 38894 4898 38946
rect 5182 38894 5234 38946
rect 7310 38894 7362 38946
rect 8206 38894 8258 38946
rect 10894 38894 10946 38946
rect 14478 38894 14530 38946
rect 14814 38894 14866 38946
rect 15374 38894 15426 38946
rect 17726 38894 17778 38946
rect 17950 38894 18002 38946
rect 18286 38894 18338 38946
rect 19518 38894 19570 38946
rect 20638 38894 20690 38946
rect 23998 38894 24050 38946
rect 27806 38894 27858 38946
rect 29150 38894 29202 38946
rect 33630 38894 33682 38946
rect 33854 38894 33906 38946
rect 40798 38894 40850 38946
rect 52222 38894 52274 38946
rect 58494 38894 58546 38946
rect 2046 38782 2098 38834
rect 2606 38782 2658 38834
rect 3166 38782 3218 38834
rect 6078 38782 6130 38834
rect 6414 38782 6466 38834
rect 6750 38782 6802 38834
rect 7646 38782 7698 38834
rect 7758 38782 7810 38834
rect 10334 38782 10386 38834
rect 10670 38782 10722 38834
rect 11790 38782 11842 38834
rect 12014 38782 12066 38834
rect 12350 38782 12402 38834
rect 12686 38782 12738 38834
rect 14254 38782 14306 38834
rect 19182 38782 19234 38834
rect 19406 38782 19458 38834
rect 20526 38782 20578 38834
rect 21534 38782 21586 38834
rect 23550 38782 23602 38834
rect 25790 38782 25842 38834
rect 26014 38782 26066 38834
rect 29710 38782 29762 38834
rect 30046 38782 30098 38834
rect 30718 38782 30770 38834
rect 31726 38782 31778 38834
rect 34190 38782 34242 38834
rect 35534 38782 35586 38834
rect 35982 38782 36034 38834
rect 40126 38782 40178 38834
rect 44942 38782 44994 38834
rect 48078 38782 48130 38834
rect 49870 38782 49922 38834
rect 50430 38782 50482 38834
rect 50542 38782 50594 38834
rect 51326 38782 51378 38834
rect 53790 38782 53842 38834
rect 54798 38782 54850 38834
rect 56702 38782 56754 38834
rect 57934 38782 57986 38834
rect 2494 38670 2546 38722
rect 3390 38670 3442 38722
rect 5070 38670 5122 38722
rect 5630 38670 5682 38722
rect 6302 38670 6354 38722
rect 7982 38670 8034 38722
rect 8094 38670 8146 38722
rect 9774 38670 9826 38722
rect 10782 38670 10834 38722
rect 12574 38670 12626 38722
rect 16606 38670 16658 38722
rect 18174 38670 18226 38722
rect 21198 38670 21250 38722
rect 21310 38670 21362 38722
rect 24558 38670 24610 38722
rect 25006 38670 25058 38722
rect 29822 38670 29874 38722
rect 31502 38670 31554 38722
rect 32622 38670 32674 38722
rect 35198 38670 35250 38722
rect 38334 38670 38386 38722
rect 39342 38670 39394 38722
rect 40350 38670 40402 38722
rect 46286 38670 46338 38722
rect 47966 38670 48018 38722
rect 48750 38670 48802 38722
rect 51438 38670 51490 38722
rect 53902 38670 53954 38722
rect 55582 38670 55634 38722
rect 56366 38670 56418 38722
rect 57598 38670 57650 38722
rect 19966 38558 20018 38610
rect 31390 38558 31442 38610
rect 38446 38558 38498 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 8990 38222 9042 38274
rect 10110 38222 10162 38274
rect 11230 38222 11282 38274
rect 16270 38222 16322 38274
rect 18510 38222 18562 38274
rect 19294 38222 19346 38274
rect 35422 38222 35474 38274
rect 39230 38222 39282 38274
rect 50318 38222 50370 38274
rect 2382 38110 2434 38162
rect 5070 38110 5122 38162
rect 7422 38110 7474 38162
rect 8654 38110 8706 38162
rect 10334 38110 10386 38162
rect 11566 38110 11618 38162
rect 15038 38110 15090 38162
rect 17614 38110 17666 38162
rect 18174 38110 18226 38162
rect 18510 38110 18562 38162
rect 22654 38110 22706 38162
rect 26350 38110 26402 38162
rect 27246 38110 27298 38162
rect 30606 38110 30658 38162
rect 31838 38110 31890 38162
rect 36318 38110 36370 38162
rect 2942 37998 2994 38050
rect 3502 37998 3554 38050
rect 4062 37998 4114 38050
rect 5742 37998 5794 38050
rect 6750 37998 6802 38050
rect 7646 37998 7698 38050
rect 8542 37998 8594 38050
rect 9102 37998 9154 38050
rect 13918 37998 13970 38050
rect 14814 37998 14866 38050
rect 15934 37998 15986 38050
rect 19406 37998 19458 38050
rect 20526 37998 20578 38050
rect 20750 37998 20802 38050
rect 21646 37998 21698 38050
rect 21870 37998 21922 38050
rect 22766 37998 22818 38050
rect 24110 37998 24162 38050
rect 24446 37998 24498 38050
rect 26574 37998 26626 38050
rect 28142 37998 28194 38050
rect 30718 37998 30770 38050
rect 34190 37998 34242 38050
rect 35198 37998 35250 38050
rect 38110 37998 38162 38050
rect 38334 37998 38386 38050
rect 39006 37998 39058 38050
rect 3054 37886 3106 37938
rect 3950 37886 4002 37938
rect 4286 37886 4338 37938
rect 4510 37886 4562 37938
rect 6862 37886 6914 37938
rect 7534 37886 7586 37938
rect 8766 37886 8818 37938
rect 9774 37886 9826 37938
rect 14366 37886 14418 37938
rect 15038 37886 15090 37938
rect 20638 37886 20690 37938
rect 22990 37886 23042 37938
rect 25566 37886 25618 37938
rect 27806 37886 27858 37938
rect 33294 37886 33346 37938
rect 33406 37886 33458 37938
rect 33630 37886 33682 37938
rect 34526 37886 34578 37938
rect 1934 37774 1986 37826
rect 3278 37774 3330 37826
rect 10670 37774 10722 37826
rect 11118 37774 11170 37826
rect 12014 37774 12066 37826
rect 12574 37774 12626 37826
rect 12910 37774 12962 37826
rect 16158 37774 16210 37826
rect 16718 37774 16770 37826
rect 17166 37774 17218 37826
rect 19070 37774 19122 37826
rect 27918 37774 27970 37826
rect 28814 37774 28866 37826
rect 29598 37774 29650 37826
rect 30046 37774 30098 37826
rect 32622 37774 32674 37826
rect 34078 37774 34130 37826
rect 34302 37774 34354 37826
rect 35758 37774 35810 37826
rect 36654 37774 36706 37826
rect 40126 38110 40178 38162
rect 46734 38110 46786 38162
rect 50766 38110 50818 38162
rect 53902 38110 53954 38162
rect 55246 38110 55298 38162
rect 56366 38110 56418 38162
rect 57822 38110 57874 38162
rect 39566 37998 39618 38050
rect 40238 37998 40290 38050
rect 43598 37998 43650 38050
rect 44158 37998 44210 38050
rect 50430 37998 50482 38050
rect 51550 37998 51602 38050
rect 51886 37998 51938 38050
rect 53566 37998 53618 38050
rect 54126 37998 54178 38050
rect 56142 37998 56194 38050
rect 56478 37998 56530 38050
rect 57710 37998 57762 38050
rect 58382 37998 58434 38050
rect 51774 37886 51826 37938
rect 53678 37886 53730 37938
rect 54910 37886 54962 37938
rect 37438 37774 37490 37826
rect 39230 37774 39282 37826
rect 40014 37774 40066 37826
rect 40798 37774 40850 37826
rect 41246 37774 41298 37826
rect 42142 37774 42194 37826
rect 44046 37774 44098 37826
rect 44270 37774 44322 37826
rect 45726 37774 45778 37826
rect 46622 37774 46674 37826
rect 46846 37774 46898 37826
rect 47070 37774 47122 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 1934 37438 1986 37490
rect 10558 37438 10610 37490
rect 12126 37438 12178 37490
rect 17838 37438 17890 37490
rect 17950 37438 18002 37490
rect 19966 37438 20018 37490
rect 21870 37438 21922 37490
rect 22094 37438 22146 37490
rect 23102 37438 23154 37490
rect 23550 37438 23602 37490
rect 23998 37438 24050 37490
rect 24446 37438 24498 37490
rect 24894 37438 24946 37490
rect 25902 37438 25954 37490
rect 29710 37438 29762 37490
rect 32062 37438 32114 37490
rect 35310 37438 35362 37490
rect 38782 37438 38834 37490
rect 39006 37438 39058 37490
rect 41470 37438 41522 37490
rect 54350 37438 54402 37490
rect 54910 37438 54962 37490
rect 57486 37438 57538 37490
rect 3838 37326 3890 37378
rect 4398 37326 4450 37378
rect 8430 37326 8482 37378
rect 9998 37326 10050 37378
rect 11118 37326 11170 37378
rect 11230 37326 11282 37378
rect 13134 37326 13186 37378
rect 14926 37326 14978 37378
rect 18062 37326 18114 37378
rect 18174 37326 18226 37378
rect 18398 37326 18450 37378
rect 20974 37326 21026 37378
rect 21310 37326 21362 37378
rect 27358 37326 27410 37378
rect 29150 37326 29202 37378
rect 29262 37326 29314 37378
rect 34414 37326 34466 37378
rect 36206 37326 36258 37378
rect 38110 37326 38162 37378
rect 38670 37326 38722 37378
rect 45054 37326 45106 37378
rect 57710 37326 57762 37378
rect 57822 37326 57874 37378
rect 3278 37214 3330 37266
rect 3726 37214 3778 37266
rect 4734 37214 4786 37266
rect 7086 37214 7138 37266
rect 7422 37214 7474 37266
rect 8206 37214 8258 37266
rect 9774 37214 9826 37266
rect 10558 37214 10610 37266
rect 12686 37214 12738 37266
rect 12798 37214 12850 37266
rect 13358 37214 13410 37266
rect 13582 37214 13634 37266
rect 14814 37214 14866 37266
rect 15822 37214 15874 37266
rect 16494 37214 16546 37266
rect 20750 37214 20802 37266
rect 21086 37214 21138 37266
rect 21982 37214 22034 37266
rect 22430 37214 22482 37266
rect 26350 37214 26402 37266
rect 27470 37214 27522 37266
rect 27806 37214 27858 37266
rect 29038 37214 29090 37266
rect 31502 37214 31554 37266
rect 31726 37214 31778 37266
rect 34302 37214 34354 37266
rect 37438 37214 37490 37266
rect 39790 37214 39842 37266
rect 42590 37214 42642 37266
rect 44382 37214 44434 37266
rect 46398 37214 46450 37266
rect 46846 37214 46898 37266
rect 47518 37214 47570 37266
rect 2382 37102 2434 37154
rect 3054 37102 3106 37154
rect 3502 37102 3554 37154
rect 5182 37102 5234 37154
rect 5630 37102 5682 37154
rect 6078 37102 6130 37154
rect 6526 37102 6578 37154
rect 7982 37102 8034 37154
rect 13694 37102 13746 37154
rect 14590 37102 14642 37154
rect 19406 37102 19458 37154
rect 27582 37102 27634 37154
rect 30158 37102 30210 37154
rect 30718 37102 30770 37154
rect 32174 37102 32226 37154
rect 32846 37102 32898 37154
rect 33518 37102 33570 37154
rect 34862 37102 34914 37154
rect 35982 37102 36034 37154
rect 39902 37102 39954 37154
rect 40574 37102 40626 37154
rect 42702 37102 42754 37154
rect 43374 37102 43426 37154
rect 44158 37102 44210 37154
rect 48302 37102 48354 37154
rect 56366 37102 56418 37154
rect 56702 37102 56754 37154
rect 4734 36990 4786 37042
rect 5294 36990 5346 37042
rect 6414 36990 6466 37042
rect 10222 36990 10274 37042
rect 11230 36990 11282 37042
rect 16382 36990 16434 37042
rect 16718 36990 16770 37042
rect 16830 36990 16882 37042
rect 19406 36990 19458 37042
rect 19966 36990 20018 37042
rect 20526 36990 20578 37042
rect 24110 36990 24162 37042
rect 24894 36990 24946 37042
rect 55918 36990 55970 37042
rect 56366 36990 56418 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 1822 36654 1874 36706
rect 2382 36654 2434 36706
rect 9998 36654 10050 36706
rect 16718 36654 16770 36706
rect 17390 36654 17442 36706
rect 19406 36654 19458 36706
rect 20190 36654 20242 36706
rect 20526 36654 20578 36706
rect 23662 36654 23714 36706
rect 24334 36654 24386 36706
rect 28366 36654 28418 36706
rect 31054 36654 31106 36706
rect 1822 36542 1874 36594
rect 6190 36542 6242 36594
rect 7870 36542 7922 36594
rect 10894 36542 10946 36594
rect 12126 36542 12178 36594
rect 17838 36542 17890 36594
rect 23662 36542 23714 36594
rect 30046 36542 30098 36594
rect 42926 36654 42978 36706
rect 43262 36654 43314 36706
rect 43934 36654 43986 36706
rect 46286 36654 46338 36706
rect 31502 36542 31554 36594
rect 31950 36542 32002 36594
rect 32958 36542 33010 36594
rect 33966 36542 34018 36594
rect 34526 36542 34578 36594
rect 35870 36542 35922 36594
rect 36430 36542 36482 36594
rect 38782 36542 38834 36594
rect 41694 36542 41746 36594
rect 43822 36542 43874 36594
rect 46510 36542 46562 36594
rect 47854 36542 47906 36594
rect 50654 36542 50706 36594
rect 53902 36542 53954 36594
rect 55022 36542 55074 36594
rect 57486 36542 57538 36594
rect 57822 36542 57874 36594
rect 2830 36430 2882 36482
rect 4062 36430 4114 36482
rect 4510 36430 4562 36482
rect 5966 36430 6018 36482
rect 6526 36430 6578 36482
rect 7534 36430 7586 36482
rect 7982 36430 8034 36482
rect 8766 36430 8818 36482
rect 9326 36430 9378 36482
rect 9438 36430 9490 36482
rect 10110 36430 10162 36482
rect 11566 36430 11618 36482
rect 13918 36430 13970 36482
rect 14590 36430 14642 36482
rect 15486 36430 15538 36482
rect 17614 36430 17666 36482
rect 18174 36430 18226 36482
rect 18286 36430 18338 36482
rect 18958 36430 19010 36482
rect 19182 36430 19234 36482
rect 21534 36430 21586 36482
rect 21870 36430 21922 36482
rect 22766 36430 22818 36482
rect 25342 36430 25394 36482
rect 25902 36430 25954 36482
rect 26126 36430 26178 36482
rect 26574 36430 26626 36482
rect 28478 36430 28530 36482
rect 29486 36430 29538 36482
rect 29934 36430 29986 36482
rect 31838 36430 31890 36482
rect 33406 36430 33458 36482
rect 33854 36430 33906 36482
rect 35310 36430 35362 36482
rect 37886 36430 37938 36482
rect 39678 36430 39730 36482
rect 40014 36430 40066 36482
rect 41134 36430 41186 36482
rect 41358 36430 41410 36482
rect 47070 36430 47122 36482
rect 47406 36430 47458 36482
rect 50878 36430 50930 36482
rect 53342 36430 53394 36482
rect 57374 36430 57426 36482
rect 3950 36318 4002 36370
rect 4846 36318 4898 36370
rect 6414 36318 6466 36370
rect 7646 36318 7698 36370
rect 10670 36318 10722 36370
rect 10894 36318 10946 36370
rect 13806 36318 13858 36370
rect 14478 36318 14530 36370
rect 16718 36318 16770 36370
rect 16830 36318 16882 36370
rect 19966 36318 20018 36370
rect 22206 36318 22258 36370
rect 25006 36318 25058 36370
rect 26014 36318 26066 36370
rect 28814 36318 28866 36370
rect 30158 36318 30210 36370
rect 31614 36318 31666 36370
rect 32062 36318 32114 36370
rect 34078 36318 34130 36370
rect 39790 36318 39842 36370
rect 42702 36318 42754 36370
rect 50206 36318 50258 36370
rect 50430 36318 50482 36370
rect 54574 36318 54626 36370
rect 54798 36318 54850 36370
rect 55134 36318 55186 36370
rect 2270 36206 2322 36258
rect 3838 36206 3890 36258
rect 9214 36206 9266 36258
rect 10446 36206 10498 36258
rect 12910 36206 12962 36258
rect 14814 36206 14866 36258
rect 18062 36206 18114 36258
rect 19070 36206 19122 36258
rect 20414 36206 20466 36258
rect 20862 36206 20914 36258
rect 21758 36206 21810 36258
rect 22878 36206 22930 36258
rect 23102 36206 23154 36258
rect 23998 36206 24050 36258
rect 24446 36206 24498 36258
rect 25118 36206 25170 36258
rect 31054 36206 31106 36258
rect 32622 36206 32674 36258
rect 35758 36206 35810 36258
rect 35982 36206 36034 36258
rect 37438 36206 37490 36258
rect 38334 36206 38386 36258
rect 40462 36206 40514 36258
rect 42254 36206 42306 36258
rect 44382 36206 44434 36258
rect 45502 36206 45554 36258
rect 46510 36206 46562 36258
rect 47294 36206 47346 36258
rect 51214 36206 51266 36258
rect 53790 36206 53842 36258
rect 54014 36206 54066 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 7198 35870 7250 35922
rect 8542 35870 8594 35922
rect 8990 35870 9042 35922
rect 10894 35870 10946 35922
rect 11790 35870 11842 35922
rect 13022 35870 13074 35922
rect 13470 35870 13522 35922
rect 14254 35870 14306 35922
rect 15038 35870 15090 35922
rect 16942 35870 16994 35922
rect 18622 35870 18674 35922
rect 19406 35870 19458 35922
rect 20302 35870 20354 35922
rect 22206 35870 22258 35922
rect 26014 35870 26066 35922
rect 26126 35870 26178 35922
rect 26798 35870 26850 35922
rect 33854 35870 33906 35922
rect 34974 35870 35026 35922
rect 38558 35870 38610 35922
rect 39678 35870 39730 35922
rect 44494 35870 44546 35922
rect 45502 35870 45554 35922
rect 46734 35870 46786 35922
rect 49758 35870 49810 35922
rect 51998 35870 52050 35922
rect 57710 35870 57762 35922
rect 5518 35758 5570 35810
rect 13694 35758 13746 35810
rect 15150 35758 15202 35810
rect 16046 35758 16098 35810
rect 16270 35758 16322 35810
rect 17726 35758 17778 35810
rect 20078 35758 20130 35810
rect 30830 35758 30882 35810
rect 40686 35758 40738 35810
rect 43486 35758 43538 35810
rect 44942 35758 44994 35810
rect 45390 35758 45442 35810
rect 53902 35758 53954 35810
rect 56590 35758 56642 35810
rect 57486 35758 57538 35810
rect 3390 35646 3442 35698
rect 4174 35646 4226 35698
rect 4734 35646 4786 35698
rect 5406 35646 5458 35698
rect 5742 35646 5794 35698
rect 6750 35646 6802 35698
rect 10110 35646 10162 35698
rect 10558 35646 10610 35698
rect 10782 35646 10834 35698
rect 11006 35646 11058 35698
rect 11902 35646 11954 35698
rect 12350 35646 12402 35698
rect 13806 35646 13858 35698
rect 14926 35646 14978 35698
rect 16606 35646 16658 35698
rect 16830 35646 16882 35698
rect 17950 35646 18002 35698
rect 18286 35646 18338 35698
rect 20526 35646 20578 35698
rect 21086 35646 21138 35698
rect 21310 35646 21362 35698
rect 21758 35646 21810 35698
rect 23326 35646 23378 35698
rect 23886 35646 23938 35698
rect 25790 35646 25842 35698
rect 25902 35646 25954 35698
rect 26350 35646 26402 35698
rect 27470 35646 27522 35698
rect 27806 35646 27858 35698
rect 29486 35646 29538 35698
rect 30270 35646 30322 35698
rect 31614 35646 31666 35698
rect 31838 35646 31890 35698
rect 32174 35646 32226 35698
rect 34638 35646 34690 35698
rect 34862 35646 34914 35698
rect 35086 35646 35138 35698
rect 35310 35646 35362 35698
rect 36878 35646 36930 35698
rect 37326 35646 37378 35698
rect 37550 35646 37602 35698
rect 39902 35646 39954 35698
rect 41806 35646 41858 35698
rect 42030 35646 42082 35698
rect 45726 35646 45778 35698
rect 49534 35646 49586 35698
rect 51102 35646 51154 35698
rect 53006 35646 53058 35698
rect 53230 35646 53282 35698
rect 54798 35646 54850 35698
rect 55582 35646 55634 35698
rect 57710 35646 57762 35698
rect 57934 35646 57986 35698
rect 2158 35534 2210 35586
rect 2606 35534 2658 35586
rect 3502 35534 3554 35586
rect 6302 35534 6354 35586
rect 7646 35534 7698 35586
rect 8206 35534 8258 35586
rect 20414 35534 20466 35586
rect 21534 35534 21586 35586
rect 22654 35534 22706 35586
rect 24782 35534 24834 35586
rect 28926 35534 28978 35586
rect 30382 35534 30434 35586
rect 31950 35534 32002 35586
rect 32510 35534 32562 35586
rect 33966 35534 34018 35586
rect 35758 35534 35810 35586
rect 36206 35534 36258 35586
rect 37102 35534 37154 35586
rect 37438 35534 37490 35586
rect 38110 35534 38162 35586
rect 39118 35534 39170 35586
rect 40798 35534 40850 35586
rect 41582 35534 41634 35586
rect 43038 35534 43090 35586
rect 44046 35534 44098 35586
rect 46174 35534 46226 35586
rect 47742 35534 47794 35586
rect 48190 35534 48242 35586
rect 50766 35534 50818 35586
rect 51550 35534 51602 35586
rect 54686 35534 54738 35586
rect 56702 35534 56754 35586
rect 3726 35422 3778 35474
rect 7870 35422 7922 35474
rect 8206 35422 8258 35474
rect 10334 35422 10386 35474
rect 18510 35422 18562 35474
rect 33630 35422 33682 35474
rect 39566 35422 39618 35474
rect 40462 35422 40514 35474
rect 49870 35422 49922 35474
rect 56366 35422 56418 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 15150 35086 15202 35138
rect 15710 35086 15762 35138
rect 16830 35086 16882 35138
rect 20974 35086 21026 35138
rect 22654 35086 22706 35138
rect 23886 35086 23938 35138
rect 28254 35086 28306 35138
rect 41694 35086 41746 35138
rect 1822 34974 1874 35026
rect 2382 34974 2434 35026
rect 4398 34974 4450 35026
rect 7198 34974 7250 35026
rect 9662 34974 9714 35026
rect 12126 34974 12178 35026
rect 14254 34974 14306 35026
rect 15486 34974 15538 35026
rect 16046 34974 16098 35026
rect 17502 34974 17554 35026
rect 18398 34974 18450 35026
rect 20526 34974 20578 35026
rect 21534 34974 21586 35026
rect 22654 34974 22706 35026
rect 27022 34974 27074 35026
rect 28030 34974 28082 35026
rect 30382 34974 30434 35026
rect 37998 34974 38050 35026
rect 3390 34862 3442 34914
rect 3502 34862 3554 34914
rect 6862 34862 6914 34914
rect 7310 34862 7362 34914
rect 10558 34862 10610 34914
rect 11006 34862 11058 34914
rect 11902 34862 11954 34914
rect 13918 34862 13970 34914
rect 16494 34862 16546 34914
rect 18958 34862 19010 34914
rect 20078 34862 20130 34914
rect 20302 34862 20354 34914
rect 24222 34862 24274 34914
rect 24558 34862 24610 34914
rect 27470 34862 27522 34914
rect 30046 34862 30098 34914
rect 30270 34862 30322 34914
rect 3838 34750 3890 34802
rect 4062 34750 4114 34802
rect 4286 34750 4338 34802
rect 6190 34750 6242 34802
rect 7982 34750 8034 34802
rect 8318 34750 8370 34802
rect 8430 34750 8482 34802
rect 10334 34750 10386 34802
rect 14478 34750 14530 34802
rect 19182 34750 19234 34802
rect 25678 34750 25730 34802
rect 29710 34750 29762 34802
rect 40798 34974 40850 35026
rect 42030 34974 42082 35026
rect 45614 34974 45666 35026
rect 47518 34974 47570 35026
rect 50542 34974 50594 35026
rect 51774 34974 51826 35026
rect 54462 34974 54514 35026
rect 56478 34974 56530 35026
rect 57374 34974 57426 35026
rect 30830 34862 30882 34914
rect 31054 34862 31106 34914
rect 31166 34862 31218 34914
rect 32174 34862 32226 34914
rect 32398 34862 32450 34914
rect 32846 34862 32898 34914
rect 33182 34862 33234 34914
rect 34526 34862 34578 34914
rect 34974 34862 35026 34914
rect 35870 34862 35922 34914
rect 37550 34862 37602 34914
rect 37886 34862 37938 34914
rect 38222 34862 38274 34914
rect 42590 34862 42642 34914
rect 43262 34862 43314 34914
rect 43598 34862 43650 34914
rect 43934 34862 43986 34914
rect 45838 34862 45890 34914
rect 46958 34862 47010 34914
rect 49086 34862 49138 34914
rect 49870 34862 49922 34914
rect 51662 34862 51714 34914
rect 52558 34862 52610 34914
rect 53566 34862 53618 34914
rect 53790 34862 53842 34914
rect 56702 34862 56754 34914
rect 30718 34750 30770 34802
rect 33518 34750 33570 34802
rect 35086 34750 35138 34802
rect 36094 34750 36146 34802
rect 36206 34750 36258 34802
rect 38782 34750 38834 34802
rect 39006 34750 39058 34802
rect 42702 34750 42754 34802
rect 46510 34750 46562 34802
rect 48974 34750 49026 34802
rect 2830 34638 2882 34690
rect 5070 34638 5122 34690
rect 5966 34638 6018 34690
rect 6078 34638 6130 34690
rect 6974 34638 7026 34690
rect 7198 34638 7250 34690
rect 8094 34638 8146 34690
rect 8206 34638 8258 34690
rect 11118 34638 11170 34690
rect 12350 34638 12402 34690
rect 12462 34638 12514 34690
rect 12574 34638 12626 34690
rect 15150 34638 15202 34690
rect 16718 34638 16770 34690
rect 17950 34638 18002 34690
rect 19070 34638 19122 34690
rect 19406 34638 19458 34690
rect 21982 34638 22034 34690
rect 23102 34638 23154 34690
rect 23550 34638 23602 34690
rect 26350 34638 26402 34690
rect 28590 34638 28642 34690
rect 29934 34638 29986 34690
rect 31614 34638 31666 34690
rect 32286 34638 32338 34690
rect 33406 34638 33458 34690
rect 34190 34638 34242 34690
rect 36766 34638 36818 34690
rect 38894 34638 38946 34690
rect 39566 34638 39618 34690
rect 39902 34638 39954 34690
rect 40462 34638 40514 34690
rect 41918 34638 41970 34690
rect 42814 34638 42866 34690
rect 43822 34638 43874 34690
rect 44382 34638 44434 34690
rect 47406 34638 47458 34690
rect 47630 34638 47682 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 4174 34302 4226 34354
rect 4510 34302 4562 34354
rect 5406 34302 5458 34354
rect 8542 34302 8594 34354
rect 11902 34302 11954 34354
rect 12238 34302 12290 34354
rect 19182 34302 19234 34354
rect 23550 34302 23602 34354
rect 23998 34302 24050 34354
rect 24446 34302 24498 34354
rect 26014 34302 26066 34354
rect 29822 34302 29874 34354
rect 30606 34302 30658 34354
rect 36654 34302 36706 34354
rect 44942 34302 44994 34354
rect 51214 34302 51266 34354
rect 52110 34302 52162 34354
rect 52334 34302 52386 34354
rect 52670 34302 52722 34354
rect 54014 34302 54066 34354
rect 56366 34302 56418 34354
rect 2942 34190 2994 34242
rect 5294 34190 5346 34242
rect 5966 34190 6018 34242
rect 7310 34190 7362 34242
rect 7534 34190 7586 34242
rect 8206 34190 8258 34242
rect 12798 34190 12850 34242
rect 14142 34190 14194 34242
rect 15598 34190 15650 34242
rect 17838 34190 17890 34242
rect 17950 34190 18002 34242
rect 26462 34190 26514 34242
rect 35310 34190 35362 34242
rect 39230 34190 39282 34242
rect 39902 34190 39954 34242
rect 40798 34190 40850 34242
rect 42590 34190 42642 34242
rect 46958 34190 47010 34242
rect 49534 34190 49586 34242
rect 51998 34190 52050 34242
rect 57486 34190 57538 34242
rect 3502 34078 3554 34130
rect 4062 34078 4114 34130
rect 4286 34078 4338 34130
rect 6414 34078 6466 34130
rect 8094 34078 8146 34130
rect 10110 34078 10162 34130
rect 10782 34078 10834 34130
rect 13022 34078 13074 34130
rect 13694 34078 13746 34130
rect 14366 34078 14418 34130
rect 14814 34078 14866 34130
rect 15822 34078 15874 34130
rect 16046 34078 16098 34130
rect 16158 34078 16210 34130
rect 17614 34078 17666 34130
rect 21086 34078 21138 34130
rect 21534 34078 21586 34130
rect 21646 34078 21698 34130
rect 28590 34078 28642 34130
rect 31726 34078 31778 34130
rect 31950 34078 32002 34130
rect 34414 34078 34466 34130
rect 34638 34078 34690 34130
rect 35758 34078 35810 34130
rect 38110 34078 38162 34130
rect 39454 34078 39506 34130
rect 40014 34078 40066 34130
rect 41470 34078 41522 34130
rect 43934 34078 43986 34130
rect 46062 34078 46114 34130
rect 47854 34078 47906 34130
rect 49758 34078 49810 34130
rect 49982 34078 50034 34130
rect 53454 34078 53506 34130
rect 53678 34078 53730 34130
rect 55918 34078 55970 34130
rect 56142 34078 56194 34130
rect 56478 34078 56530 34130
rect 57934 34078 57986 34130
rect 1934 33966 1986 34018
rect 2494 33966 2546 34018
rect 8990 33966 9042 34018
rect 10558 33966 10610 34018
rect 15934 33966 15986 34018
rect 16942 33966 16994 34018
rect 18734 33966 18786 34018
rect 19742 33966 19794 34018
rect 20190 33966 20242 34018
rect 20638 33966 20690 34018
rect 21310 33966 21362 34018
rect 22318 33966 22370 34018
rect 22654 33966 22706 34018
rect 23102 33966 23154 34018
rect 24894 33966 24946 34018
rect 25566 33966 25618 34018
rect 28030 33966 28082 34018
rect 29038 33966 29090 34018
rect 32062 33966 32114 34018
rect 33518 33966 33570 34018
rect 36206 33966 36258 34018
rect 37102 33966 37154 34018
rect 37550 33966 37602 34018
rect 40238 33966 40290 34018
rect 42366 33966 42418 34018
rect 44494 33966 44546 34018
rect 46510 33966 46562 34018
rect 47630 33966 47682 34018
rect 48526 33966 48578 34018
rect 58270 33966 58322 34018
rect 5518 33854 5570 33906
rect 5742 33854 5794 33906
rect 6190 33854 6242 33906
rect 10110 33854 10162 33906
rect 22318 33854 22370 33906
rect 22542 33854 22594 33906
rect 23326 33854 23378 33906
rect 23662 33854 23714 33906
rect 24558 33854 24610 33906
rect 27134 33854 27186 33906
rect 27246 33854 27298 33906
rect 27470 33854 27522 33906
rect 30382 33854 30434 33906
rect 30718 33854 30770 33906
rect 32510 33854 32562 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 9886 33518 9938 33570
rect 10782 33518 10834 33570
rect 34750 33518 34802 33570
rect 35198 33518 35250 33570
rect 39118 33518 39170 33570
rect 42478 33518 42530 33570
rect 43374 33518 43426 33570
rect 48974 33518 49026 33570
rect 49534 33518 49586 33570
rect 2270 33406 2322 33458
rect 6078 33406 6130 33458
rect 6638 33406 6690 33458
rect 8094 33406 8146 33458
rect 12910 33406 12962 33458
rect 14254 33406 14306 33458
rect 14814 33406 14866 33458
rect 16046 33406 16098 33458
rect 19630 33406 19682 33458
rect 20414 33406 20466 33458
rect 22430 33406 22482 33458
rect 26798 33406 26850 33458
rect 27694 33406 27746 33458
rect 29822 33406 29874 33458
rect 32958 33406 33010 33458
rect 34302 33406 34354 33458
rect 35198 33406 35250 33458
rect 42478 33406 42530 33458
rect 43374 33406 43426 33458
rect 45502 33406 45554 33458
rect 56478 33406 56530 33458
rect 57934 33406 57986 33458
rect 3390 33294 3442 33346
rect 5630 33294 5682 33346
rect 6414 33294 6466 33346
rect 9998 33294 10050 33346
rect 14366 33294 14418 33346
rect 15038 33294 15090 33346
rect 15822 33294 15874 33346
rect 16270 33294 16322 33346
rect 17838 33294 17890 33346
rect 17950 33294 18002 33346
rect 18398 33294 18450 33346
rect 18846 33294 18898 33346
rect 18958 33294 19010 33346
rect 19966 33294 20018 33346
rect 21646 33294 21698 33346
rect 22878 33294 22930 33346
rect 23214 33294 23266 33346
rect 24222 33294 24274 33346
rect 24558 33294 24610 33346
rect 27582 33294 27634 33346
rect 28478 33294 28530 33346
rect 31166 33294 31218 33346
rect 32062 33294 32114 33346
rect 35982 33294 36034 33346
rect 37438 33294 37490 33346
rect 38446 33294 38498 33346
rect 41246 33294 41298 33346
rect 46398 33294 46450 33346
rect 46734 33294 46786 33346
rect 56254 33294 56306 33346
rect 57486 33294 57538 33346
rect 58046 33294 58098 33346
rect 4286 33182 4338 33234
rect 11790 33182 11842 33234
rect 17390 33182 17442 33234
rect 17614 33182 17666 33234
rect 18622 33182 18674 33234
rect 21982 33182 22034 33234
rect 22094 33182 22146 33234
rect 25790 33182 25842 33234
rect 27918 33182 27970 33234
rect 30718 33182 30770 33234
rect 32510 33182 32562 33234
rect 34750 33182 34802 33234
rect 36318 33182 36370 33234
rect 40014 33182 40066 33234
rect 40910 33182 40962 33234
rect 56926 33182 56978 33234
rect 2830 33070 2882 33122
rect 8542 33070 8594 33122
rect 9214 33070 9266 33122
rect 9886 33070 9938 33122
rect 12462 33070 12514 33122
rect 16382 33070 16434 33122
rect 16494 33070 16546 33122
rect 17726 33070 17778 33122
rect 19742 33070 19794 33122
rect 20862 33070 20914 33122
rect 21870 33070 21922 33122
rect 23102 33070 23154 33122
rect 26350 33070 26402 33122
rect 33406 33070 33458 33122
rect 33854 33070 33906 33122
rect 36430 33070 36482 33122
rect 36542 33070 36594 33122
rect 40126 33070 40178 33122
rect 40238 33070 40290 33122
rect 41022 33070 41074 33122
rect 41582 33070 41634 33122
rect 42030 33070 42082 33122
rect 43038 33070 43090 33122
rect 43822 33070 43874 33122
rect 44382 33070 44434 33122
rect 46510 33070 46562 33122
rect 47070 33070 47122 33122
rect 48974 33070 49026 33122
rect 49422 33070 49474 33122
rect 54798 33070 54850 33122
rect 57822 33070 57874 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 1934 32734 1986 32786
rect 2382 32734 2434 32786
rect 5518 32734 5570 32786
rect 6414 32734 6466 32786
rect 13806 32734 13858 32786
rect 15822 32734 15874 32786
rect 18398 32734 18450 32786
rect 19406 32734 19458 32786
rect 22990 32734 23042 32786
rect 31502 32734 31554 32786
rect 31726 32734 31778 32786
rect 32398 32734 32450 32786
rect 34526 32734 34578 32786
rect 39118 32734 39170 32786
rect 44046 32734 44098 32786
rect 49870 32734 49922 32786
rect 50878 32734 50930 32786
rect 57486 32734 57538 32786
rect 4286 32622 4338 32674
rect 6078 32622 6130 32674
rect 6190 32622 6242 32674
rect 8542 32622 8594 32674
rect 12126 32622 12178 32674
rect 13470 32622 13522 32674
rect 13582 32622 13634 32674
rect 14366 32622 14418 32674
rect 14590 32622 14642 32674
rect 16382 32622 16434 32674
rect 20302 32622 20354 32674
rect 20750 32622 20802 32674
rect 22766 32622 22818 32674
rect 23326 32622 23378 32674
rect 25678 32622 25730 32674
rect 30830 32622 30882 32674
rect 31838 32622 31890 32674
rect 35422 32622 35474 32674
rect 38334 32622 38386 32674
rect 44830 32622 44882 32674
rect 44942 32622 44994 32674
rect 54462 32622 54514 32674
rect 56030 32622 56082 32674
rect 57710 32622 57762 32674
rect 4510 32510 4562 32562
rect 5070 32510 5122 32562
rect 7422 32510 7474 32562
rect 7646 32510 7698 32562
rect 9102 32510 9154 32562
rect 10222 32510 10274 32562
rect 11230 32510 11282 32562
rect 11678 32510 11730 32562
rect 12574 32510 12626 32562
rect 14254 32510 14306 32562
rect 14702 32510 14754 32562
rect 16718 32510 16770 32562
rect 16942 32510 16994 32562
rect 18622 32510 18674 32562
rect 20190 32510 20242 32562
rect 21086 32510 21138 32562
rect 21758 32510 21810 32562
rect 23214 32510 23266 32562
rect 24334 32510 24386 32562
rect 26014 32510 26066 32562
rect 26910 32510 26962 32562
rect 28142 32510 28194 32562
rect 28702 32510 28754 32562
rect 29934 32510 29986 32562
rect 30494 32510 30546 32562
rect 34414 32510 34466 32562
rect 34750 32510 34802 32562
rect 35310 32510 35362 32562
rect 36990 32510 37042 32562
rect 38222 32510 38274 32562
rect 38558 32510 38610 32562
rect 39230 32510 39282 32562
rect 39902 32510 39954 32562
rect 40126 32510 40178 32562
rect 41918 32510 41970 32562
rect 42926 32510 42978 32562
rect 45166 32510 45218 32562
rect 50430 32510 50482 32562
rect 50766 32510 50818 32562
rect 50990 32510 51042 32562
rect 53790 32510 53842 32562
rect 55358 32510 55410 32562
rect 57822 32510 57874 32562
rect 2942 32398 2994 32450
rect 3390 32398 3442 32450
rect 4062 32398 4114 32450
rect 8094 32398 8146 32450
rect 9998 32398 10050 32450
rect 12350 32398 12402 32450
rect 15374 32398 15426 32450
rect 16494 32398 16546 32450
rect 17950 32398 18002 32450
rect 18174 32398 18226 32450
rect 18510 32398 18562 32450
rect 19966 32398 20018 32450
rect 23326 32398 23378 32450
rect 24110 32398 24162 32450
rect 25902 32398 25954 32450
rect 27918 32398 27970 32450
rect 32734 32398 32786 32450
rect 33630 32398 33682 32450
rect 37438 32398 37490 32450
rect 40798 32398 40850 32450
rect 42702 32398 42754 32450
rect 43598 32398 43650 32450
rect 45502 32398 45554 32450
rect 51550 32398 51602 32450
rect 54014 32398 54066 32450
rect 55134 32398 55186 32450
rect 6974 32286 7026 32338
rect 10110 32286 10162 32338
rect 17726 32286 17778 32338
rect 24558 32286 24610 32338
rect 25006 32286 25058 32338
rect 27582 32286 27634 32338
rect 36094 32286 36146 32338
rect 36430 32286 36482 32338
rect 39118 32286 39170 32338
rect 42030 32286 42082 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 2046 31950 2098 32002
rect 2494 31950 2546 32002
rect 18510 31950 18562 32002
rect 19294 31950 19346 32002
rect 28142 31950 28194 32002
rect 28478 31950 28530 32002
rect 58158 31950 58210 32002
rect 2382 31838 2434 31890
rect 3390 31838 3442 31890
rect 5070 31838 5122 31890
rect 5854 31838 5906 31890
rect 6302 31838 6354 31890
rect 12910 31838 12962 31890
rect 16830 31838 16882 31890
rect 17726 31838 17778 31890
rect 18286 31838 18338 31890
rect 19070 31838 19122 31890
rect 20190 31838 20242 31890
rect 22878 31838 22930 31890
rect 23550 31838 23602 31890
rect 24446 31838 24498 31890
rect 25006 31838 25058 31890
rect 26574 31838 26626 31890
rect 27918 31838 27970 31890
rect 34190 31838 34242 31890
rect 40014 31838 40066 31890
rect 44382 31838 44434 31890
rect 47070 31838 47122 31890
rect 48302 31838 48354 31890
rect 53902 31838 53954 31890
rect 54462 31838 54514 31890
rect 55470 31838 55522 31890
rect 55806 31838 55858 31890
rect 57710 31838 57762 31890
rect 6750 31726 6802 31778
rect 7086 31726 7138 31778
rect 7758 31726 7810 31778
rect 7870 31726 7922 31778
rect 9326 31726 9378 31778
rect 11118 31726 11170 31778
rect 13582 31726 13634 31778
rect 13918 31726 13970 31778
rect 15150 31726 15202 31778
rect 15822 31726 15874 31778
rect 18734 31726 18786 31778
rect 19966 31726 20018 31778
rect 20526 31726 20578 31778
rect 21758 31726 21810 31778
rect 21982 31726 22034 31778
rect 22430 31726 22482 31778
rect 23774 31726 23826 31778
rect 25902 31726 25954 31778
rect 26686 31726 26738 31778
rect 29934 31726 29986 31778
rect 31838 31726 31890 31778
rect 32622 31726 32674 31778
rect 34078 31726 34130 31778
rect 34414 31726 34466 31778
rect 36430 31726 36482 31778
rect 39230 31726 39282 31778
rect 41694 31726 41746 31778
rect 42254 31726 42306 31778
rect 43822 31726 43874 31778
rect 45390 31726 45442 31778
rect 46062 31726 46114 31778
rect 48414 31726 48466 31778
rect 49758 31726 49810 31778
rect 49982 31726 50034 31778
rect 51774 31726 51826 31778
rect 52446 31726 52498 31778
rect 53342 31726 53394 31778
rect 55246 31726 55298 31778
rect 57598 31726 57650 31778
rect 2830 31614 2882 31666
rect 8654 31614 8706 31666
rect 9214 31614 9266 31666
rect 11454 31614 11506 31666
rect 14142 31614 14194 31666
rect 14590 31614 14642 31666
rect 15262 31614 15314 31666
rect 15486 31614 15538 31666
rect 20414 31614 20466 31666
rect 27358 31614 27410 31666
rect 29598 31614 29650 31666
rect 31726 31614 31778 31666
rect 35870 31614 35922 31666
rect 37774 31614 37826 31666
rect 38894 31614 38946 31666
rect 42814 31614 42866 31666
rect 44718 31614 44770 31666
rect 45838 31614 45890 31666
rect 49086 31614 49138 31666
rect 50654 31614 50706 31666
rect 52670 31614 52722 31666
rect 54014 31614 54066 31666
rect 1934 31502 1986 31554
rect 3838 31502 3890 31554
rect 4622 31502 4674 31554
rect 7646 31502 7698 31554
rect 8094 31502 8146 31554
rect 12014 31502 12066 31554
rect 12462 31502 12514 31554
rect 14254 31502 14306 31554
rect 16158 31502 16210 31554
rect 17278 31502 17330 31554
rect 19518 31502 19570 31554
rect 22206 31502 22258 31554
rect 25566 31502 25618 31554
rect 28366 31502 28418 31554
rect 28814 31502 28866 31554
rect 30158 31502 30210 31554
rect 30718 31502 30770 31554
rect 31166 31502 31218 31554
rect 31950 31502 32002 31554
rect 37438 31502 37490 31554
rect 37662 31502 37714 31554
rect 42926 31502 42978 31554
rect 43150 31502 43202 31554
rect 45950 31502 46002 31554
rect 47518 31502 47570 31554
rect 53790 31502 53842 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 2382 31166 2434 31218
rect 2718 31166 2770 31218
rect 12126 31166 12178 31218
rect 12686 31166 12738 31218
rect 13134 31166 13186 31218
rect 13694 31166 13746 31218
rect 17054 31166 17106 31218
rect 17838 31166 17890 31218
rect 18846 31166 18898 31218
rect 21422 31166 21474 31218
rect 21646 31166 21698 31218
rect 23998 31166 24050 31218
rect 25006 31166 25058 31218
rect 35310 31166 35362 31218
rect 35982 31166 36034 31218
rect 38110 31166 38162 31218
rect 40574 31166 40626 31218
rect 43822 31166 43874 31218
rect 44270 31166 44322 31218
rect 44718 31166 44770 31218
rect 47182 31166 47234 31218
rect 47630 31166 47682 31218
rect 48750 31166 48802 31218
rect 52782 31166 52834 31218
rect 54798 31166 54850 31218
rect 55246 31166 55298 31218
rect 7198 31054 7250 31106
rect 16494 31054 16546 31106
rect 19406 31054 19458 31106
rect 21870 31054 21922 31106
rect 29374 31054 29426 31106
rect 32622 31054 32674 31106
rect 32734 31054 32786 31106
rect 33742 31054 33794 31106
rect 35646 31054 35698 31106
rect 39118 31054 39170 31106
rect 39790 31054 39842 31106
rect 40014 31054 40066 31106
rect 42702 31054 42754 31106
rect 48190 31054 48242 31106
rect 49534 31054 49586 31106
rect 49758 31054 49810 31106
rect 51550 31054 51602 31106
rect 52446 31054 52498 31106
rect 52558 31054 52610 31106
rect 3726 30942 3778 30994
rect 4846 30942 4898 30994
rect 5182 30942 5234 30994
rect 6638 30942 6690 30994
rect 7086 30942 7138 30994
rect 8542 30942 8594 30994
rect 8766 30942 8818 30994
rect 8990 30942 9042 30994
rect 9662 30942 9714 30994
rect 10110 30942 10162 30994
rect 10334 30942 10386 30994
rect 10782 30942 10834 30994
rect 11230 30942 11282 30994
rect 11454 30942 11506 30994
rect 13806 30942 13858 30994
rect 15150 30942 15202 30994
rect 15374 30942 15426 30994
rect 19294 30942 19346 30994
rect 20302 30942 20354 30994
rect 25902 30942 25954 30994
rect 26126 30942 26178 30994
rect 27582 30942 27634 30994
rect 28478 30942 28530 30994
rect 31838 30942 31890 30994
rect 34190 30942 34242 30994
rect 34638 30942 34690 30994
rect 34974 30942 35026 30994
rect 36766 30942 36818 30994
rect 36990 30942 37042 30994
rect 41806 30942 41858 30994
rect 43150 30942 43202 30994
rect 43598 30942 43650 30994
rect 45838 30942 45890 30994
rect 50878 30942 50930 30994
rect 1934 30830 1986 30882
rect 7310 30830 7362 30882
rect 8878 30830 8930 30882
rect 10222 30830 10274 30882
rect 11006 30830 11058 30882
rect 13918 30830 13970 30882
rect 18286 30830 18338 30882
rect 19854 30830 19906 30882
rect 20078 30830 20130 30882
rect 21534 30830 21586 30882
rect 22654 30830 22706 30882
rect 23214 30830 23266 30882
rect 23662 30830 23714 30882
rect 24446 30830 24498 30882
rect 25678 30830 25730 30882
rect 30494 30830 30546 30882
rect 37662 30830 37714 30882
rect 39230 30830 39282 30882
rect 39902 30830 39954 30882
rect 42142 30830 42194 30882
rect 43710 30830 43762 30882
rect 46062 30830 46114 30882
rect 49870 30830 49922 30882
rect 51102 30830 51154 30882
rect 53118 30830 53170 30882
rect 56366 30830 56418 30882
rect 56814 30830 56866 30882
rect 57486 30830 57538 30882
rect 3614 30718 3666 30770
rect 15710 30718 15762 30770
rect 17502 30718 17554 30770
rect 18174 30718 18226 30770
rect 26574 30718 26626 30770
rect 29822 30718 29874 30770
rect 30718 30718 30770 30770
rect 31054 30718 31106 30770
rect 32734 30718 32786 30770
rect 38894 30718 38946 30770
rect 44046 30718 44098 30770
rect 44382 30718 44434 30770
rect 46398 30718 46450 30770
rect 48414 30718 48466 30770
rect 57710 30718 57762 30770
rect 58046 30718 58098 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 6862 30382 6914 30434
rect 16830 30382 16882 30434
rect 19630 30382 19682 30434
rect 35534 30382 35586 30434
rect 37886 30382 37938 30434
rect 42030 30382 42082 30434
rect 43598 30382 43650 30434
rect 8430 30270 8482 30322
rect 9774 30270 9826 30322
rect 12014 30270 12066 30322
rect 12574 30270 12626 30322
rect 15262 30270 15314 30322
rect 16606 30270 16658 30322
rect 26014 30270 26066 30322
rect 28366 30270 28418 30322
rect 31726 30270 31778 30322
rect 44046 30270 44098 30322
rect 47406 30270 47458 30322
rect 48414 30270 48466 30322
rect 49870 30270 49922 30322
rect 56590 30270 56642 30322
rect 57374 30270 57426 30322
rect 3054 30158 3106 30210
rect 3278 30158 3330 30210
rect 4622 30158 4674 30210
rect 4958 30102 5010 30154
rect 7198 30158 7250 30210
rect 7982 30158 8034 30210
rect 9550 30158 9602 30210
rect 11006 30158 11058 30210
rect 11118 30158 11170 30210
rect 11902 30158 11954 30210
rect 13694 30158 13746 30210
rect 14366 30158 14418 30210
rect 16382 30158 16434 30210
rect 17278 30158 17330 30210
rect 18174 30158 18226 30210
rect 18398 30158 18450 30210
rect 19182 30158 19234 30210
rect 19406 30158 19458 30210
rect 19742 30158 19794 30210
rect 22654 30158 22706 30210
rect 22990 30158 23042 30210
rect 25230 30158 25282 30210
rect 25342 30158 25394 30210
rect 25902 30158 25954 30210
rect 26798 30158 26850 30210
rect 27806 30158 27858 30210
rect 30382 30158 30434 30210
rect 32398 30158 32450 30210
rect 33294 30158 33346 30210
rect 33630 30158 33682 30210
rect 34078 30158 34130 30210
rect 35870 30158 35922 30210
rect 36094 30158 36146 30210
rect 36206 30158 36258 30210
rect 36766 30158 36818 30210
rect 39454 30158 39506 30210
rect 42254 30158 42306 30210
rect 46398 30158 46450 30210
rect 46846 30158 46898 30210
rect 50094 30158 50146 30210
rect 52670 30158 52722 30210
rect 53678 30158 53730 30210
rect 54126 30158 54178 30210
rect 55470 30158 55522 30210
rect 55694 30158 55746 30210
rect 57262 30158 57314 30210
rect 2382 30046 2434 30098
rect 6302 30046 6354 30098
rect 6526 30046 6578 30098
rect 9214 30046 9266 30098
rect 11678 30046 11730 30098
rect 14142 30046 14194 30098
rect 17726 30046 17778 30098
rect 24222 30046 24274 30098
rect 25118 30046 25170 30098
rect 25678 30046 25730 30098
rect 27582 30046 27634 30098
rect 30718 30046 30770 30098
rect 37550 30046 37602 30098
rect 39230 30046 39282 30098
rect 40574 30046 40626 30098
rect 43486 30046 43538 30098
rect 48078 30046 48130 30098
rect 49198 30046 49250 30098
rect 50766 30046 50818 30098
rect 53454 30046 53506 30098
rect 58158 30046 58210 30098
rect 1822 29934 1874 29986
rect 4846 29934 4898 29986
rect 10446 29934 10498 29986
rect 11454 29934 11506 29986
rect 12910 29934 12962 29986
rect 17950 29934 18002 29986
rect 18062 29934 18114 29986
rect 19966 29934 20018 29986
rect 20414 29934 20466 29986
rect 20862 29934 20914 29986
rect 21534 29934 21586 29986
rect 22094 29934 22146 29986
rect 29598 29934 29650 29986
rect 35982 29934 36034 29986
rect 37774 29934 37826 29986
rect 40462 29934 40514 29986
rect 41246 29934 41298 29986
rect 41694 29934 41746 29986
rect 42590 29934 42642 29986
rect 43038 29934 43090 29986
rect 46062 29934 46114 29986
rect 47294 29934 47346 29986
rect 47518 29934 47570 29986
rect 48302 29934 48354 29986
rect 51214 29934 51266 29986
rect 53790 29934 53842 29986
rect 54910 29934 54962 29986
rect 56030 29934 56082 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 3502 29598 3554 29650
rect 4286 29598 4338 29650
rect 6078 29598 6130 29650
rect 9886 29598 9938 29650
rect 11342 29598 11394 29650
rect 12126 29598 12178 29650
rect 12686 29598 12738 29650
rect 14590 29598 14642 29650
rect 15262 29598 15314 29650
rect 19518 29598 19570 29650
rect 22430 29598 22482 29650
rect 25678 29598 25730 29650
rect 25790 29598 25842 29650
rect 25902 29598 25954 29650
rect 32062 29598 32114 29650
rect 32734 29598 32786 29650
rect 33854 29598 33906 29650
rect 34974 29598 35026 29650
rect 35870 29598 35922 29650
rect 36430 29598 36482 29650
rect 38894 29598 38946 29650
rect 45166 29598 45218 29650
rect 46286 29598 46338 29650
rect 46398 29598 46450 29650
rect 46958 29598 47010 29650
rect 47742 29598 47794 29650
rect 57822 29598 57874 29650
rect 2718 29486 2770 29538
rect 5294 29486 5346 29538
rect 8878 29486 8930 29538
rect 10782 29486 10834 29538
rect 11678 29486 11730 29538
rect 13246 29486 13298 29538
rect 14030 29486 14082 29538
rect 17950 29486 18002 29538
rect 18174 29486 18226 29538
rect 19294 29486 19346 29538
rect 20414 29486 20466 29538
rect 24558 29486 24610 29538
rect 27134 29486 27186 29538
rect 27246 29486 27298 29538
rect 29150 29486 29202 29538
rect 30382 29486 30434 29538
rect 32510 29486 32562 29538
rect 33630 29486 33682 29538
rect 44382 29486 44434 29538
rect 53006 29486 53058 29538
rect 57486 29486 57538 29538
rect 4622 29374 4674 29426
rect 5406 29374 5458 29426
rect 6750 29374 6802 29426
rect 7870 29374 7922 29426
rect 9774 29374 9826 29426
rect 11342 29374 11394 29426
rect 13806 29374 13858 29426
rect 14366 29374 14418 29426
rect 15150 29374 15202 29426
rect 16158 29374 16210 29426
rect 20302 29374 20354 29426
rect 21310 29374 21362 29426
rect 23438 29374 23490 29426
rect 26126 29374 26178 29426
rect 26462 29374 26514 29426
rect 26910 29374 26962 29426
rect 28142 29374 28194 29426
rect 28478 29374 28530 29426
rect 30830 29374 30882 29426
rect 31166 29374 31218 29426
rect 31950 29374 32002 29426
rect 34526 29374 34578 29426
rect 34750 29374 34802 29426
rect 35086 29374 35138 29426
rect 35758 29374 35810 29426
rect 36094 29374 36146 29426
rect 37774 29374 37826 29426
rect 39790 29374 39842 29426
rect 40014 29374 40066 29426
rect 40238 29374 40290 29426
rect 40462 29374 40514 29426
rect 40686 29374 40738 29426
rect 41694 29374 41746 29426
rect 41918 29374 41970 29426
rect 43486 29374 43538 29426
rect 52110 29374 52162 29426
rect 52446 29374 52498 29426
rect 53902 29374 53954 29426
rect 57710 29374 57762 29426
rect 58046 29374 58098 29426
rect 2718 29262 2770 29314
rect 8318 29262 8370 29314
rect 11006 29262 11058 29314
rect 16494 29262 16546 29314
rect 16942 29262 16994 29314
rect 18846 29262 18898 29314
rect 19630 29262 19682 29314
rect 20526 29262 20578 29314
rect 21086 29262 21138 29314
rect 23550 29262 23602 29314
rect 28590 29262 28642 29314
rect 29822 29262 29874 29314
rect 34862 29262 34914 29314
rect 37550 29262 37602 29314
rect 40574 29262 40626 29314
rect 42590 29262 42642 29314
rect 44046 29262 44098 29314
rect 45726 29262 45778 29314
rect 46174 29262 46226 29314
rect 54126 29262 54178 29314
rect 54574 29262 54626 29314
rect 55134 29262 55186 29314
rect 55358 29262 55410 29314
rect 56142 29262 56194 29314
rect 56702 29262 56754 29314
rect 9886 29150 9938 29202
rect 11230 29150 11282 29202
rect 14366 29150 14418 29202
rect 15262 29150 15314 29202
rect 18286 29150 18338 29202
rect 33966 29150 34018 29202
rect 38334 29150 38386 29202
rect 43150 29150 43202 29202
rect 43486 29150 43538 29202
rect 55694 29150 55746 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 3950 28814 4002 28866
rect 10334 28814 10386 28866
rect 18846 28814 18898 28866
rect 28030 28814 28082 28866
rect 34750 28814 34802 28866
rect 36430 28814 36482 28866
rect 36654 28814 36706 28866
rect 40014 28814 40066 28866
rect 48078 28814 48130 28866
rect 52334 28814 52386 28866
rect 52670 28814 52722 28866
rect 2046 28702 2098 28754
rect 3166 28702 3218 28754
rect 4510 28702 4562 28754
rect 5854 28702 5906 28754
rect 6414 28702 6466 28754
rect 10894 28702 10946 28754
rect 11790 28702 11842 28754
rect 13694 28702 13746 28754
rect 14926 28702 14978 28754
rect 16942 28702 16994 28754
rect 23550 28702 23602 28754
rect 24558 28702 24610 28754
rect 25230 28702 25282 28754
rect 25790 28702 25842 28754
rect 35870 28702 35922 28754
rect 36654 28702 36706 28754
rect 37438 28702 37490 28754
rect 37886 28702 37938 28754
rect 38334 28702 38386 28754
rect 38782 28702 38834 28754
rect 40350 28702 40402 28754
rect 40798 28702 40850 28754
rect 43934 28702 43986 28754
rect 45390 28702 45442 28754
rect 45838 28702 45890 28754
rect 46286 28702 46338 28754
rect 47070 28702 47122 28754
rect 49310 28702 49362 28754
rect 54350 28702 54402 28754
rect 55134 28702 55186 28754
rect 57822 28702 57874 28754
rect 3054 28590 3106 28642
rect 4958 28590 5010 28642
rect 8318 28590 8370 28642
rect 9102 28590 9154 28642
rect 9550 28590 9602 28642
rect 10670 28590 10722 28642
rect 12686 28590 12738 28642
rect 12910 28590 12962 28642
rect 14142 28590 14194 28642
rect 15374 28590 15426 28642
rect 17166 28590 17218 28642
rect 17502 28590 17554 28642
rect 19070 28590 19122 28642
rect 19294 28590 19346 28642
rect 20526 28590 20578 28642
rect 20974 28590 21026 28642
rect 21982 28590 22034 28642
rect 23662 28590 23714 28642
rect 26238 28590 26290 28642
rect 27694 28590 27746 28642
rect 27806 28590 27858 28642
rect 30158 28590 30210 28642
rect 31390 28590 31442 28642
rect 31614 28590 31666 28642
rect 32286 28590 32338 28642
rect 35086 28590 35138 28642
rect 35982 28590 36034 28642
rect 42926 28590 42978 28642
rect 43486 28590 43538 28642
rect 47182 28590 47234 28642
rect 48302 28590 48354 28642
rect 49870 28590 49922 28642
rect 50094 28590 50146 28642
rect 50430 28590 50482 28642
rect 52110 28590 52162 28642
rect 53342 28590 53394 28642
rect 55022 28590 55074 28642
rect 56366 28590 56418 28642
rect 57934 28590 57986 28642
rect 58270 28590 58322 28642
rect 7086 28478 7138 28530
rect 9662 28478 9714 28530
rect 12350 28478 12402 28530
rect 14478 28478 14530 28530
rect 14926 28478 14978 28530
rect 18622 28478 18674 28530
rect 22206 28478 22258 28530
rect 27022 28478 27074 28530
rect 28590 28478 28642 28530
rect 29934 28478 29986 28530
rect 30942 28478 30994 28530
rect 32846 28478 32898 28530
rect 34190 28478 34242 28530
rect 34526 28478 34578 28530
rect 36094 28478 36146 28530
rect 39454 28478 39506 28530
rect 39678 28478 39730 28530
rect 41582 28478 41634 28530
rect 41918 28478 41970 28530
rect 43710 28478 43762 28530
rect 44046 28478 44098 28530
rect 57150 28478 57202 28530
rect 57710 28478 57762 28530
rect 7982 28366 8034 28418
rect 9774 28366 9826 28418
rect 10782 28366 10834 28418
rect 11006 28366 11058 28418
rect 12574 28366 12626 28418
rect 17838 28366 17890 28418
rect 19742 28366 19794 28418
rect 30158 28366 30210 28418
rect 32510 28366 32562 28418
rect 33182 28366 33234 28418
rect 39902 28366 39954 28418
rect 41694 28366 41746 28418
rect 42366 28366 42418 28418
rect 44606 28366 44658 28418
rect 48638 28366 48690 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 5294 28030 5346 28082
rect 6078 28030 6130 28082
rect 13246 28030 13298 28082
rect 13806 28030 13858 28082
rect 14254 28030 14306 28082
rect 15710 28030 15762 28082
rect 16606 28030 16658 28082
rect 20862 28030 20914 28082
rect 22318 28030 22370 28082
rect 23214 28030 23266 28082
rect 23662 28030 23714 28082
rect 24110 28030 24162 28082
rect 25006 28030 25058 28082
rect 29374 28030 29426 28082
rect 32734 28030 32786 28082
rect 34190 28030 34242 28082
rect 38110 28030 38162 28082
rect 41918 28030 41970 28082
rect 4174 27918 4226 27970
rect 8990 27918 9042 27970
rect 14702 27918 14754 27970
rect 18510 27918 18562 27970
rect 25902 27918 25954 27970
rect 30270 27918 30322 27970
rect 31838 27918 31890 27970
rect 33630 27918 33682 27970
rect 36318 27918 36370 27970
rect 36990 27918 37042 27970
rect 37662 27918 37714 27970
rect 45614 27918 45666 27970
rect 47406 27918 47458 27970
rect 48638 27918 48690 27970
rect 49870 27918 49922 27970
rect 2494 27806 2546 27858
rect 3054 27806 3106 27858
rect 6974 27806 7026 27858
rect 8430 27806 8482 27858
rect 9774 27806 9826 27858
rect 9998 27806 10050 27858
rect 11902 27806 11954 27858
rect 15150 27806 15202 27858
rect 15598 27806 15650 27858
rect 19854 27806 19906 27858
rect 20302 27806 20354 27858
rect 22766 27806 22818 27858
rect 24558 27806 24610 27858
rect 27694 27806 27746 27858
rect 28030 27806 28082 27858
rect 29934 27806 29986 27858
rect 32174 27806 32226 27858
rect 35422 27806 35474 27858
rect 35646 27806 35698 27858
rect 37102 27806 37154 27858
rect 39566 27806 39618 27858
rect 43038 27806 43090 27858
rect 44158 27806 44210 27858
rect 45950 27806 46002 27858
rect 46510 27806 46562 27858
rect 51102 27806 51154 27858
rect 52670 27806 52722 27858
rect 1934 27694 1986 27746
rect 8094 27694 8146 27746
rect 17054 27694 17106 27746
rect 18062 27694 18114 27746
rect 18846 27694 18898 27746
rect 19966 27694 20018 27746
rect 21310 27694 21362 27746
rect 26014 27694 26066 27746
rect 26462 27694 26514 27746
rect 28590 27694 28642 27746
rect 39118 27694 39170 27746
rect 40014 27694 40066 27746
rect 40462 27694 40514 27746
rect 41470 27694 41522 27746
rect 43150 27694 43202 27746
rect 44942 27694 44994 27746
rect 48190 27694 48242 27746
rect 49646 27694 49698 27746
rect 51774 27694 51826 27746
rect 52446 27694 52498 27746
rect 53342 27694 53394 27746
rect 10110 27582 10162 27634
rect 25678 27582 25730 27634
rect 33854 27582 33906 27634
rect 45950 27582 46002 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 14590 27246 14642 27298
rect 22990 27246 23042 27298
rect 45614 27246 45666 27298
rect 48414 27246 48466 27298
rect 50654 27246 50706 27298
rect 4174 27134 4226 27186
rect 5742 27134 5794 27186
rect 8430 27134 8482 27186
rect 9438 27134 9490 27186
rect 10334 27134 10386 27186
rect 12126 27134 12178 27186
rect 20862 27134 20914 27186
rect 23998 27134 24050 27186
rect 26014 27134 26066 27186
rect 27134 27134 27186 27186
rect 28702 27134 28754 27186
rect 29486 27134 29538 27186
rect 29934 27134 29986 27186
rect 38894 27134 38946 27186
rect 41358 27134 41410 27186
rect 41806 27134 41858 27186
rect 42702 27134 42754 27186
rect 43598 27134 43650 27186
rect 46174 27134 46226 27186
rect 48974 27134 49026 27186
rect 49534 27134 49586 27186
rect 49758 27134 49810 27186
rect 50430 27134 50482 27186
rect 50878 27134 50930 27186
rect 51214 27134 51266 27186
rect 57374 27134 57426 27186
rect 3054 27022 3106 27074
rect 3390 27022 3442 27074
rect 6750 27022 6802 27074
rect 7310 27022 7362 27074
rect 11230 27022 11282 27074
rect 11454 27022 11506 27074
rect 12014 27022 12066 27074
rect 13918 27022 13970 27074
rect 15374 27022 15426 27074
rect 17950 27022 18002 27074
rect 18510 27022 18562 27074
rect 22206 27022 22258 27074
rect 24222 27022 24274 27074
rect 25790 27022 25842 27074
rect 27022 27022 27074 27074
rect 28142 27022 28194 27074
rect 30942 27022 30994 27074
rect 32510 27022 32562 27074
rect 34190 27022 34242 27074
rect 34750 27022 34802 27074
rect 36206 27022 36258 27074
rect 36318 27022 36370 27074
rect 36542 27022 36594 27074
rect 37774 27022 37826 27074
rect 39230 27022 39282 27074
rect 40574 27022 40626 27074
rect 40910 27022 40962 27074
rect 45838 27022 45890 27074
rect 46062 27022 46114 27074
rect 47518 27022 47570 27074
rect 47742 27022 47794 27074
rect 51102 27022 51154 27074
rect 52782 27022 52834 27074
rect 53678 27022 53730 27074
rect 58046 27022 58098 27074
rect 4958 26910 5010 26962
rect 10894 26910 10946 26962
rect 12462 26910 12514 26962
rect 15822 26910 15874 26962
rect 16382 26910 16434 26962
rect 18958 26910 19010 26962
rect 21870 26910 21922 26962
rect 24894 26910 24946 26962
rect 26462 26910 26514 26962
rect 27246 26910 27298 26962
rect 28254 26910 28306 26962
rect 31278 26910 31330 26962
rect 32398 26910 32450 26962
rect 36654 26910 36706 26962
rect 39454 26910 39506 26962
rect 42254 26910 42306 26962
rect 43150 26910 43202 26962
rect 44046 26910 44098 26962
rect 47182 26910 47234 26962
rect 48302 26910 48354 26962
rect 51326 26910 51378 26962
rect 51998 26910 52050 26962
rect 53454 26910 53506 26962
rect 54014 26910 54066 26962
rect 57150 26910 57202 26962
rect 1934 26798 1986 26850
rect 7982 26798 8034 26850
rect 8990 26798 9042 26850
rect 11006 26798 11058 26850
rect 12238 26798 12290 26850
rect 19854 26798 19906 26850
rect 27470 26798 27522 26850
rect 32510 26798 32562 26850
rect 36430 26798 36482 26850
rect 40798 26798 40850 26850
rect 44494 26798 44546 26850
rect 46286 26798 46338 26850
rect 48414 26798 48466 26850
rect 49758 26798 49810 26850
rect 53678 26798 53730 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 1934 26462 1986 26514
rect 2942 26462 2994 26514
rect 3726 26462 3778 26514
rect 10334 26462 10386 26514
rect 20862 26462 20914 26514
rect 23886 26462 23938 26514
rect 24558 26462 24610 26514
rect 26238 26462 26290 26514
rect 28590 26462 28642 26514
rect 30830 26462 30882 26514
rect 32174 26462 32226 26514
rect 32958 26462 33010 26514
rect 35198 26462 35250 26514
rect 35310 26462 35362 26514
rect 37326 26462 37378 26514
rect 37774 26462 37826 26514
rect 38110 26462 38162 26514
rect 38558 26462 38610 26514
rect 40462 26462 40514 26514
rect 41806 26462 41858 26514
rect 43710 26462 43762 26514
rect 45390 26462 45442 26514
rect 46958 26462 47010 26514
rect 47406 26462 47458 26514
rect 50430 26462 50482 26514
rect 52110 26462 52162 26514
rect 54462 26462 54514 26514
rect 56478 26462 56530 26514
rect 56590 26462 56642 26514
rect 4846 26350 4898 26402
rect 11678 26350 11730 26402
rect 14030 26350 14082 26402
rect 21758 26350 21810 26402
rect 22766 26350 22818 26402
rect 23662 26350 23714 26402
rect 24894 26350 24946 26402
rect 25678 26350 25730 26402
rect 29486 26350 29538 26402
rect 30046 26350 30098 26402
rect 33966 26350 34018 26402
rect 34974 26350 35026 26402
rect 39230 26350 39282 26402
rect 43598 26350 43650 26402
rect 46062 26350 46114 26402
rect 54574 26350 54626 26402
rect 56254 26350 56306 26402
rect 2382 26238 2434 26290
rect 4174 26238 4226 26290
rect 5406 26238 5458 26290
rect 5966 26238 6018 26290
rect 8654 26238 8706 26290
rect 10670 26238 10722 26290
rect 11006 26238 11058 26290
rect 11230 26238 11282 26290
rect 12574 26238 12626 26290
rect 14142 26238 14194 26290
rect 15374 26238 15426 26290
rect 18734 26238 18786 26290
rect 21982 26238 22034 26290
rect 23550 26238 23602 26290
rect 26910 26238 26962 26290
rect 27134 26238 27186 26290
rect 27358 26238 27410 26290
rect 27582 26238 27634 26290
rect 28254 26238 28306 26290
rect 28366 26238 28418 26290
rect 28702 26238 28754 26290
rect 29710 26238 29762 26290
rect 33742 26238 33794 26290
rect 33854 26238 33906 26290
rect 34078 26238 34130 26290
rect 34190 26238 34242 26290
rect 35422 26238 35474 26290
rect 39566 26238 39618 26290
rect 40126 26238 40178 26290
rect 41694 26238 41746 26290
rect 41918 26238 41970 26290
rect 43150 26238 43202 26290
rect 43822 26238 43874 26290
rect 45614 26238 45666 26290
rect 48302 26238 48354 26290
rect 52894 26238 52946 26290
rect 56702 26238 56754 26290
rect 57598 26238 57650 26290
rect 57934 26238 57986 26290
rect 3278 26126 3330 26178
rect 7534 26126 7586 26178
rect 8542 26126 8594 26178
rect 9774 26126 9826 26178
rect 11454 26126 11506 26178
rect 11566 26126 11618 26178
rect 12910 26126 12962 26178
rect 15262 26126 15314 26178
rect 18622 26126 18674 26178
rect 20078 26126 20130 26178
rect 27470 26126 27522 26178
rect 28478 26126 28530 26178
rect 29374 26126 29426 26178
rect 31278 26126 31330 26178
rect 31726 26126 31778 26178
rect 35870 26126 35922 26178
rect 36430 26126 36482 26178
rect 36878 26126 36930 26178
rect 39902 26126 39954 26178
rect 42142 26126 42194 26178
rect 42366 26126 42418 26178
rect 44270 26126 44322 26178
rect 44718 26126 44770 26178
rect 45502 26126 45554 26178
rect 46510 26126 46562 26178
rect 47854 26126 47906 26178
rect 48750 26126 48802 26178
rect 49422 26126 49474 26178
rect 49870 26126 49922 26178
rect 53454 26126 53506 26178
rect 57486 26126 57538 26178
rect 12798 26014 12850 26066
rect 16494 26014 16546 26066
rect 25902 26014 25954 26066
rect 30270 26014 30322 26066
rect 30382 26014 30434 26066
rect 31166 26014 31218 26066
rect 31726 26014 31778 26066
rect 35982 26014 36034 26066
rect 36430 26014 36482 26066
rect 36878 26014 36930 26066
rect 42590 26014 42642 26066
rect 44046 26014 44098 26066
rect 44718 26014 44770 26066
rect 45838 26014 45890 26066
rect 46510 26014 46562 26066
rect 47518 26014 47570 26066
rect 47854 26014 47906 26066
rect 53678 26014 53730 26066
rect 54350 26014 54402 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 8990 25678 9042 25730
rect 9550 25678 9602 25730
rect 22094 25678 22146 25730
rect 22430 25678 22482 25730
rect 43822 25678 43874 25730
rect 2046 25566 2098 25618
rect 2942 25566 2994 25618
rect 4062 25566 4114 25618
rect 5854 25566 5906 25618
rect 6750 25566 6802 25618
rect 7870 25566 7922 25618
rect 8766 25566 8818 25618
rect 9214 25566 9266 25618
rect 9662 25566 9714 25618
rect 11678 25566 11730 25618
rect 13022 25566 13074 25618
rect 13806 25566 13858 25618
rect 14142 25566 14194 25618
rect 15262 25566 15314 25618
rect 16942 25566 16994 25618
rect 19070 25566 19122 25618
rect 20078 25566 20130 25618
rect 21870 25566 21922 25618
rect 22990 25566 23042 25618
rect 23550 25566 23602 25618
rect 26126 25566 26178 25618
rect 26910 25566 26962 25618
rect 33182 25566 33234 25618
rect 33966 25566 34018 25618
rect 36542 25566 36594 25618
rect 37438 25566 37490 25618
rect 38446 25566 38498 25618
rect 38782 25566 38834 25618
rect 39678 25566 39730 25618
rect 41022 25566 41074 25618
rect 41470 25566 41522 25618
rect 42366 25566 42418 25618
rect 43150 25566 43202 25618
rect 48862 25566 48914 25618
rect 51326 25566 51378 25618
rect 54350 25566 54402 25618
rect 55806 25566 55858 25618
rect 57150 25566 57202 25618
rect 6414 25454 6466 25506
rect 10110 25454 10162 25506
rect 10558 25454 10610 25506
rect 11790 25454 11842 25506
rect 12574 25454 12626 25506
rect 15374 25454 15426 25506
rect 18174 25454 18226 25506
rect 18398 25454 18450 25506
rect 24110 25454 24162 25506
rect 24670 25454 24722 25506
rect 27358 25454 27410 25506
rect 32174 25454 32226 25506
rect 32846 25454 32898 25506
rect 34190 25454 34242 25506
rect 40686 25454 40738 25506
rect 42814 25454 42866 25506
rect 43934 25454 43986 25506
rect 45838 25454 45890 25506
rect 46846 25454 46898 25506
rect 47630 25454 47682 25506
rect 49086 25454 49138 25506
rect 50542 25454 50594 25506
rect 50766 25454 50818 25506
rect 53902 25454 53954 25506
rect 55694 25454 55746 25506
rect 56926 25454 56978 25506
rect 57822 25454 57874 25506
rect 4062 25342 4114 25394
rect 10782 25342 10834 25394
rect 11342 25342 11394 25394
rect 16270 25342 16322 25394
rect 28254 25342 28306 25394
rect 30382 25342 30434 25394
rect 32062 25342 32114 25394
rect 34862 25342 34914 25394
rect 35534 25342 35586 25394
rect 37886 25342 37938 25394
rect 45502 25342 45554 25394
rect 47966 25342 48018 25394
rect 49758 25342 49810 25394
rect 50318 25342 50370 25394
rect 50878 25342 50930 25394
rect 53454 25342 53506 25394
rect 56030 25342 56082 25394
rect 2382 25230 2434 25282
rect 4846 25230 4898 25282
rect 7422 25230 7474 25282
rect 10446 25230 10498 25282
rect 11566 25230 11618 25282
rect 11902 25230 11954 25282
rect 20526 25230 20578 25282
rect 29822 25230 29874 25282
rect 31166 25230 31218 25282
rect 35758 25230 35810 25282
rect 35870 25230 35922 25282
rect 35982 25230 36034 25282
rect 39230 25230 39282 25282
rect 44046 25230 44098 25282
rect 44606 25230 44658 25282
rect 45614 25230 45666 25282
rect 46846 25230 46898 25282
rect 47854 25230 47906 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 2270 24894 2322 24946
rect 2718 24894 2770 24946
rect 3726 24894 3778 24946
rect 9886 24894 9938 24946
rect 11902 24894 11954 24946
rect 15710 24894 15762 24946
rect 16606 24894 16658 24946
rect 17054 24894 17106 24946
rect 19854 24894 19906 24946
rect 30382 24894 30434 24946
rect 30830 24894 30882 24946
rect 32062 24894 32114 24946
rect 34750 24894 34802 24946
rect 34862 24894 34914 24946
rect 36094 24894 36146 24946
rect 36654 24894 36706 24946
rect 40014 24894 40066 24946
rect 40462 24894 40514 24946
rect 41470 24894 41522 24946
rect 44382 24894 44434 24946
rect 45054 24894 45106 24946
rect 47742 24894 47794 24946
rect 48414 24894 48466 24946
rect 48638 24894 48690 24946
rect 49982 24894 50034 24946
rect 50094 24894 50146 24946
rect 57486 24894 57538 24946
rect 5742 24782 5794 24834
rect 8878 24782 8930 24834
rect 10446 24782 10498 24834
rect 11006 24782 11058 24834
rect 12238 24782 12290 24834
rect 13246 24782 13298 24834
rect 18734 24782 18786 24834
rect 21982 24782 22034 24834
rect 24446 24782 24498 24834
rect 26350 24782 26402 24834
rect 27582 24782 27634 24834
rect 29486 24782 29538 24834
rect 29934 24782 29986 24834
rect 33966 24782 34018 24834
rect 35870 24782 35922 24834
rect 47182 24782 47234 24834
rect 52782 24782 52834 24834
rect 55582 24782 55634 24834
rect 55694 24782 55746 24834
rect 4734 24670 4786 24722
rect 6974 24670 7026 24722
rect 7086 24670 7138 24722
rect 11566 24670 11618 24722
rect 11902 24670 11954 24722
rect 14142 24670 14194 24722
rect 14702 24670 14754 24722
rect 18062 24670 18114 24722
rect 20862 24670 20914 24722
rect 21422 24670 21474 24722
rect 23102 24670 23154 24722
rect 23774 24670 23826 24722
rect 26238 24670 26290 24722
rect 28366 24670 28418 24722
rect 31278 24670 31330 24722
rect 34190 24670 34242 24722
rect 34526 24670 34578 24722
rect 35646 24670 35698 24722
rect 36318 24670 36370 24722
rect 37438 24670 37490 24722
rect 38782 24670 38834 24722
rect 43038 24670 43090 24722
rect 43262 24670 43314 24722
rect 45390 24670 45442 24722
rect 47070 24670 47122 24722
rect 48750 24670 48802 24722
rect 53006 24670 53058 24722
rect 53342 24670 53394 24722
rect 57822 24670 57874 24722
rect 1934 24558 1986 24610
rect 3166 24558 3218 24610
rect 4958 24558 5010 24610
rect 16158 24558 16210 24610
rect 18398 24558 18450 24610
rect 19294 24558 19346 24610
rect 25790 24558 25842 24610
rect 32510 24558 32562 24610
rect 37326 24558 37378 24610
rect 42366 24558 42418 24610
rect 43934 24558 43986 24610
rect 53230 24558 53282 24610
rect 58046 24558 58098 24610
rect 2046 24446 2098 24498
rect 2718 24446 2770 24498
rect 3278 24446 3330 24498
rect 10222 24446 10274 24498
rect 19518 24446 19570 24498
rect 28590 24446 28642 24498
rect 28926 24446 28978 24498
rect 39454 24446 39506 24498
rect 40014 24446 40066 24498
rect 40462 24446 40514 24498
rect 44158 24446 44210 24498
rect 44830 24446 44882 24498
rect 46062 24446 46114 24498
rect 46398 24446 46450 24498
rect 50206 24446 50258 24498
rect 55582 24446 55634 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 3390 24110 3442 24162
rect 4510 24110 4562 24162
rect 11790 24110 11842 24162
rect 32398 24110 32450 24162
rect 41134 24110 41186 24162
rect 1822 23998 1874 24050
rect 2382 23998 2434 24050
rect 2718 23998 2770 24050
rect 3278 23998 3330 24050
rect 3726 23998 3778 24050
rect 4062 23998 4114 24050
rect 4510 23998 4562 24050
rect 7646 23998 7698 24050
rect 12462 23998 12514 24050
rect 13022 23998 13074 24050
rect 15150 23998 15202 24050
rect 18286 23998 18338 24050
rect 18734 23998 18786 24050
rect 19182 23998 19234 24050
rect 19518 23998 19570 24050
rect 22094 23998 22146 24050
rect 23662 23998 23714 24050
rect 26798 23998 26850 24050
rect 28478 23998 28530 24050
rect 33406 23998 33458 24050
rect 33854 23998 33906 24050
rect 34750 23998 34802 24050
rect 37774 23998 37826 24050
rect 39006 23998 39058 24050
rect 39566 23998 39618 24050
rect 39902 23998 39954 24050
rect 40462 23998 40514 24050
rect 44382 23998 44434 24050
rect 45614 23998 45666 24050
rect 46958 23998 47010 24050
rect 48526 23998 48578 24050
rect 54686 23998 54738 24050
rect 6750 23886 6802 23938
rect 7086 23886 7138 23938
rect 8654 23886 8706 23938
rect 8766 23886 8818 23938
rect 11230 23886 11282 23938
rect 11454 23886 11506 23938
rect 13918 23886 13970 23938
rect 14590 23886 14642 23938
rect 20190 23886 20242 23938
rect 20638 23886 20690 23938
rect 21758 23886 21810 23938
rect 21870 23886 21922 23938
rect 22206 23886 22258 23938
rect 25454 23886 25506 23938
rect 26014 23886 26066 23938
rect 27470 23886 27522 23938
rect 28030 23886 28082 23938
rect 29598 23886 29650 23938
rect 30942 23886 30994 23938
rect 31950 23886 32002 23938
rect 36094 23886 36146 23938
rect 37550 23886 37602 23938
rect 37998 23886 38050 23938
rect 38334 23886 38386 23938
rect 40910 23886 40962 23938
rect 42926 23886 42978 23938
rect 43150 23886 43202 23938
rect 45838 23886 45890 23938
rect 50206 23886 50258 23938
rect 54126 23886 54178 23938
rect 54462 23886 54514 23938
rect 56366 23886 56418 23938
rect 57262 23886 57314 23938
rect 4958 23774 5010 23826
rect 10558 23774 10610 23826
rect 11678 23774 11730 23826
rect 17614 23774 17666 23826
rect 23774 23774 23826 23826
rect 25118 23774 25170 23826
rect 28366 23774 28418 23826
rect 32174 23774 32226 23826
rect 34974 23774 35026 23826
rect 36766 23774 36818 23826
rect 38222 23774 38274 23826
rect 41470 23774 41522 23826
rect 42478 23774 42530 23826
rect 42702 23774 42754 23826
rect 46510 23774 46562 23826
rect 49086 23774 49138 23826
rect 50654 23774 50706 23826
rect 55134 23774 55186 23826
rect 56142 23774 56194 23826
rect 57934 23774 57986 23826
rect 16382 23662 16434 23714
rect 16830 23662 16882 23714
rect 20750 23662 20802 23714
rect 22990 23662 23042 23714
rect 23550 23662 23602 23714
rect 38446 23662 38498 23714
rect 47518 23662 47570 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 2046 23326 2098 23378
rect 2830 23326 2882 23378
rect 3838 23326 3890 23378
rect 5630 23326 5682 23378
rect 5966 23326 6018 23378
rect 9662 23326 9714 23378
rect 11790 23326 11842 23378
rect 12126 23326 12178 23378
rect 13470 23326 13522 23378
rect 14030 23326 14082 23378
rect 14478 23326 14530 23378
rect 14926 23326 14978 23378
rect 17950 23326 18002 23378
rect 19854 23326 19906 23378
rect 26574 23326 26626 23378
rect 30606 23326 30658 23378
rect 32062 23326 32114 23378
rect 32398 23326 32450 23378
rect 33630 23326 33682 23378
rect 36206 23326 36258 23378
rect 39902 23326 39954 23378
rect 40014 23326 40066 23378
rect 46398 23326 46450 23378
rect 55694 23326 55746 23378
rect 56142 23326 56194 23378
rect 4622 23214 4674 23266
rect 5070 23214 5122 23266
rect 8990 23214 9042 23266
rect 10894 23214 10946 23266
rect 12798 23214 12850 23266
rect 18510 23214 18562 23266
rect 22318 23214 22370 23266
rect 24670 23214 24722 23266
rect 24782 23214 24834 23266
rect 26126 23214 26178 23266
rect 32174 23214 32226 23266
rect 35086 23214 35138 23266
rect 36766 23214 36818 23266
rect 36990 23214 37042 23266
rect 37214 23214 37266 23266
rect 37550 23214 37602 23266
rect 51102 23214 51154 23266
rect 51326 23214 51378 23266
rect 6638 23102 6690 23154
rect 8094 23102 8146 23154
rect 11230 23102 11282 23154
rect 12910 23102 12962 23154
rect 15486 23102 15538 23154
rect 16718 23102 16770 23154
rect 16942 23102 16994 23154
rect 17838 23102 17890 23154
rect 21310 23102 21362 23154
rect 26014 23102 26066 23154
rect 27470 23102 27522 23154
rect 30718 23102 30770 23154
rect 30942 23102 30994 23154
rect 31166 23102 31218 23154
rect 31390 23102 31442 23154
rect 32622 23102 32674 23154
rect 34638 23102 34690 23154
rect 34750 23102 34802 23154
rect 35870 23102 35922 23154
rect 38222 23102 38274 23154
rect 39678 23102 39730 23154
rect 40126 23102 40178 23154
rect 40238 23102 40290 23154
rect 41694 23102 41746 23154
rect 42030 23102 42082 23154
rect 42590 23102 42642 23154
rect 43262 23102 43314 23154
rect 43486 23102 43538 23154
rect 44830 23102 44882 23154
rect 45054 23102 45106 23154
rect 47182 23102 47234 23154
rect 50990 23102 51042 23154
rect 52670 23102 52722 23154
rect 53342 23102 53394 23154
rect 54350 23102 54402 23154
rect 2382 22990 2434 23042
rect 3278 22990 3330 23042
rect 4174 22990 4226 23042
rect 6974 22990 7026 23042
rect 8654 22990 8706 23042
rect 10110 22990 10162 23042
rect 16046 22990 16098 23042
rect 18958 22990 19010 23042
rect 19518 22990 19570 23042
rect 20414 22990 20466 23042
rect 20750 22990 20802 23042
rect 23102 22990 23154 23042
rect 23662 22990 23714 23042
rect 29262 22990 29314 23042
rect 32174 22990 32226 23042
rect 33966 22990 34018 23042
rect 35646 22990 35698 23042
rect 37102 22990 37154 23042
rect 38446 22990 38498 23042
rect 38782 22990 38834 23042
rect 40798 22990 40850 23042
rect 44158 22990 44210 23042
rect 45726 22990 45778 23042
rect 47070 22990 47122 23042
rect 47854 22990 47906 23042
rect 48302 22990 48354 23042
rect 53454 22990 53506 23042
rect 54462 22990 54514 23042
rect 1934 22878 1986 22930
rect 2382 22878 2434 22930
rect 2942 22878 2994 22930
rect 3278 22878 3330 22930
rect 4958 22878 5010 22930
rect 11566 22878 11618 22930
rect 11902 22878 11954 22930
rect 12126 22878 12178 22930
rect 12798 22878 12850 22930
rect 17950 22878 18002 22930
rect 24782 22878 24834 22930
rect 34974 22878 35026 22930
rect 54686 22878 54738 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 3502 22542 3554 22594
rect 3726 22542 3778 22594
rect 4398 22542 4450 22594
rect 4958 22542 5010 22594
rect 30158 22542 30210 22594
rect 41134 22542 41186 22594
rect 41918 22542 41970 22594
rect 46734 22542 46786 22594
rect 2158 22430 2210 22482
rect 2606 22430 2658 22482
rect 3502 22430 3554 22482
rect 4062 22430 4114 22482
rect 4398 22430 4450 22482
rect 5966 22430 6018 22482
rect 8206 22430 8258 22482
rect 9550 22430 9602 22482
rect 10222 22430 10274 22482
rect 10670 22430 10722 22482
rect 11566 22430 11618 22482
rect 14814 22430 14866 22482
rect 15598 22430 15650 22482
rect 17278 22430 17330 22482
rect 18734 22430 18786 22482
rect 21646 22430 21698 22482
rect 21982 22430 22034 22482
rect 22542 22430 22594 22482
rect 23550 22430 23602 22482
rect 25790 22430 25842 22482
rect 27358 22430 27410 22482
rect 28478 22430 28530 22482
rect 29710 22430 29762 22482
rect 30382 22430 30434 22482
rect 31614 22430 31666 22482
rect 32286 22430 32338 22482
rect 32622 22430 32674 22482
rect 34862 22430 34914 22482
rect 35646 22430 35698 22482
rect 36094 22430 36146 22482
rect 37438 22430 37490 22482
rect 39342 22430 39394 22482
rect 41918 22430 41970 22482
rect 42814 22430 42866 22482
rect 43262 22430 43314 22482
rect 43934 22430 43986 22482
rect 48190 22430 48242 22482
rect 56366 22430 56418 22482
rect 4846 22318 4898 22370
rect 7870 22318 7922 22370
rect 12798 22318 12850 22370
rect 13918 22318 13970 22370
rect 17054 22318 17106 22370
rect 18398 22318 18450 22370
rect 20190 22318 20242 22370
rect 20862 22318 20914 22370
rect 22990 22318 23042 22370
rect 24222 22318 24274 22370
rect 25902 22318 25954 22370
rect 27582 22318 27634 22370
rect 30606 22318 30658 22370
rect 30830 22318 30882 22370
rect 33518 22318 33570 22370
rect 33854 22318 33906 22370
rect 33966 22318 34018 22370
rect 44494 22318 44546 22370
rect 44830 22318 44882 22370
rect 45502 22318 45554 22370
rect 46062 22318 46114 22370
rect 50542 22318 50594 22370
rect 50990 22318 51042 22370
rect 54014 22318 54066 22370
rect 54462 22318 54514 22370
rect 57262 22318 57314 22370
rect 6414 22206 6466 22258
rect 7422 22206 7474 22258
rect 11118 22206 11170 22258
rect 13806 22206 13858 22258
rect 16382 22206 16434 22258
rect 17950 22206 18002 22258
rect 24782 22206 24834 22258
rect 27918 22206 27970 22258
rect 40126 22206 40178 22258
rect 40574 22206 40626 22258
rect 47742 22206 47794 22258
rect 51214 22206 51266 22258
rect 51774 22206 51826 22258
rect 51998 22206 52050 22258
rect 52222 22206 52274 22258
rect 52334 22206 52386 22258
rect 55134 22206 55186 22258
rect 56030 22206 56082 22258
rect 1822 22094 1874 22146
rect 3054 22094 3106 22146
rect 6862 22094 6914 22146
rect 9102 22094 9154 22146
rect 12126 22094 12178 22146
rect 12238 22094 12290 22146
rect 12350 22094 12402 22146
rect 13582 22094 13634 22146
rect 15150 22094 15202 22146
rect 19518 22094 19570 22146
rect 19630 22094 19682 22146
rect 19742 22094 19794 22146
rect 20526 22094 20578 22146
rect 20750 22094 20802 22146
rect 23438 22094 23490 22146
rect 23662 22094 23714 22146
rect 28814 22094 28866 22146
rect 30718 22094 30770 22146
rect 34078 22094 34130 22146
rect 34190 22094 34242 22146
rect 35198 22094 35250 22146
rect 36542 22094 36594 22146
rect 37886 22094 37938 22146
rect 38334 22094 38386 22146
rect 38782 22094 38834 22146
rect 40350 22094 40402 22146
rect 40686 22094 40738 22146
rect 41022 22094 41074 22146
rect 41470 22094 41522 22146
rect 42366 22094 42418 22146
rect 44606 22094 44658 22146
rect 45950 22094 46002 22146
rect 46174 22094 46226 22146
rect 46846 22094 46898 22146
rect 46958 22094 47010 22146
rect 47630 22094 47682 22146
rect 48638 22094 48690 22146
rect 58158 22094 58210 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 2158 21758 2210 21810
rect 2718 21758 2770 21810
rect 3502 21758 3554 21810
rect 5406 21758 5458 21810
rect 7310 21758 7362 21810
rect 8990 21758 9042 21810
rect 9998 21758 10050 21810
rect 11454 21758 11506 21810
rect 14478 21758 14530 21810
rect 17838 21758 17890 21810
rect 17950 21758 18002 21810
rect 18622 21758 18674 21810
rect 25678 21758 25730 21810
rect 29150 21758 29202 21810
rect 29486 21758 29538 21810
rect 30382 21758 30434 21810
rect 30830 21758 30882 21810
rect 34862 21758 34914 21810
rect 35310 21758 35362 21810
rect 37214 21758 37266 21810
rect 37774 21758 37826 21810
rect 38222 21758 38274 21810
rect 40574 21758 40626 21810
rect 43374 21758 43426 21810
rect 47406 21758 47458 21810
rect 51662 21758 51714 21810
rect 54126 21758 54178 21810
rect 1822 21646 1874 21698
rect 5854 21646 5906 21698
rect 6190 21646 6242 21698
rect 7982 21646 8034 21698
rect 10558 21646 10610 21698
rect 16606 21646 16658 21698
rect 16942 21646 16994 21698
rect 20526 21646 20578 21698
rect 23102 21646 23154 21698
rect 24558 21646 24610 21698
rect 28926 21646 28978 21698
rect 30606 21646 30658 21698
rect 32510 21646 32562 21698
rect 32734 21646 32786 21698
rect 36318 21646 36370 21698
rect 43486 21646 43538 21698
rect 45054 21646 45106 21698
rect 48302 21646 48354 21698
rect 48414 21646 48466 21698
rect 50542 21646 50594 21698
rect 53566 21646 53618 21698
rect 3054 21534 3106 21586
rect 4846 21534 4898 21586
rect 6638 21534 6690 21586
rect 7870 21534 7922 21586
rect 10334 21534 10386 21586
rect 10670 21534 10722 21586
rect 12238 21534 12290 21586
rect 12910 21534 12962 21586
rect 13246 21534 13298 21586
rect 15598 21534 15650 21586
rect 15822 21534 15874 21586
rect 18062 21534 18114 21586
rect 18846 21534 18898 21586
rect 19294 21534 19346 21586
rect 20078 21534 20130 21586
rect 20302 21534 20354 21586
rect 21310 21534 21362 21586
rect 22206 21534 22258 21586
rect 24446 21534 24498 21586
rect 24670 21534 24722 21586
rect 26350 21534 26402 21586
rect 26686 21534 26738 21586
rect 29374 21534 29426 21586
rect 33854 21534 33906 21586
rect 35870 21534 35922 21586
rect 36094 21534 36146 21586
rect 36542 21534 36594 21586
rect 37102 21534 37154 21586
rect 37438 21534 37490 21586
rect 39230 21534 39282 21586
rect 39790 21534 39842 21586
rect 41470 21534 41522 21586
rect 43150 21534 43202 21586
rect 43822 21534 43874 21586
rect 45726 21534 45778 21586
rect 45950 21534 46002 21586
rect 47182 21534 47234 21586
rect 47294 21534 47346 21586
rect 47854 21534 47906 21586
rect 49646 21534 49698 21586
rect 49870 21534 49922 21586
rect 51102 21534 51154 21586
rect 53790 21534 53842 21586
rect 55358 21534 55410 21586
rect 57486 21534 57538 21586
rect 57710 21534 57762 21586
rect 58046 21534 58098 21586
rect 58494 21534 58546 21586
rect 3950 21422 4002 21474
rect 4398 21422 4450 21474
rect 8542 21422 8594 21474
rect 11790 21422 11842 21474
rect 12574 21422 12626 21474
rect 14926 21422 14978 21474
rect 18734 21422 18786 21474
rect 22318 21422 22370 21474
rect 23550 21422 23602 21474
rect 27806 21422 27858 21474
rect 28366 21422 28418 21474
rect 29262 21422 29314 21474
rect 30494 21422 30546 21474
rect 31614 21422 31666 21474
rect 32846 21422 32898 21474
rect 33966 21422 34018 21474
rect 34414 21422 34466 21474
rect 36654 21422 36706 21474
rect 41918 21422 41970 21474
rect 42590 21422 42642 21474
rect 43934 21422 43986 21474
rect 44494 21422 44546 21474
rect 44718 21422 44770 21474
rect 46622 21422 46674 21474
rect 47854 21422 47906 21474
rect 48078 21422 48130 21474
rect 52110 21422 52162 21474
rect 55582 21422 55634 21474
rect 56702 21422 56754 21474
rect 57598 21422 57650 21474
rect 3502 21310 3554 21362
rect 4174 21310 4226 21362
rect 11790 21310 11842 21362
rect 12014 21310 12066 21362
rect 20638 21310 20690 21362
rect 22206 21310 22258 21362
rect 38894 21310 38946 21362
rect 39230 21310 39282 21362
rect 48414 21310 48466 21362
rect 51326 21310 51378 21362
rect 55022 21310 55074 21362
rect 56142 21310 56194 21362
rect 56478 21310 56530 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 3950 20974 4002 21026
rect 4510 20974 4562 21026
rect 12910 20974 12962 21026
rect 13694 20974 13746 21026
rect 21870 20974 21922 21026
rect 23326 20974 23378 21026
rect 30942 20974 30994 21026
rect 31614 20974 31666 21026
rect 31950 20974 32002 21026
rect 34750 20974 34802 21026
rect 39118 20974 39170 21026
rect 39902 20974 39954 21026
rect 40686 20974 40738 21026
rect 2270 20862 2322 20914
rect 2718 20862 2770 20914
rect 3166 20862 3218 20914
rect 4062 20862 4114 20914
rect 4510 20862 4562 20914
rect 4958 20862 5010 20914
rect 5630 20862 5682 20914
rect 6078 20862 6130 20914
rect 7534 20862 7586 20914
rect 9774 20862 9826 20914
rect 15822 20862 15874 20914
rect 17166 20862 17218 20914
rect 18062 20862 18114 20914
rect 19070 20862 19122 20914
rect 20190 20862 20242 20914
rect 24334 20862 24386 20914
rect 25902 20862 25954 20914
rect 26574 20862 26626 20914
rect 26686 20862 26738 20914
rect 36094 20862 36146 20914
rect 36766 20862 36818 20914
rect 39902 20862 39954 20914
rect 43038 20862 43090 20914
rect 45726 20862 45778 20914
rect 46398 20862 46450 20914
rect 49310 20862 49362 20914
rect 50542 20862 50594 20914
rect 57374 20862 57426 20914
rect 7310 20750 7362 20802
rect 9438 20750 9490 20802
rect 11790 20750 11842 20802
rect 15150 20750 15202 20802
rect 16494 20750 16546 20802
rect 17726 20750 17778 20802
rect 19518 20750 19570 20802
rect 21758 20750 21810 20802
rect 22094 20750 22146 20802
rect 26910 20750 26962 20802
rect 27358 20750 27410 20802
rect 27806 20750 27858 20802
rect 28366 20750 28418 20802
rect 28590 20750 28642 20802
rect 30270 20750 30322 20802
rect 32510 20750 32562 20802
rect 32958 20750 33010 20802
rect 33630 20750 33682 20802
rect 34078 20750 34130 20802
rect 34190 20750 34242 20802
rect 35534 20750 35586 20802
rect 35758 20750 35810 20802
rect 37550 20750 37602 20802
rect 37886 20750 37938 20802
rect 38110 20750 38162 20802
rect 41022 20750 41074 20802
rect 42030 20750 42082 20802
rect 42366 20750 42418 20802
rect 42590 20750 42642 20802
rect 46510 20750 46562 20802
rect 47854 20750 47906 20802
rect 50878 20750 50930 20802
rect 54350 20750 54402 20802
rect 56366 20750 56418 20802
rect 57262 20750 57314 20802
rect 6638 20638 6690 20690
rect 8990 20638 9042 20690
rect 10894 20638 10946 20690
rect 11566 20638 11618 20690
rect 12798 20638 12850 20690
rect 13918 20638 13970 20690
rect 22654 20638 22706 20690
rect 23214 20638 23266 20690
rect 23998 20638 24050 20690
rect 25006 20638 25058 20690
rect 26462 20638 26514 20690
rect 27134 20638 27186 20690
rect 28142 20638 28194 20690
rect 28814 20638 28866 20690
rect 29822 20638 29874 20690
rect 40462 20638 40514 20690
rect 48638 20638 48690 20690
rect 51326 20638 51378 20690
rect 54686 20638 54738 20690
rect 56030 20638 56082 20690
rect 56702 20638 56754 20690
rect 1934 20526 1986 20578
rect 3614 20526 3666 20578
rect 8430 20526 8482 20578
rect 11678 20526 11730 20578
rect 12238 20526 12290 20578
rect 13806 20526 13858 20578
rect 14814 20526 14866 20578
rect 16270 20526 16322 20578
rect 18510 20526 18562 20578
rect 23326 20526 23378 20578
rect 24222 20526 24274 20578
rect 25454 20526 25506 20578
rect 28366 20526 28418 20578
rect 31838 20526 31890 20578
rect 35982 20526 36034 20578
rect 36094 20526 36146 20578
rect 37998 20526 38050 20578
rect 38558 20526 38610 20578
rect 39006 20526 39058 20578
rect 39454 20526 39506 20578
rect 42478 20526 42530 20578
rect 53790 20526 53842 20578
rect 54462 20526 54514 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 2718 20190 2770 20242
rect 5294 20190 5346 20242
rect 5854 20190 5906 20242
rect 7870 20190 7922 20242
rect 17838 20190 17890 20242
rect 20526 20190 20578 20242
rect 21422 20190 21474 20242
rect 23662 20190 23714 20242
rect 23886 20190 23938 20242
rect 24446 20190 24498 20242
rect 30830 20190 30882 20242
rect 31838 20190 31890 20242
rect 40014 20190 40066 20242
rect 40910 20190 40962 20242
rect 46062 20190 46114 20242
rect 47854 20190 47906 20242
rect 48302 20190 48354 20242
rect 56478 20190 56530 20242
rect 4510 20078 4562 20130
rect 4958 20078 5010 20130
rect 6190 20078 6242 20130
rect 11678 20078 11730 20130
rect 14478 20078 14530 20130
rect 18286 20078 18338 20130
rect 18846 20078 18898 20130
rect 21310 20078 21362 20130
rect 21646 20078 21698 20130
rect 22094 20078 22146 20130
rect 23550 20078 23602 20130
rect 25006 20078 25058 20130
rect 27246 20078 27298 20130
rect 27806 20078 27858 20130
rect 28030 20078 28082 20130
rect 30158 20078 30210 20130
rect 32062 20078 32114 20130
rect 32734 20078 32786 20130
rect 35870 20078 35922 20130
rect 36542 20078 36594 20130
rect 36766 20078 36818 20130
rect 37550 20078 37602 20130
rect 39118 20078 39170 20130
rect 53454 20078 53506 20130
rect 54798 20078 54850 20130
rect 56590 20078 56642 20130
rect 57486 20078 57538 20130
rect 3054 19966 3106 20018
rect 3502 19966 3554 20018
rect 7086 19966 7138 20018
rect 7198 19966 7250 20018
rect 7646 19966 7698 20018
rect 10670 19966 10722 20018
rect 12014 19966 12066 20018
rect 12574 19966 12626 20018
rect 13246 19966 13298 20018
rect 16494 19966 16546 20018
rect 19742 19966 19794 20018
rect 28702 19966 28754 20018
rect 28926 19966 28978 20018
rect 29822 19966 29874 20018
rect 30942 19966 30994 20018
rect 31726 19966 31778 20018
rect 33854 19966 33906 20018
rect 34862 19966 34914 20018
rect 36430 19966 36482 20018
rect 42254 19966 42306 20018
rect 56030 19966 56082 20018
rect 56254 19966 56306 20018
rect 57598 19966 57650 20018
rect 57822 19966 57874 20018
rect 1822 19854 1874 19906
rect 2270 19854 2322 19906
rect 3950 19854 4002 19906
rect 6862 19854 6914 19906
rect 8206 19854 8258 19906
rect 8990 19854 9042 19906
rect 9998 19854 10050 19906
rect 10782 19854 10834 19906
rect 13358 19854 13410 19906
rect 15262 19854 15314 19906
rect 15598 19854 15650 19906
rect 16046 19854 16098 19906
rect 17054 19854 17106 19906
rect 19182 19854 19234 19906
rect 23102 19854 23154 19906
rect 25678 19854 25730 19906
rect 26014 19854 26066 19906
rect 26462 19854 26514 19906
rect 28142 19854 28194 19906
rect 32846 19854 32898 19906
rect 34190 19854 34242 19906
rect 34638 19854 34690 19906
rect 37438 19854 37490 19906
rect 39454 19854 39506 19906
rect 40350 19854 40402 19906
rect 42478 19854 42530 19906
rect 42926 19854 42978 19906
rect 52222 19854 52274 19906
rect 52894 19854 52946 19906
rect 55022 19854 55074 19906
rect 55470 19854 55522 19906
rect 56590 19854 56642 19906
rect 16046 19742 16098 19794
rect 16718 19742 16770 19794
rect 22206 19742 22258 19794
rect 29262 19742 29314 19794
rect 32510 19742 32562 19794
rect 34974 19742 35026 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 6862 19406 6914 19458
rect 7422 19406 7474 19458
rect 12798 19406 12850 19458
rect 13134 19406 13186 19458
rect 19070 19406 19122 19458
rect 19294 19406 19346 19458
rect 20526 19406 20578 19458
rect 20862 19406 20914 19458
rect 30382 19406 30434 19458
rect 30718 19406 30770 19458
rect 33854 19406 33906 19458
rect 34078 19406 34130 19458
rect 34862 19406 34914 19458
rect 2382 19294 2434 19346
rect 5070 19294 5122 19346
rect 5854 19294 5906 19346
rect 6302 19294 6354 19346
rect 6750 19294 6802 19346
rect 7086 19294 7138 19346
rect 7534 19294 7586 19346
rect 7982 19294 8034 19346
rect 8990 19294 9042 19346
rect 10558 19294 10610 19346
rect 11006 19294 11058 19346
rect 11454 19294 11506 19346
rect 12126 19294 12178 19346
rect 12574 19294 12626 19346
rect 14366 19294 14418 19346
rect 19406 19294 19458 19346
rect 20414 19294 20466 19346
rect 23774 19294 23826 19346
rect 26462 19294 26514 19346
rect 27134 19294 27186 19346
rect 27582 19294 27634 19346
rect 28366 19294 28418 19346
rect 28814 19294 28866 19346
rect 30382 19294 30434 19346
rect 31166 19294 31218 19346
rect 32958 19294 33010 19346
rect 33406 19294 33458 19346
rect 33854 19294 33906 19346
rect 34302 19294 34354 19346
rect 34750 19294 34802 19346
rect 35758 19294 35810 19346
rect 38446 19294 38498 19346
rect 9886 19182 9938 19234
rect 15374 19182 15426 19234
rect 16046 19182 16098 19234
rect 22318 19182 22370 19234
rect 39118 19406 39170 19458
rect 46062 19406 46114 19458
rect 38782 19294 38834 19346
rect 39342 19294 39394 19346
rect 40910 19294 40962 19346
rect 42926 19294 42978 19346
rect 46398 19294 46450 19346
rect 23102 19182 23154 19234
rect 25006 19182 25058 19234
rect 32622 19182 32674 19234
rect 36206 19182 36258 19234
rect 37886 19182 37938 19234
rect 38670 19182 38722 19234
rect 41470 19182 41522 19234
rect 41806 19182 41858 19234
rect 42590 19182 42642 19234
rect 44046 19182 44098 19234
rect 46846 19182 46898 19234
rect 49086 19182 49138 19234
rect 49422 19182 49474 19234
rect 49870 19182 49922 19234
rect 53678 19182 53730 19234
rect 54350 19182 54402 19234
rect 55470 19182 55522 19234
rect 57934 19182 57986 19234
rect 58382 19182 58434 19234
rect 22094 19070 22146 19122
rect 22990 19070 23042 19122
rect 24334 19070 24386 19122
rect 26126 19070 26178 19122
rect 36654 19070 36706 19122
rect 41582 19070 41634 19122
rect 43486 19070 43538 19122
rect 44158 19070 44210 19122
rect 44718 19070 44770 19122
rect 45838 19070 45890 19122
rect 47406 19070 47458 19122
rect 49198 19070 49250 19122
rect 51326 19070 51378 19122
rect 52670 19070 52722 19122
rect 53902 19070 53954 19122
rect 55358 19070 55410 19122
rect 2718 18958 2770 19010
rect 3166 18958 3218 19010
rect 3614 18958 3666 19010
rect 4062 18958 4114 19010
rect 4510 18958 4562 19010
rect 8430 18958 8482 19010
rect 9550 18958 9602 19010
rect 12910 18958 12962 19010
rect 13582 18958 13634 19010
rect 14702 18958 14754 19010
rect 18286 18958 18338 19010
rect 19966 18958 20018 19010
rect 20862 18958 20914 19010
rect 22206 18958 22258 19010
rect 22766 18958 22818 19010
rect 27918 18958 27970 19010
rect 29486 18958 29538 19010
rect 30718 18958 30770 19010
rect 31614 18958 31666 19010
rect 32062 18958 32114 19010
rect 37438 18958 37490 19010
rect 40238 18958 40290 19010
rect 44382 18958 44434 19010
rect 47294 18958 47346 19010
rect 47518 18958 47570 19010
rect 50318 18958 50370 19010
rect 50430 18958 50482 19010
rect 50542 18958 50594 19010
rect 51438 18958 51490 19010
rect 51662 18958 51714 19010
rect 54126 18958 54178 19010
rect 56030 18958 56082 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 4174 18622 4226 18674
rect 10558 18622 10610 18674
rect 11342 18622 11394 18674
rect 17054 18622 17106 18674
rect 21086 18622 21138 18674
rect 25678 18622 25730 18674
rect 27022 18622 27074 18674
rect 27806 18622 27858 18674
rect 33518 18622 33570 18674
rect 35310 18622 35362 18674
rect 37438 18622 37490 18674
rect 39678 18622 39730 18674
rect 40910 18622 40962 18674
rect 42926 18622 42978 18674
rect 43486 18622 43538 18674
rect 57598 18622 57650 18674
rect 57710 18622 57762 18674
rect 3726 18510 3778 18562
rect 7982 18510 8034 18562
rect 16270 18510 16322 18562
rect 22654 18510 22706 18562
rect 23550 18510 23602 18562
rect 23886 18510 23938 18562
rect 25902 18510 25954 18562
rect 26910 18510 26962 18562
rect 27918 18510 27970 18562
rect 29598 18510 29650 18562
rect 29822 18510 29874 18562
rect 30158 18510 30210 18562
rect 32174 18510 32226 18562
rect 34414 18510 34466 18562
rect 34750 18510 34802 18562
rect 38782 18510 38834 18562
rect 39006 18510 39058 18562
rect 41582 18510 41634 18562
rect 52782 18510 52834 18562
rect 54014 18510 54066 18562
rect 57822 18510 57874 18562
rect 3390 18398 3442 18450
rect 5070 18398 5122 18450
rect 5742 18398 5794 18450
rect 8766 18398 8818 18450
rect 10110 18398 10162 18450
rect 12126 18398 12178 18450
rect 12574 18398 12626 18450
rect 13582 18398 13634 18450
rect 14030 18398 14082 18450
rect 17838 18398 17890 18450
rect 21310 18398 21362 18450
rect 24558 18398 24610 18450
rect 24782 18398 24834 18450
rect 24894 18398 24946 18450
rect 26350 18398 26402 18450
rect 27582 18398 27634 18450
rect 28366 18398 28418 18450
rect 31502 18398 31554 18450
rect 32286 18398 32338 18450
rect 34190 18398 34242 18450
rect 36094 18398 36146 18450
rect 37102 18398 37154 18450
rect 38558 18398 38610 18450
rect 39118 18398 39170 18450
rect 40238 18398 40290 18450
rect 43598 18398 43650 18450
rect 43710 18398 43762 18450
rect 44158 18398 44210 18450
rect 45614 18398 45666 18450
rect 46510 18398 46562 18450
rect 47854 18398 47906 18450
rect 48078 18398 48130 18450
rect 49982 18398 50034 18450
rect 51662 18398 51714 18450
rect 52110 18398 52162 18450
rect 54910 18398 54962 18450
rect 57934 18398 57986 18450
rect 4622 18286 4674 18338
rect 11678 18286 11730 18338
rect 18398 18286 18450 18338
rect 18734 18286 18786 18338
rect 19182 18286 19234 18338
rect 19630 18286 19682 18338
rect 20078 18286 20130 18338
rect 22878 18286 22930 18338
rect 25790 18286 25842 18338
rect 28814 18286 28866 18338
rect 29486 18286 29538 18338
rect 30382 18286 30434 18338
rect 31054 18286 31106 18338
rect 32734 18286 32786 18338
rect 34638 18286 34690 18338
rect 35758 18286 35810 18338
rect 36542 18286 36594 18338
rect 37886 18286 37938 18338
rect 44494 18286 44546 18338
rect 46062 18286 46114 18338
rect 48750 18286 48802 18338
rect 50094 18286 50146 18338
rect 52222 18286 52274 18338
rect 53454 18286 53506 18338
rect 56030 18286 56082 18338
rect 11118 18174 11170 18226
rect 11342 18174 11394 18226
rect 11678 18174 11730 18226
rect 17726 18174 17778 18226
rect 18510 18174 18562 18226
rect 18734 18174 18786 18226
rect 20190 18174 20242 18226
rect 27134 18174 27186 18226
rect 30494 18174 30546 18226
rect 34974 18174 35026 18226
rect 36542 18174 36594 18226
rect 41806 18174 41858 18226
rect 42142 18174 42194 18226
rect 50318 18174 50370 18226
rect 58270 18174 58322 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 13022 17838 13074 17890
rect 13582 17838 13634 17890
rect 15374 17838 15426 17890
rect 22990 17838 23042 17890
rect 23774 17838 23826 17890
rect 24446 17838 24498 17890
rect 27582 17838 27634 17890
rect 28030 17838 28082 17890
rect 30830 17838 30882 17890
rect 33070 17838 33122 17890
rect 37662 17838 37714 17890
rect 37998 17838 38050 17890
rect 48974 17838 49026 17890
rect 50094 17838 50146 17890
rect 4062 17726 4114 17778
rect 4510 17726 4562 17778
rect 4958 17726 5010 17778
rect 5742 17726 5794 17778
rect 6526 17726 6578 17778
rect 7086 17726 7138 17778
rect 7870 17726 7922 17778
rect 8430 17726 8482 17778
rect 14142 17726 14194 17778
rect 19630 17726 19682 17778
rect 19966 17726 20018 17778
rect 20526 17726 20578 17778
rect 20974 17726 21026 17778
rect 23774 17726 23826 17778
rect 24894 17726 24946 17778
rect 25342 17726 25394 17778
rect 26574 17726 26626 17778
rect 27582 17726 27634 17778
rect 28590 17726 28642 17778
rect 38894 17726 38946 17778
rect 40910 17726 40962 17778
rect 41358 17726 41410 17778
rect 43822 17726 43874 17778
rect 44494 17726 44546 17778
rect 46622 17726 46674 17778
rect 49982 17726 50034 17778
rect 51326 17726 51378 17778
rect 53454 17726 53506 17778
rect 53790 17726 53842 17778
rect 9550 17614 9602 17666
rect 9886 17614 9938 17666
rect 13582 17614 13634 17666
rect 15486 17614 15538 17666
rect 16158 17614 16210 17666
rect 19182 17614 19234 17666
rect 22094 17614 22146 17666
rect 22542 17614 22594 17666
rect 23102 17614 23154 17666
rect 24446 17614 24498 17666
rect 25678 17614 25730 17666
rect 26350 17614 26402 17666
rect 26686 17614 26738 17666
rect 33406 17614 33458 17666
rect 34190 17614 34242 17666
rect 34526 17614 34578 17666
rect 35870 17614 35922 17666
rect 36094 17614 36146 17666
rect 36318 17614 36370 17666
rect 38782 17614 38834 17666
rect 40238 17614 40290 17666
rect 42590 17614 42642 17666
rect 42814 17614 42866 17666
rect 43710 17614 43762 17666
rect 46510 17614 46562 17666
rect 48862 17614 48914 17666
rect 51438 17614 51490 17666
rect 51998 17614 52050 17666
rect 55470 17614 55522 17666
rect 57038 17614 57090 17666
rect 57374 17614 57426 17666
rect 25902 17502 25954 17554
rect 27022 17502 27074 17554
rect 30046 17502 30098 17554
rect 30606 17502 30658 17554
rect 32286 17502 32338 17554
rect 32734 17502 32786 17554
rect 35086 17502 35138 17554
rect 35646 17502 35698 17554
rect 36766 17502 36818 17554
rect 39678 17502 39730 17554
rect 42926 17502 42978 17554
rect 47406 17502 47458 17554
rect 48974 17502 49026 17554
rect 55694 17502 55746 17554
rect 6078 17390 6130 17442
rect 7422 17390 7474 17442
rect 8990 17390 9042 17442
rect 12238 17390 12290 17442
rect 14590 17390 14642 17442
rect 15038 17390 15090 17442
rect 18510 17390 18562 17442
rect 21870 17390 21922 17442
rect 21982 17390 22034 17442
rect 28142 17390 28194 17442
rect 28702 17390 28754 17442
rect 31166 17390 31218 17442
rect 35982 17390 36034 17442
rect 37886 17390 37938 17442
rect 40350 17390 40402 17442
rect 40574 17390 40626 17442
rect 56926 17390 56978 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 4622 17054 4674 17106
rect 5070 17054 5122 17106
rect 8542 17054 8594 17106
rect 9102 17054 9154 17106
rect 9774 17054 9826 17106
rect 10222 17054 10274 17106
rect 10670 17054 10722 17106
rect 12126 17054 12178 17106
rect 15710 17054 15762 17106
rect 16158 17054 16210 17106
rect 16606 17054 16658 17106
rect 17726 17054 17778 17106
rect 18062 17054 18114 17106
rect 19182 17054 19234 17106
rect 19854 17054 19906 17106
rect 20526 17054 20578 17106
rect 20974 17054 21026 17106
rect 21422 17054 21474 17106
rect 22990 17054 23042 17106
rect 23550 17054 23602 17106
rect 23998 17054 24050 17106
rect 25006 17054 25058 17106
rect 26238 17054 26290 17106
rect 28366 17054 28418 17106
rect 29374 17054 29426 17106
rect 29934 17054 29986 17106
rect 30046 17054 30098 17106
rect 31054 17054 31106 17106
rect 31390 17054 31442 17106
rect 31838 17054 31890 17106
rect 32734 17054 32786 17106
rect 33854 17054 33906 17106
rect 34078 17054 34130 17106
rect 34750 17054 34802 17106
rect 38894 17054 38946 17106
rect 39566 17054 39618 17106
rect 40350 17054 40402 17106
rect 40574 17054 40626 17106
rect 41470 17054 41522 17106
rect 41918 17054 41970 17106
rect 43038 17054 43090 17106
rect 43150 17054 43202 17106
rect 43262 17054 43314 17106
rect 44382 17054 44434 17106
rect 45166 17054 45218 17106
rect 45614 17054 45666 17106
rect 53790 17054 53842 17106
rect 58270 17054 58322 17106
rect 17054 16942 17106 16994
rect 18846 16942 18898 16994
rect 21870 16942 21922 16994
rect 22206 16942 22258 16994
rect 24446 16942 24498 16994
rect 32622 16942 32674 16994
rect 34190 16942 34242 16994
rect 35646 16942 35698 16994
rect 36542 16942 36594 16994
rect 38334 16942 38386 16994
rect 40126 16942 40178 16994
rect 44718 16942 44770 16994
rect 53902 16942 53954 16994
rect 56366 16942 56418 16994
rect 57822 16942 57874 16994
rect 58158 16942 58210 16994
rect 58382 16942 58434 16994
rect 5406 16830 5458 16882
rect 5966 16830 6018 16882
rect 11230 16830 11282 16882
rect 14478 16830 14530 16882
rect 15038 16830 15090 16882
rect 26686 16830 26738 16882
rect 27246 16830 27298 16882
rect 28702 16830 28754 16882
rect 30158 16830 30210 16882
rect 30606 16830 30658 16882
rect 32958 16830 33010 16882
rect 33742 16830 33794 16882
rect 35310 16830 35362 16882
rect 35534 16830 35586 16882
rect 37438 16830 37490 16882
rect 37886 16830 37938 16882
rect 42814 16830 42866 16882
rect 42926 16830 42978 16882
rect 43822 16830 43874 16882
rect 50094 16830 50146 16882
rect 51998 16830 52050 16882
rect 52334 16830 52386 16882
rect 53342 16830 53394 16882
rect 54014 16830 54066 16882
rect 55246 16830 55298 16882
rect 55582 16830 55634 16882
rect 56254 16830 56306 16882
rect 25678 16718 25730 16770
rect 27470 16718 27522 16770
rect 30606 16718 30658 16770
rect 34190 16718 34242 16770
rect 50318 16718 50370 16770
rect 50766 16718 50818 16770
rect 10334 16606 10386 16658
rect 10894 16606 10946 16658
rect 18958 16606 19010 16658
rect 19518 16606 19570 16658
rect 28366 16606 28418 16658
rect 28478 16606 28530 16658
rect 52894 16718 52946 16770
rect 55918 16718 55970 16770
rect 31278 16606 31330 16658
rect 36094 16606 36146 16658
rect 40686 16606 40738 16658
rect 57486 16606 57538 16658
rect 57598 16606 57650 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 11790 16270 11842 16322
rect 13582 16270 13634 16322
rect 14366 16270 14418 16322
rect 19070 16270 19122 16322
rect 27582 16270 27634 16322
rect 27806 16270 27858 16322
rect 28366 16270 28418 16322
rect 29710 16270 29762 16322
rect 30606 16270 30658 16322
rect 31278 16270 31330 16322
rect 42814 16270 42866 16322
rect 45726 16270 45778 16322
rect 6414 16158 6466 16210
rect 7646 16158 7698 16210
rect 12574 16158 12626 16210
rect 13022 16158 13074 16210
rect 14590 16158 14642 16210
rect 19518 16158 19570 16210
rect 19854 16158 19906 16210
rect 20414 16158 20466 16210
rect 20862 16158 20914 16210
rect 21646 16158 21698 16210
rect 22318 16158 22370 16210
rect 23214 16158 23266 16210
rect 23662 16158 23714 16210
rect 24894 16158 24946 16210
rect 26238 16158 26290 16210
rect 27470 16158 27522 16210
rect 28254 16158 28306 16210
rect 29598 16158 29650 16210
rect 31838 16158 31890 16210
rect 32286 16158 32338 16210
rect 32734 16158 32786 16210
rect 33182 16158 33234 16210
rect 34750 16158 34802 16210
rect 37438 16158 37490 16210
rect 37886 16158 37938 16210
rect 38446 16158 38498 16210
rect 41246 16158 41298 16210
rect 41694 16158 41746 16210
rect 42142 16158 42194 16210
rect 46062 16158 46114 16210
rect 46622 16158 46674 16210
rect 53678 16158 53730 16210
rect 55918 16158 55970 16210
rect 8094 16046 8146 16098
rect 8766 16046 8818 16098
rect 15374 16046 15426 16098
rect 16046 16046 16098 16098
rect 22430 16046 22482 16098
rect 26014 16046 26066 16098
rect 31166 16046 31218 16098
rect 34078 16046 34130 16098
rect 35982 16046 36034 16098
rect 39006 16046 39058 16098
rect 40238 16046 40290 16098
rect 40686 16046 40738 16098
rect 43374 16046 43426 16098
rect 43710 16046 43762 16098
rect 52782 16046 52834 16098
rect 55022 16046 55074 16098
rect 56142 16046 56194 16098
rect 58494 16046 58546 16098
rect 18286 15934 18338 15986
rect 22206 15934 22258 15986
rect 22766 15934 22818 15986
rect 25342 15934 25394 15986
rect 27358 15934 27410 15986
rect 30382 15934 30434 15986
rect 31278 15934 31330 15986
rect 34190 15934 34242 15986
rect 35422 15934 35474 15986
rect 35646 15934 35698 15986
rect 36430 15934 36482 15986
rect 39118 15934 39170 15986
rect 39790 15934 39842 15986
rect 42702 15934 42754 15986
rect 42814 15934 42866 15986
rect 44046 15934 44098 15986
rect 44606 15934 44658 15986
rect 45950 15934 46002 15986
rect 52446 15934 52498 15986
rect 53454 15934 53506 15986
rect 55246 15934 55298 15986
rect 57822 15934 57874 15986
rect 5854 15822 5906 15874
rect 6750 15822 6802 15874
rect 7198 15822 7250 15874
rect 11118 15822 11170 15874
rect 13582 15822 13634 15874
rect 14030 15822 14082 15874
rect 15038 15822 15090 15874
rect 24446 15822 24498 15874
rect 28590 15822 28642 15874
rect 30494 15822 30546 15874
rect 34414 15822 34466 15874
rect 35870 15822 35922 15874
rect 39342 15822 39394 15874
rect 43710 15822 43762 15874
rect 46734 15822 46786 15874
rect 49198 15822 49250 15874
rect 52558 15822 52610 15874
rect 53678 15822 53730 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 10558 15486 10610 15538
rect 11006 15486 11058 15538
rect 18062 15486 18114 15538
rect 19742 15486 19794 15538
rect 24558 15486 24610 15538
rect 26238 15486 26290 15538
rect 26574 15486 26626 15538
rect 27022 15486 27074 15538
rect 28030 15486 28082 15538
rect 28478 15486 28530 15538
rect 28926 15486 28978 15538
rect 29374 15486 29426 15538
rect 30718 15486 30770 15538
rect 31390 15486 31442 15538
rect 32286 15486 32338 15538
rect 33630 15486 33682 15538
rect 34526 15486 34578 15538
rect 35198 15486 35250 15538
rect 38894 15486 38946 15538
rect 42926 15486 42978 15538
rect 43934 15486 43986 15538
rect 45838 15486 45890 15538
rect 48638 15486 48690 15538
rect 49758 15486 49810 15538
rect 55694 15486 55746 15538
rect 5406 15374 5458 15426
rect 16606 15374 16658 15426
rect 17614 15374 17666 15426
rect 22206 15374 22258 15426
rect 23886 15374 23938 15426
rect 24894 15374 24946 15426
rect 31614 15374 31666 15426
rect 37438 15374 37490 15426
rect 37998 15374 38050 15426
rect 39230 15374 39282 15426
rect 40798 15374 40850 15426
rect 41806 15374 41858 15426
rect 42366 15374 42418 15426
rect 43710 15374 43762 15426
rect 45054 15374 45106 15426
rect 45614 15374 45666 15426
rect 45950 15374 46002 15426
rect 46174 15374 46226 15426
rect 47182 15374 47234 15426
rect 49982 15374 50034 15426
rect 52558 15374 52610 15426
rect 56366 15374 56418 15426
rect 57486 15374 57538 15426
rect 8318 15262 8370 15314
rect 11790 15262 11842 15314
rect 18510 15262 18562 15314
rect 21198 15262 21250 15314
rect 21422 15262 21474 15314
rect 22878 15262 22930 15314
rect 23774 15262 23826 15314
rect 25678 15262 25730 15314
rect 27470 15262 27522 15314
rect 30494 15262 30546 15314
rect 30606 15262 30658 15314
rect 30830 15262 30882 15314
rect 31726 15262 31778 15314
rect 33966 15262 34018 15314
rect 35870 15262 35922 15314
rect 35982 15262 36034 15314
rect 36206 15262 36258 15314
rect 36766 15262 36818 15314
rect 37214 15262 37266 15314
rect 38334 15262 38386 15314
rect 39902 15262 39954 15314
rect 40350 15262 40402 15314
rect 42590 15262 42642 15314
rect 43486 15262 43538 15314
rect 49534 15262 49586 15314
rect 49646 15262 49698 15314
rect 52446 15262 52498 15314
rect 52670 15262 52722 15314
rect 53342 15262 53394 15314
rect 54238 15262 54290 15314
rect 54798 15262 54850 15314
rect 55582 15262 55634 15314
rect 56702 15262 56754 15314
rect 57598 15262 57650 15314
rect 57934 15262 57986 15314
rect 9662 15150 9714 15202
rect 19294 15150 19346 15202
rect 21646 15150 21698 15202
rect 22990 15150 23042 15202
rect 32622 15150 32674 15202
rect 37326 15150 37378 15202
rect 43598 15150 43650 15202
rect 47294 15150 47346 15202
rect 48414 15150 48466 15202
rect 30158 15038 30210 15090
rect 36318 15038 36370 15090
rect 38334 15038 38386 15090
rect 46958 15038 47010 15090
rect 48750 15038 48802 15090
rect 54462 15038 54514 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 7198 14702 7250 14754
rect 8206 14702 8258 14754
rect 13022 14702 13074 14754
rect 19070 14702 19122 14754
rect 27694 14702 27746 14754
rect 30158 14702 30210 14754
rect 30606 14702 30658 14754
rect 31614 14702 31666 14754
rect 33854 14702 33906 14754
rect 35086 14702 35138 14754
rect 35422 14702 35474 14754
rect 35646 14702 35698 14754
rect 36430 14702 36482 14754
rect 43150 14702 43202 14754
rect 43486 14702 43538 14754
rect 51886 14702 51938 14754
rect 52222 14702 52274 14754
rect 4958 14590 5010 14642
rect 5630 14590 5682 14642
rect 6414 14590 6466 14642
rect 6862 14590 6914 14642
rect 7310 14590 7362 14642
rect 7758 14590 7810 14642
rect 8766 14590 8818 14642
rect 13694 14590 13746 14642
rect 14030 14590 14082 14642
rect 22766 14590 22818 14642
rect 23886 14590 23938 14642
rect 26574 14590 26626 14642
rect 31054 14590 31106 14642
rect 31390 14590 31442 14642
rect 35982 14590 36034 14642
rect 36766 14590 36818 14642
rect 43150 14590 43202 14642
rect 44270 14590 44322 14642
rect 44718 14590 44770 14642
rect 46510 14590 46562 14642
rect 48862 14590 48914 14642
rect 49646 14590 49698 14642
rect 50318 14590 50370 14642
rect 54686 14590 54738 14642
rect 55582 14590 55634 14642
rect 56478 14590 56530 14642
rect 57262 14590 57314 14642
rect 9550 14478 9602 14530
rect 9998 14478 10050 14530
rect 15374 14478 15426 14530
rect 16046 14478 16098 14530
rect 21870 14478 21922 14530
rect 25118 14478 25170 14530
rect 27134 14478 27186 14530
rect 30494 14478 30546 14530
rect 32510 14478 32562 14530
rect 32734 14478 32786 14530
rect 34078 14478 34130 14530
rect 34526 14478 34578 14530
rect 38334 14478 38386 14530
rect 44046 14478 44098 14530
rect 46846 14478 46898 14530
rect 49982 14478 50034 14530
rect 51662 14478 51714 14530
rect 54238 14478 54290 14530
rect 54462 14478 54514 14530
rect 56254 14478 56306 14530
rect 18286 14366 18338 14418
rect 22766 14366 22818 14418
rect 22990 14366 23042 14418
rect 27582 14366 27634 14418
rect 29710 14366 29762 14418
rect 29934 14366 29986 14418
rect 35310 14366 35362 14418
rect 36318 14366 36370 14418
rect 38110 14366 38162 14418
rect 39566 14366 39618 14418
rect 47406 14366 47458 14418
rect 8206 14254 8258 14306
rect 12462 14254 12514 14306
rect 14478 14254 14530 14306
rect 14926 14254 14978 14306
rect 19406 14254 19458 14306
rect 21646 14254 21698 14306
rect 24222 14254 24274 14306
rect 24782 14254 24834 14306
rect 25902 14254 25954 14306
rect 26462 14254 26514 14306
rect 26686 14254 26738 14306
rect 27694 14254 27746 14306
rect 28366 14254 28418 14306
rect 28814 14254 28866 14306
rect 30046 14254 30098 14306
rect 31838 14254 31890 14306
rect 32846 14254 32898 14306
rect 32958 14254 33010 14306
rect 33070 14254 33122 14306
rect 39678 14254 39730 14306
rect 42030 14254 42082 14306
rect 47854 14254 47906 14306
rect 58494 14254 58546 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 8094 13918 8146 13970
rect 8878 13918 8930 13970
rect 9662 13918 9714 13970
rect 10110 13918 10162 13970
rect 13694 13918 13746 13970
rect 22542 13918 22594 13970
rect 23438 13918 23490 13970
rect 28590 13918 28642 13970
rect 29150 13918 29202 13970
rect 29598 13918 29650 13970
rect 31502 13918 31554 13970
rect 39790 13918 39842 13970
rect 44158 13918 44210 13970
rect 46062 13918 46114 13970
rect 48190 13918 48242 13970
rect 55358 13918 55410 13970
rect 55806 13918 55858 13970
rect 30830 13806 30882 13858
rect 34302 13806 34354 13858
rect 34638 13806 34690 13858
rect 35422 13806 35474 13858
rect 37774 13806 37826 13858
rect 37998 13806 38050 13858
rect 38334 13806 38386 13858
rect 42702 13806 42754 13858
rect 43038 13806 43090 13858
rect 46622 13806 46674 13858
rect 46846 13806 46898 13858
rect 47630 13806 47682 13858
rect 47742 13806 47794 13858
rect 52670 13806 52722 13858
rect 53790 13806 53842 13858
rect 4286 13694 4338 13746
rect 5406 13694 5458 13746
rect 5742 13694 5794 13746
rect 10558 13694 10610 13746
rect 11230 13694 11282 13746
rect 16270 13694 16322 13746
rect 22430 13694 22482 13746
rect 22654 13694 22706 13746
rect 23102 13694 23154 13746
rect 24334 13694 24386 13746
rect 26126 13694 26178 13746
rect 27694 13694 27746 13746
rect 32174 13694 32226 13746
rect 32398 13694 32450 13746
rect 32622 13694 32674 13746
rect 32846 13694 32898 13746
rect 33742 13694 33794 13746
rect 43262 13694 43314 13746
rect 47406 13694 47458 13746
rect 3950 13582 4002 13634
rect 14926 13582 14978 13634
rect 15374 13582 15426 13634
rect 15822 13582 15874 13634
rect 19182 13582 19234 13634
rect 19742 13582 19794 13634
rect 24894 13582 24946 13634
rect 26462 13582 26514 13634
rect 30046 13582 30098 13634
rect 32510 13582 32562 13634
rect 34078 13582 34130 13634
rect 38222 13582 38274 13634
rect 41470 13582 41522 13634
rect 45614 13582 45666 13634
rect 51998 13582 52050 13634
rect 4286 13470 4338 13522
rect 14254 13470 14306 13522
rect 27582 13470 27634 13522
rect 29710 13470 29762 13522
rect 29934 13470 29986 13522
rect 30942 13470 30994 13522
rect 43598 13470 43650 13522
rect 46958 13470 47010 13522
rect 54798 13470 54850 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 10222 13134 10274 13186
rect 19070 13134 19122 13186
rect 26574 13134 26626 13186
rect 30046 13134 30098 13186
rect 52334 13134 52386 13186
rect 52670 13134 52722 13186
rect 10894 13022 10946 13074
rect 11342 13022 11394 13074
rect 12350 13022 12402 13074
rect 13582 13022 13634 13074
rect 14590 13022 14642 13074
rect 19630 13022 19682 13074
rect 23662 13022 23714 13074
rect 25454 13022 25506 13074
rect 26462 13022 26514 13074
rect 28030 13022 28082 13074
rect 31166 13022 31218 13074
rect 31726 13022 31778 13074
rect 32174 13022 32226 13074
rect 32734 13022 32786 13074
rect 33742 13022 33794 13074
rect 34974 13022 35026 13074
rect 37662 13022 37714 13074
rect 38894 13022 38946 13074
rect 41918 13022 41970 13074
rect 43822 13022 43874 13074
rect 45726 13022 45778 13074
rect 46622 13022 46674 13074
rect 49310 13022 49362 13074
rect 51214 13022 51266 13074
rect 52110 13022 52162 13074
rect 3838 12910 3890 12962
rect 5630 12910 5682 12962
rect 6190 12910 6242 12962
rect 10446 12910 10498 12962
rect 11902 12910 11954 12962
rect 12910 12910 12962 12962
rect 15374 12910 15426 12962
rect 16046 12910 16098 12962
rect 20526 12910 20578 12962
rect 22318 12910 22370 12962
rect 27470 12910 27522 12962
rect 29710 12910 29762 12962
rect 29822 12910 29874 12962
rect 31390 12910 31442 12962
rect 33518 12910 33570 12962
rect 37774 12910 37826 12962
rect 40126 12910 40178 12962
rect 40798 12910 40850 12962
rect 41246 12910 41298 12962
rect 43150 12910 43202 12962
rect 43598 12910 43650 12962
rect 46398 12910 46450 12962
rect 47742 12910 47794 12962
rect 49758 12910 49810 12962
rect 50990 12910 51042 12962
rect 56478 12910 56530 12962
rect 3502 12798 3554 12850
rect 4286 12798 4338 12850
rect 4734 12798 4786 12850
rect 9886 12798 9938 12850
rect 18286 12798 18338 12850
rect 23214 12798 23266 12850
rect 24782 12798 24834 12850
rect 26350 12798 26402 12850
rect 30158 12798 30210 12850
rect 30718 12798 30770 12850
rect 30942 12798 30994 12850
rect 34414 12798 34466 12850
rect 37550 12798 37602 12850
rect 39566 12798 39618 12850
rect 41358 12798 41410 12850
rect 48526 12798 48578 12850
rect 50206 12798 50258 12850
rect 50766 12798 50818 12850
rect 51326 12798 51378 12850
rect 3614 12686 3666 12738
rect 4510 12686 4562 12738
rect 4846 12686 4898 12738
rect 8766 12686 8818 12738
rect 9326 12686 9378 12738
rect 14142 12686 14194 12738
rect 21758 12686 21810 12738
rect 24334 12686 24386 12738
rect 27134 12686 27186 12738
rect 28366 12686 28418 12738
rect 28814 12686 28866 12738
rect 37998 12686 38050 12738
rect 38446 12686 38498 12738
rect 39454 12686 39506 12738
rect 40238 12686 40290 12738
rect 40350 12686 40402 12738
rect 41582 12686 41634 12738
rect 56254 12686 56306 12738
rect 56366 12686 56418 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 6190 12350 6242 12402
rect 9662 12350 9714 12402
rect 10110 12350 10162 12402
rect 10670 12350 10722 12402
rect 20190 12350 20242 12402
rect 22654 12350 22706 12402
rect 22766 12350 22818 12402
rect 23326 12350 23378 12402
rect 23550 12350 23602 12402
rect 26014 12350 26066 12402
rect 27246 12350 27298 12402
rect 28030 12350 28082 12402
rect 28702 12350 28754 12402
rect 31950 12350 32002 12402
rect 32398 12350 32450 12402
rect 32958 12350 33010 12402
rect 33518 12350 33570 12402
rect 33966 12350 34018 12402
rect 35422 12350 35474 12402
rect 40462 12350 40514 12402
rect 42030 12350 42082 12402
rect 43038 12350 43090 12402
rect 43486 12350 43538 12402
rect 43934 12350 43986 12402
rect 45950 12350 46002 12402
rect 47630 12350 47682 12402
rect 49646 12350 49698 12402
rect 49758 12350 49810 12402
rect 56590 12350 56642 12402
rect 15150 12238 15202 12290
rect 21422 12238 21474 12290
rect 21758 12238 21810 12290
rect 22878 12238 22930 12290
rect 23662 12238 23714 12290
rect 24334 12238 24386 12290
rect 30494 12238 30546 12290
rect 31054 12238 31106 12290
rect 34974 12238 35026 12290
rect 36878 12238 36930 12290
rect 36990 12238 37042 12290
rect 38894 12238 38946 12290
rect 39454 12238 39506 12290
rect 41806 12238 41858 12290
rect 42590 12238 42642 12290
rect 47182 12238 47234 12290
rect 47406 12238 47458 12290
rect 47742 12238 47794 12290
rect 49534 12238 49586 12290
rect 53902 12238 53954 12290
rect 56030 12238 56082 12290
rect 57598 12238 57650 12290
rect 4174 12126 4226 12178
rect 5406 12126 5458 12178
rect 8430 12126 8482 12178
rect 9102 12126 9154 12178
rect 11230 12126 11282 12178
rect 11678 12126 11730 12178
rect 18734 12126 18786 12178
rect 28814 12126 28866 12178
rect 29598 12126 29650 12178
rect 30046 12126 30098 12178
rect 31278 12126 31330 12178
rect 34638 12126 34690 12178
rect 36654 12126 36706 12178
rect 37326 12126 37378 12178
rect 39230 12126 39282 12178
rect 40238 12126 40290 12178
rect 40686 12126 40738 12178
rect 41582 12126 41634 12178
rect 55582 12126 55634 12178
rect 56478 12126 56530 12178
rect 57374 12126 57426 12178
rect 57710 12126 57762 12178
rect 4286 12014 4338 12066
rect 4622 12014 4674 12066
rect 19182 12014 19234 12066
rect 24446 12014 24498 12066
rect 26462 12014 26514 12066
rect 27582 12014 27634 12066
rect 37438 12014 37490 12066
rect 37886 12014 37938 12066
rect 38334 12014 38386 12066
rect 39006 12014 39058 12066
rect 40574 12014 40626 12066
rect 41694 12014 41746 12066
rect 45166 12014 45218 12066
rect 28926 11902 28978 11954
rect 32286 11902 32338 11954
rect 32846 11902 32898 11954
rect 33854 11902 33906 11954
rect 34414 11902 34466 11954
rect 34638 11902 34690 11954
rect 40014 11902 40066 11954
rect 53678 11902 53730 11954
rect 54014 11902 54066 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 10894 11566 10946 11618
rect 11678 11566 11730 11618
rect 24670 11566 24722 11618
rect 26574 11566 26626 11618
rect 33518 11566 33570 11618
rect 35310 11566 35362 11618
rect 41246 11566 41298 11618
rect 41470 11566 41522 11618
rect 41806 11566 41858 11618
rect 42814 11566 42866 11618
rect 5070 11454 5122 11506
rect 8094 11454 8146 11506
rect 10558 11454 10610 11506
rect 11118 11454 11170 11506
rect 11678 11454 11730 11506
rect 19070 11454 19122 11506
rect 19630 11454 19682 11506
rect 21646 11454 21698 11506
rect 22318 11454 22370 11506
rect 23214 11454 23266 11506
rect 28366 11454 28418 11506
rect 30606 11454 30658 11506
rect 32958 11454 33010 11506
rect 39006 11454 39058 11506
rect 41134 11454 41186 11506
rect 41806 11454 41858 11506
rect 42142 11454 42194 11506
rect 45502 11454 45554 11506
rect 51326 11454 51378 11506
rect 56478 11454 56530 11506
rect 5742 11342 5794 11394
rect 6638 11342 6690 11394
rect 8990 11342 9042 11394
rect 10334 11342 10386 11394
rect 15486 11342 15538 11394
rect 16046 11342 16098 11394
rect 22094 11342 22146 11394
rect 22430 11342 22482 11394
rect 25342 11342 25394 11394
rect 27470 11342 27522 11394
rect 30158 11342 30210 11394
rect 30494 11342 30546 11394
rect 33854 11342 33906 11394
rect 34190 11342 34242 11394
rect 38782 11342 38834 11394
rect 40462 11342 40514 11394
rect 44046 11342 44098 11394
rect 44606 11342 44658 11394
rect 45726 11342 45778 11394
rect 50990 11342 51042 11394
rect 54014 11342 54066 11394
rect 54910 11342 54962 11394
rect 55358 11342 55410 11394
rect 57038 11342 57090 11394
rect 6078 11230 6130 11282
rect 6974 11230 7026 11282
rect 8542 11230 8594 11282
rect 9662 11230 9714 11282
rect 18286 11230 18338 11282
rect 22766 11230 22818 11282
rect 25902 11230 25954 11282
rect 26014 11230 26066 11282
rect 26126 11230 26178 11282
rect 27134 11230 27186 11282
rect 32174 11230 32226 11282
rect 35646 11230 35698 11282
rect 35870 11230 35922 11282
rect 38110 11230 38162 11282
rect 40126 11230 40178 11282
rect 43038 11230 43090 11282
rect 44718 11230 44770 11282
rect 47070 11230 47122 11282
rect 51662 11230 51714 11282
rect 54126 11230 54178 11282
rect 54686 11230 54738 11282
rect 56590 11230 56642 11282
rect 14926 11118 14978 11170
rect 24222 11118 24274 11170
rect 24782 11118 24834 11170
rect 25006 11118 25058 11170
rect 27246 11118 27298 11170
rect 27806 11118 27858 11170
rect 28926 11118 28978 11170
rect 31054 11118 31106 11170
rect 33966 11118 34018 11170
rect 34078 11118 34130 11170
rect 34974 11118 35026 11170
rect 40350 11118 40402 11170
rect 42926 11118 42978 11170
rect 46062 11118 46114 11170
rect 46622 11118 46674 11170
rect 46734 11118 46786 11170
rect 46846 11118 46898 11170
rect 56366 11118 56418 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 9102 10782 9154 10834
rect 16494 10782 16546 10834
rect 17054 10782 17106 10834
rect 18062 10782 18114 10834
rect 24446 10782 24498 10834
rect 25566 10782 25618 10834
rect 25678 10782 25730 10834
rect 25902 10782 25954 10834
rect 29262 10782 29314 10834
rect 29710 10782 29762 10834
rect 31502 10782 31554 10834
rect 33630 10782 33682 10834
rect 39342 10782 39394 10834
rect 39790 10782 39842 10834
rect 40686 10782 40738 10834
rect 41582 10782 41634 10834
rect 42366 10782 42418 10834
rect 42702 10782 42754 10834
rect 44158 10782 44210 10834
rect 48750 10782 48802 10834
rect 49758 10782 49810 10834
rect 9998 10670 10050 10722
rect 10334 10670 10386 10722
rect 19630 10670 19682 10722
rect 22094 10670 22146 10722
rect 23774 10670 23826 10722
rect 26126 10670 26178 10722
rect 26798 10670 26850 10722
rect 32622 10670 32674 10722
rect 34302 10670 34354 10722
rect 43710 10670 43762 10722
rect 43934 10670 43986 10722
rect 49534 10670 49586 10722
rect 55806 10670 55858 10722
rect 4846 10558 4898 10610
rect 13582 10558 13634 10610
rect 14030 10558 14082 10610
rect 17614 10558 17666 10610
rect 19966 10558 20018 10610
rect 20526 10558 20578 10610
rect 21198 10558 21250 10610
rect 22654 10558 22706 10610
rect 23662 10558 23714 10610
rect 24670 10558 24722 10610
rect 25006 10558 25058 10610
rect 31390 10558 31442 10610
rect 31614 10558 31666 10610
rect 32062 10558 32114 10610
rect 32510 10558 32562 10610
rect 35086 10558 35138 10610
rect 35310 10558 35362 10610
rect 36542 10558 36594 10610
rect 37550 10558 37602 10610
rect 37774 10558 37826 10610
rect 44270 10558 44322 10610
rect 44718 10558 44770 10610
rect 46622 10558 46674 10610
rect 47406 10558 47458 10610
rect 50990 10558 51042 10610
rect 51326 10558 51378 10610
rect 53118 10558 53170 10610
rect 53342 10558 53394 10610
rect 54798 10558 54850 10610
rect 55694 10558 55746 10610
rect 56030 10558 56082 10610
rect 5070 10446 5122 10498
rect 18510 10446 18562 10498
rect 21422 10446 21474 10498
rect 22990 10446 23042 10498
rect 24334 10446 24386 10498
rect 26686 10446 26738 10498
rect 27470 10446 27522 10498
rect 27918 10446 27970 10498
rect 28478 10446 28530 10498
rect 28814 10446 28866 10498
rect 30158 10446 30210 10498
rect 30718 10446 30770 10498
rect 35982 10446 36034 10498
rect 40238 10446 40290 10498
rect 43150 10446 43202 10498
rect 45166 10446 45218 10498
rect 45614 10446 45666 10498
rect 47070 10446 47122 10498
rect 51550 10446 51602 10498
rect 54014 10446 54066 10498
rect 54574 10446 54626 10498
rect 5294 10334 5346 10386
rect 27022 10334 27074 10386
rect 32622 10334 32674 10386
rect 34078 10334 34130 10386
rect 34414 10334 34466 10386
rect 38110 10334 38162 10386
rect 39230 10334 39282 10386
rect 40238 10334 40290 10386
rect 49870 10334 49922 10386
rect 55134 10334 55186 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 13022 9998 13074 10050
rect 22990 9998 23042 10050
rect 26350 9998 26402 10050
rect 26686 9998 26738 10050
rect 27358 9998 27410 10050
rect 29710 9998 29762 10050
rect 38894 9998 38946 10050
rect 44270 9998 44322 10050
rect 46286 9998 46338 10050
rect 46622 9998 46674 10050
rect 55470 9998 55522 10050
rect 8430 9886 8482 9938
rect 14030 9886 14082 9938
rect 19294 9886 19346 9938
rect 22766 9886 22818 9938
rect 23550 9886 23602 9938
rect 28590 9886 28642 9938
rect 33518 9886 33570 9938
rect 43262 9886 43314 9938
rect 48302 9886 48354 9938
rect 49422 9886 49474 9938
rect 51662 9886 51714 9938
rect 56814 9886 56866 9938
rect 57486 9886 57538 9938
rect 4286 9774 4338 9826
rect 4846 9774 4898 9826
rect 9550 9774 9602 9826
rect 9886 9774 9938 9826
rect 15486 9774 15538 9826
rect 15934 9774 15986 9826
rect 22654 9774 22706 9826
rect 25790 9774 25842 9826
rect 26910 9774 26962 9826
rect 28030 9774 28082 9826
rect 29598 9774 29650 9826
rect 31502 9774 31554 9826
rect 32174 9774 32226 9826
rect 34750 9774 34802 9826
rect 35086 9774 35138 9826
rect 35310 9774 35362 9826
rect 37886 9774 37938 9826
rect 37998 9774 38050 9826
rect 39230 9774 39282 9826
rect 40014 9774 40066 9826
rect 40462 9774 40514 9826
rect 40910 9774 40962 9826
rect 41134 9774 41186 9826
rect 42030 9774 42082 9826
rect 43038 9774 43090 9826
rect 44606 9774 44658 9826
rect 46622 9774 46674 9826
rect 47070 9774 47122 9826
rect 49198 9774 49250 9826
rect 54350 9774 54402 9826
rect 54574 9774 54626 9826
rect 55246 9774 55298 9826
rect 56926 9774 56978 9826
rect 4958 9662 5010 9714
rect 5742 9662 5794 9714
rect 18958 9662 19010 9714
rect 27694 9662 27746 9714
rect 28478 9662 28530 9714
rect 30942 9662 30994 9714
rect 34078 9662 34130 9714
rect 34974 9662 35026 9714
rect 37550 9662 37602 9714
rect 41694 9662 41746 9714
rect 43710 9662 43762 9714
rect 49870 9662 49922 9714
rect 6078 9550 6130 9602
rect 8878 9550 8930 9602
rect 12462 9550 12514 9602
rect 13582 9550 13634 9602
rect 14814 9550 14866 9602
rect 18398 9550 18450 9602
rect 25118 9550 25170 9602
rect 27470 9550 27522 9602
rect 28702 9550 28754 9602
rect 29710 9550 29762 9602
rect 32734 9550 32786 9602
rect 37774 9550 37826 9602
rect 39006 9550 39058 9602
rect 40798 9550 40850 9602
rect 41806 9550 41858 9602
rect 44382 9550 44434 9602
rect 45390 9550 45442 9602
rect 51550 9550 51602 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 4398 9214 4450 9266
rect 4846 9214 4898 9266
rect 8318 9214 8370 9266
rect 8990 9214 9042 9266
rect 13022 9214 13074 9266
rect 14030 9214 14082 9266
rect 21310 9214 21362 9266
rect 21870 9214 21922 9266
rect 22654 9214 22706 9266
rect 23550 9214 23602 9266
rect 25678 9214 25730 9266
rect 26238 9214 26290 9266
rect 26686 9214 26738 9266
rect 27134 9214 27186 9266
rect 31054 9214 31106 9266
rect 31726 9214 31778 9266
rect 33742 9214 33794 9266
rect 34638 9214 34690 9266
rect 34974 9214 35026 9266
rect 35646 9214 35698 9266
rect 36318 9214 36370 9266
rect 42030 9214 42082 9266
rect 42254 9214 42306 9266
rect 43150 9214 43202 9266
rect 45502 9214 45554 9266
rect 54686 9214 54738 9266
rect 57598 9214 57650 9266
rect 10110 9102 10162 9154
rect 11006 9102 11058 9154
rect 22990 9102 23042 9154
rect 31614 9102 31666 9154
rect 32398 9102 32450 9154
rect 32734 9102 32786 9154
rect 36206 9102 36258 9154
rect 39118 9102 39170 9154
rect 41918 9102 41970 9154
rect 42702 9102 42754 9154
rect 43822 9102 43874 9154
rect 44494 9102 44546 9154
rect 44718 9102 44770 9154
rect 44942 9102 44994 9154
rect 45054 9102 45106 9154
rect 46286 9102 46338 9154
rect 46510 9102 46562 9154
rect 47406 9102 47458 9154
rect 47630 9102 47682 9154
rect 49534 9102 49586 9154
rect 49758 9102 49810 9154
rect 50430 9102 50482 9154
rect 51662 9102 51714 9154
rect 53678 9102 53730 9154
rect 54462 9102 54514 9154
rect 54798 9102 54850 9154
rect 57486 9102 57538 9154
rect 57710 9102 57762 9154
rect 4286 8990 4338 9042
rect 5518 8990 5570 9042
rect 5966 8990 6018 9042
rect 9774 8990 9826 9042
rect 10558 8990 10610 9042
rect 16494 8990 16546 9042
rect 17054 8990 17106 9042
rect 21646 8990 21698 9042
rect 21982 8990 22034 9042
rect 22542 8990 22594 9042
rect 22766 8990 22818 9042
rect 27582 8990 27634 9042
rect 28142 8990 28194 9042
rect 30046 8990 30098 9042
rect 30270 8990 30322 9042
rect 37438 8990 37490 9042
rect 37886 8990 37938 9042
rect 38782 8990 38834 9042
rect 39230 8990 39282 9042
rect 39566 8990 39618 9042
rect 40462 8990 40514 9042
rect 40686 8990 40738 9042
rect 42926 8990 42978 9042
rect 47182 8990 47234 9042
rect 47742 8990 47794 9042
rect 50654 8990 50706 9042
rect 51550 8990 51602 9042
rect 51886 8990 51938 9042
rect 52782 8990 52834 9042
rect 53006 8990 53058 9042
rect 54238 8990 54290 9042
rect 56030 8990 56082 9042
rect 58046 8990 58098 9042
rect 13358 8878 13410 8930
rect 17614 8878 17666 8930
rect 18062 8878 18114 8930
rect 18622 8878 18674 8930
rect 23998 8878 24050 8930
rect 29150 8878 29202 8930
rect 29822 8878 29874 8930
rect 31838 8878 31890 8930
rect 37550 8878 37602 8930
rect 39006 8878 39058 8930
rect 39790 8878 39842 8930
rect 42814 8878 42866 8930
rect 46622 8878 46674 8930
rect 56254 8878 56306 8930
rect 56702 8878 56754 8930
rect 28142 8766 28194 8818
rect 28478 8766 28530 8818
rect 43934 8766 43986 8818
rect 49870 8766 49922 8818
rect 50990 8766 51042 8818
rect 57934 8766 57986 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 29710 8430 29762 8482
rect 39566 8430 39618 8482
rect 55022 8430 55074 8482
rect 56926 8430 56978 8482
rect 6750 8318 6802 8370
rect 8094 8318 8146 8370
rect 13022 8318 13074 8370
rect 19070 8318 19122 8370
rect 22878 8318 22930 8370
rect 25454 8318 25506 8370
rect 32286 8318 32338 8370
rect 33294 8318 33346 8370
rect 34078 8318 34130 8370
rect 35198 8318 35250 8370
rect 38110 8318 38162 8370
rect 41582 8318 41634 8370
rect 43150 8318 43202 8370
rect 47070 8318 47122 8370
rect 56590 8318 56642 8370
rect 7758 8206 7810 8258
rect 9550 8206 9602 8258
rect 9886 8206 9938 8258
rect 15038 8206 15090 8258
rect 15374 8206 15426 8258
rect 18622 8206 18674 8258
rect 22654 8206 22706 8258
rect 23326 8206 23378 8258
rect 24222 8206 24274 8258
rect 24670 8206 24722 8258
rect 26014 8206 26066 8258
rect 26686 8206 26738 8258
rect 27806 8206 27858 8258
rect 28254 8206 28306 8258
rect 29822 8206 29874 8258
rect 31950 8206 32002 8258
rect 32174 8206 32226 8258
rect 32510 8206 32562 8258
rect 34302 8206 34354 8258
rect 35534 8206 35586 8258
rect 35982 8206 36034 8258
rect 37886 8206 37938 8258
rect 39118 8206 39170 8258
rect 39342 8206 39394 8258
rect 39678 8206 39730 8258
rect 40798 8206 40850 8258
rect 42478 8206 42530 8258
rect 42702 8206 42754 8258
rect 42926 8206 42978 8258
rect 44158 8206 44210 8258
rect 44606 8206 44658 8258
rect 46958 8206 47010 8258
rect 49086 8206 49138 8258
rect 49534 8206 49586 8258
rect 51102 8206 51154 8258
rect 52110 8206 52162 8258
rect 52670 8206 52722 8258
rect 53454 8206 53506 8258
rect 54238 8206 54290 8258
rect 54686 8206 54738 8258
rect 55918 8206 55970 8258
rect 56702 8206 56754 8258
rect 8206 8094 8258 8146
rect 21982 8094 22034 8146
rect 23102 8094 23154 8146
rect 23998 8094 24050 8146
rect 26238 8094 26290 8146
rect 27134 8094 27186 8146
rect 28814 8094 28866 8146
rect 30606 8094 30658 8146
rect 35310 8094 35362 8146
rect 38558 8094 38610 8146
rect 44718 8094 44770 8146
rect 47854 8094 47906 8146
rect 49758 8094 49810 8146
rect 50766 8094 50818 8146
rect 53678 8094 53730 8146
rect 55582 8094 55634 8146
rect 7198 7982 7250 8034
rect 7982 7982 8034 8034
rect 8654 7982 8706 8034
rect 12462 7982 12514 8034
rect 13582 7982 13634 8034
rect 14030 7982 14082 8034
rect 17950 7982 18002 8034
rect 19518 7982 19570 8034
rect 20862 7982 20914 8034
rect 21646 7982 21698 8034
rect 26350 7982 26402 8034
rect 27246 7982 27298 8034
rect 29710 7982 29762 8034
rect 30270 7982 30322 8034
rect 30494 7982 30546 8034
rect 31166 7982 31218 8034
rect 32846 7982 32898 8034
rect 34638 7982 34690 8034
rect 39902 7982 39954 8034
rect 40574 7982 40626 8034
rect 40910 7982 40962 8034
rect 41022 7982 41074 8034
rect 42590 7982 42642 8034
rect 45950 7982 46002 8034
rect 57710 7982 57762 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 12798 7646 12850 7698
rect 13358 7646 13410 7698
rect 18734 7646 18786 7698
rect 19182 7646 19234 7698
rect 22094 7646 22146 7698
rect 22878 7646 22930 7698
rect 27470 7646 27522 7698
rect 33630 7646 33682 7698
rect 39566 7646 39618 7698
rect 41582 7646 41634 7698
rect 42030 7646 42082 7698
rect 44494 7646 44546 7698
rect 53230 7646 53282 7698
rect 53454 7646 53506 7698
rect 54462 7646 54514 7698
rect 54686 7646 54738 7698
rect 55918 7646 55970 7698
rect 6190 7534 6242 7586
rect 8990 7534 9042 7586
rect 20862 7534 20914 7586
rect 22206 7534 22258 7586
rect 22990 7534 23042 7586
rect 23438 7534 23490 7586
rect 24670 7534 24722 7586
rect 24894 7534 24946 7586
rect 25678 7534 25730 7586
rect 25790 7534 25842 7586
rect 27358 7534 27410 7586
rect 27582 7534 27634 7586
rect 28254 7534 28306 7586
rect 34750 7534 34802 7586
rect 34974 7534 35026 7586
rect 37326 7534 37378 7586
rect 45390 7534 45442 7586
rect 46958 7534 47010 7586
rect 50654 7534 50706 7586
rect 53118 7534 53170 7586
rect 54350 7534 54402 7586
rect 5854 7422 5906 7474
rect 8318 7422 8370 7474
rect 9662 7422 9714 7474
rect 10222 7422 10274 7474
rect 21086 7422 21138 7474
rect 23214 7422 23266 7474
rect 24222 7422 24274 7474
rect 24446 7422 24498 7474
rect 26014 7422 26066 7474
rect 28814 7422 28866 7474
rect 29822 7422 29874 7474
rect 31614 7422 31666 7474
rect 32622 7422 32674 7474
rect 37662 7422 37714 7474
rect 39902 7422 39954 7474
rect 40126 7422 40178 7474
rect 43150 7422 43202 7474
rect 46062 7422 46114 7474
rect 46510 7422 46562 7474
rect 49982 7422 50034 7474
rect 50878 7422 50930 7474
rect 55358 7422 55410 7474
rect 55582 7422 55634 7474
rect 5182 7310 5234 7362
rect 8094 7310 8146 7362
rect 13694 7310 13746 7362
rect 19630 7310 19682 7362
rect 26798 7310 26850 7362
rect 30270 7310 30322 7362
rect 31278 7310 31330 7362
rect 32174 7310 32226 7362
rect 42478 7310 42530 7362
rect 42926 7310 42978 7362
rect 43934 7310 43986 7362
rect 50990 7310 51042 7362
rect 53790 7310 53842 7362
rect 29934 7198 29986 7250
rect 30158 7198 30210 7250
rect 34638 7198 34690 7250
rect 37662 7198 37714 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 18734 6862 18786 6914
rect 31838 6862 31890 6914
rect 13582 6750 13634 6802
rect 27022 6750 27074 6802
rect 28030 6750 28082 6802
rect 30718 6750 30770 6802
rect 32846 6750 32898 6802
rect 34638 6750 34690 6802
rect 43822 6750 43874 6802
rect 6750 6638 6802 6690
rect 7646 6638 7698 6690
rect 8542 6638 8594 6690
rect 8878 6638 8930 6690
rect 9550 6638 9602 6690
rect 9998 6638 10050 6690
rect 15038 6638 15090 6690
rect 15710 6638 15762 6690
rect 19630 6638 19682 6690
rect 20638 6638 20690 6690
rect 22542 6638 22594 6690
rect 24670 6638 24722 6690
rect 25790 6638 25842 6690
rect 26462 6638 26514 6690
rect 26686 6638 26738 6690
rect 28590 6638 28642 6690
rect 31614 6638 31666 6690
rect 32174 6638 32226 6690
rect 34862 6638 34914 6690
rect 35982 6638 36034 6690
rect 4734 6526 4786 6578
rect 4846 6526 4898 6578
rect 20302 6526 20354 6578
rect 21982 6526 22034 6578
rect 23998 6526 24050 6578
rect 24222 6526 24274 6578
rect 27582 6526 27634 6578
rect 28702 6526 28754 6578
rect 35534 6526 35586 6578
rect 5070 6414 5122 6466
rect 5630 6414 5682 6466
rect 6526 6414 6578 6466
rect 7982 6414 8034 6466
rect 12462 6414 12514 6466
rect 13022 6414 13074 6466
rect 14030 6414 14082 6466
rect 14478 6414 14530 6466
rect 17950 6414 18002 6466
rect 19406 6414 19458 6466
rect 21646 6414 21698 6466
rect 22990 6414 23042 6466
rect 23438 6414 23490 6466
rect 24446 6414 24498 6466
rect 25454 6414 25506 6466
rect 29822 6414 29874 6466
rect 30270 6414 30322 6466
rect 32734 6414 32786 6466
rect 32958 6414 33010 6466
rect 33182 6414 33234 6466
rect 33742 6414 33794 6466
rect 45390 6414 45442 6466
rect 55022 6414 55074 6466
rect 55470 6414 55522 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 8318 6078 8370 6130
rect 9102 6078 9154 6130
rect 13246 6078 13298 6130
rect 14366 6078 14418 6130
rect 15150 6078 15202 6130
rect 20526 6078 20578 6130
rect 23326 6078 23378 6130
rect 23550 6078 23602 6130
rect 24446 6078 24498 6130
rect 26014 6078 26066 6130
rect 27022 6078 27074 6130
rect 28590 6078 28642 6130
rect 30606 6078 30658 6130
rect 30830 6078 30882 6130
rect 44494 6078 44546 6130
rect 45278 6078 45330 6130
rect 47966 6078 48018 6130
rect 21982 5966 22034 6018
rect 23102 5966 23154 6018
rect 26462 5966 26514 6018
rect 29038 5966 29090 6018
rect 29374 5966 29426 6018
rect 33630 5966 33682 6018
rect 35534 5966 35586 6018
rect 41582 5966 41634 6018
rect 45502 5966 45554 6018
rect 46286 5966 46338 6018
rect 47070 5966 47122 6018
rect 5630 5854 5682 5906
rect 6078 5854 6130 5906
rect 10110 5854 10162 5906
rect 10782 5854 10834 5906
rect 15710 5854 15762 5906
rect 16158 5854 16210 5906
rect 16718 5854 16770 5906
rect 17614 5854 17666 5906
rect 18286 5854 18338 5906
rect 22206 5854 22258 5906
rect 23662 5854 23714 5906
rect 23998 5854 24050 5906
rect 24558 5854 24610 5906
rect 24670 5854 24722 5906
rect 27918 5854 27970 5906
rect 30942 5854 30994 5906
rect 32062 5854 32114 5906
rect 32398 5854 32450 5906
rect 32510 5854 32562 5906
rect 33854 5854 33906 5906
rect 34862 5854 34914 5906
rect 35086 5854 35138 5906
rect 35310 5854 35362 5906
rect 35758 5854 35810 5906
rect 36542 5854 36594 5906
rect 36990 5854 37042 5906
rect 39454 5854 39506 5906
rect 39678 5854 39730 5906
rect 43822 5854 43874 5906
rect 44382 5854 44434 5906
rect 44606 5854 44658 5906
rect 45166 5854 45218 5906
rect 46174 5854 46226 5906
rect 46958 5854 47010 5906
rect 47854 5854 47906 5906
rect 9662 5742 9714 5794
rect 27694 5742 27746 5794
rect 30270 5742 30322 5794
rect 35646 5742 35698 5794
rect 37438 5742 37490 5794
rect 39230 5742 39282 5794
rect 43262 5742 43314 5794
rect 13806 5630 13858 5682
rect 21310 5630 21362 5682
rect 27582 5630 27634 5682
rect 40126 5630 40178 5682
rect 41806 5630 41858 5682
rect 42142 5630 42194 5682
rect 44158 5630 44210 5682
rect 46286 5630 46338 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 5854 5294 5906 5346
rect 26910 5294 26962 5346
rect 41470 5294 41522 5346
rect 45502 5294 45554 5346
rect 49646 5294 49698 5346
rect 5966 5182 6018 5234
rect 9662 5182 9714 5234
rect 13582 5182 13634 5234
rect 14254 5182 14306 5234
rect 14926 5182 14978 5234
rect 19854 5182 19906 5234
rect 24782 5182 24834 5234
rect 25230 5182 25282 5234
rect 26350 5182 26402 5234
rect 28366 5182 28418 5234
rect 34190 5182 34242 5234
rect 34750 5182 34802 5234
rect 42926 5182 42978 5234
rect 45838 5182 45890 5234
rect 47294 5182 47346 5234
rect 48750 5182 48802 5234
rect 49198 5182 49250 5234
rect 6638 5070 6690 5122
rect 8318 5070 8370 5122
rect 15374 5070 15426 5122
rect 16046 5070 16098 5122
rect 19070 5070 19122 5122
rect 20302 5070 20354 5122
rect 20862 5070 20914 5122
rect 23102 5070 23154 5122
rect 25454 5070 25506 5122
rect 27470 5070 27522 5122
rect 28142 5070 28194 5122
rect 28478 5070 28530 5122
rect 29710 5070 29762 5122
rect 31950 5070 32002 5122
rect 34974 5070 35026 5122
rect 35646 5070 35698 5122
rect 36430 5070 36482 5122
rect 37662 5070 37714 5122
rect 38110 5070 38162 5122
rect 38558 5070 38610 5122
rect 39230 5070 39282 5122
rect 39678 5070 39730 5122
rect 39902 5070 39954 5122
rect 41022 5070 41074 5122
rect 41358 5070 41410 5122
rect 41694 5070 41746 5122
rect 41806 5070 41858 5122
rect 43038 5070 43090 5122
rect 44046 5070 44098 5122
rect 44606 5070 44658 5122
rect 47742 5070 47794 5122
rect 48974 5070 49026 5122
rect 21870 4958 21922 5010
rect 23214 4958 23266 5010
rect 27358 4958 27410 5010
rect 27582 4958 27634 5010
rect 28814 4958 28866 5010
rect 30382 4958 30434 5010
rect 33518 4958 33570 5010
rect 36654 4958 36706 5010
rect 41918 4958 41970 5010
rect 42478 4958 42530 5010
rect 42702 4958 42754 5010
rect 44718 4958 44770 5010
rect 48190 4958 48242 5010
rect 18286 4846 18338 4898
rect 21982 4846 22034 4898
rect 31838 4846 31890 4898
rect 36542 4846 36594 4898
rect 39790 4846 39842 4898
rect 45726 4846 45778 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 8430 4510 8482 4562
rect 20750 4510 20802 4562
rect 23214 4510 23266 4562
rect 23438 4510 23490 4562
rect 24110 4510 24162 4562
rect 24558 4510 24610 4562
rect 25006 4510 25058 4562
rect 25790 4510 25842 4562
rect 30382 4510 30434 4562
rect 32846 4510 32898 4562
rect 40686 4510 40738 4562
rect 40910 4510 40962 4562
rect 43150 4510 43202 4562
rect 45726 4510 45778 4562
rect 45950 4510 46002 4562
rect 15038 4398 15090 4450
rect 21758 4398 21810 4450
rect 23550 4398 23602 4450
rect 26014 4398 26066 4450
rect 26238 4398 26290 4450
rect 28030 4398 28082 4450
rect 28590 4398 28642 4450
rect 28926 4398 28978 4450
rect 32398 4398 32450 4450
rect 33630 4398 33682 4450
rect 35198 4398 35250 4450
rect 40574 4398 40626 4450
rect 44046 4398 44098 4450
rect 45614 4398 45666 4450
rect 48638 4398 48690 4450
rect 5630 4286 5682 4338
rect 6078 4286 6130 4338
rect 9102 4286 9154 4338
rect 9774 4286 9826 4338
rect 13022 4286 13074 4338
rect 17614 4286 17666 4338
rect 18174 4286 18226 4338
rect 21310 4286 21362 4338
rect 22206 4286 22258 4338
rect 25566 4286 25618 4338
rect 27246 4286 27298 4338
rect 28366 4286 28418 4338
rect 28478 4286 28530 4338
rect 29262 4286 29314 4338
rect 31502 4286 31554 4338
rect 33854 4286 33906 4338
rect 35534 4286 35586 4338
rect 36094 4286 36146 4338
rect 37214 4286 37266 4338
rect 37438 4286 37490 4338
rect 42030 4286 42082 4338
rect 44494 4286 44546 4338
rect 48078 4286 48130 4338
rect 48302 4286 48354 4338
rect 48526 4286 48578 4338
rect 10222 4174 10274 4226
rect 22654 4174 22706 4226
rect 26910 4174 26962 4226
rect 27470 4174 27522 4226
rect 28142 4174 28194 4226
rect 29598 4174 29650 4226
rect 31838 4174 31890 4226
rect 34414 4174 34466 4226
rect 35422 4174 35474 4226
rect 36206 4174 36258 4226
rect 36990 4174 37042 4226
rect 38782 4174 38834 4226
rect 41918 4174 41970 4226
rect 42590 4174 42642 4226
rect 44830 4174 44882 4226
rect 37886 4062 37938 4114
rect 39006 4062 39058 4114
rect 39342 4062 39394 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 25454 3726 25506 3778
rect 25902 3726 25954 3778
rect 27694 3726 27746 3778
rect 28478 3726 28530 3778
rect 6750 3614 6802 3666
rect 7310 3614 7362 3666
rect 7646 3614 7698 3666
rect 9662 3614 9714 3666
rect 10110 3614 10162 3666
rect 15038 3614 15090 3666
rect 16382 3614 16434 3666
rect 16830 3614 16882 3666
rect 18174 3614 18226 3666
rect 19630 3614 19682 3666
rect 22094 3614 22146 3666
rect 22878 3614 22930 3666
rect 23326 3614 23378 3666
rect 23774 3614 23826 3666
rect 24222 3614 24274 3666
rect 24670 3614 24722 3666
rect 25454 3614 25506 3666
rect 25902 3614 25954 3666
rect 26350 3614 26402 3666
rect 26798 3614 26850 3666
rect 27694 3614 27746 3666
rect 28590 3614 28642 3666
rect 29710 3614 29762 3666
rect 32286 3614 32338 3666
rect 33070 3614 33122 3666
rect 34078 3614 34130 3666
rect 34526 3614 34578 3666
rect 35422 3614 35474 3666
rect 35758 3614 35810 3666
rect 36206 3614 36258 3666
rect 39454 3614 39506 3666
rect 47518 3614 47570 3666
rect 5070 3502 5122 3554
rect 5854 3502 5906 3554
rect 6302 3502 6354 3554
rect 17726 3502 17778 3554
rect 18622 3502 18674 3554
rect 21310 3502 21362 3554
rect 21646 3502 21698 3554
rect 28142 3502 28194 3554
rect 29262 3502 29314 3554
rect 31614 3502 31666 3554
rect 32174 3502 32226 3554
rect 37102 3502 37154 3554
rect 37326 3502 37378 3554
rect 41022 3502 41074 3554
rect 42142 3502 42194 3554
rect 12910 3390 12962 3442
rect 13694 3390 13746 3442
rect 21534 3390 21586 3442
rect 27246 3390 27298 3442
rect 30382 3390 30434 3442
rect 34974 3390 35026 3442
rect 37550 3390 37602 3442
rect 38558 3390 38610 3442
rect 40350 3390 40402 3442
rect 41134 3390 41186 3442
rect 41358 3390 41410 3442
rect 41806 3390 41858 3442
rect 41918 3390 41970 3442
rect 48750 3390 48802 3442
rect 55694 3390 55746 3442
rect 56590 3390 56642 3442
rect 30718 3278 30770 3330
rect 37214 3278 37266 3330
rect 39006 3278 39058 3330
rect 48078 3278 48130 3330
rect 55358 3278 55410 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
rect 47406 2942 47458 2994
rect 48078 2942 48130 2994
<< metal2 >>
rect 10080 63181 10192 63981
rect 30128 63181 30240 63981
rect 50176 63181 50288 63981
rect 10108 62188 10164 63181
rect 10108 62132 10500 62188
rect 1372 60788 1428 60798
rect 1148 56980 1204 56990
rect 1036 52388 1092 52398
rect 924 49924 980 49934
rect 924 40068 980 49868
rect 1036 43316 1092 52332
rect 1036 43250 1092 43260
rect 924 40002 980 40012
rect 1036 33908 1092 33918
rect 1036 23380 1092 33852
rect 1036 23314 1092 23324
rect 1148 19796 1204 56924
rect 1260 52276 1316 52286
rect 1260 48580 1316 52220
rect 1260 48514 1316 48524
rect 1372 42868 1428 60732
rect 1708 60676 1764 60686
rect 1484 55972 1540 55982
rect 1484 48244 1540 55916
rect 1708 55636 1764 60620
rect 4476 60396 4740 60406
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4476 60330 4740 60340
rect 10444 60114 10500 62132
rect 25340 60900 25396 60910
rect 10444 60062 10446 60114
rect 10498 60062 10500 60114
rect 10444 60050 10500 60062
rect 21980 60226 22036 60238
rect 21980 60174 21982 60226
rect 22034 60174 22036 60226
rect 4620 60004 4676 60014
rect 4620 59910 4676 59948
rect 4956 60004 5012 60014
rect 3724 59780 3780 59790
rect 4172 59780 4228 59790
rect 3724 59686 3780 59724
rect 4060 59778 4228 59780
rect 4060 59726 4174 59778
rect 4226 59726 4228 59778
rect 4060 59724 4228 59726
rect 2716 59106 2772 59118
rect 2716 59054 2718 59106
rect 2770 59054 2772 59106
rect 2716 58996 2772 59054
rect 2716 58930 2772 58940
rect 3276 59106 3332 59118
rect 3276 59054 3278 59106
rect 3330 59054 3332 59106
rect 2492 58324 2548 58334
rect 1932 58212 1988 58222
rect 1596 55580 1764 55636
rect 1820 58210 1988 58212
rect 1820 58158 1934 58210
rect 1986 58158 1988 58210
rect 1820 58156 1988 58158
rect 1596 52276 1652 55580
rect 1596 52210 1652 52220
rect 1708 55412 1764 55422
rect 1820 55412 1876 58156
rect 1932 58146 1988 58156
rect 2492 58210 2548 58268
rect 2492 58158 2494 58210
rect 2546 58158 2548 58210
rect 2156 57538 2212 57550
rect 2492 57540 2548 58158
rect 2940 58210 2996 58222
rect 2940 58158 2942 58210
rect 2994 58158 2996 58210
rect 2940 57764 2996 58158
rect 3164 57876 3220 57886
rect 3276 57876 3332 59054
rect 3612 59106 3668 59118
rect 3612 59054 3614 59106
rect 3666 59054 3668 59106
rect 3612 58996 3668 59054
rect 3612 58930 3668 58940
rect 4060 58996 4116 59724
rect 4172 59714 4228 59724
rect 4620 59444 4676 59454
rect 4620 59350 4676 59388
rect 4060 58930 4116 58940
rect 4172 59106 4228 59118
rect 4172 59054 4174 59106
rect 4226 59054 4228 59106
rect 3388 58212 3444 58222
rect 3388 58118 3444 58156
rect 3948 58210 4004 58222
rect 3948 58158 3950 58210
rect 4002 58158 4004 58210
rect 2940 57698 2996 57708
rect 3052 57874 3332 57876
rect 3052 57822 3166 57874
rect 3218 57822 3332 57874
rect 3052 57820 3332 57822
rect 2828 57540 2884 57550
rect 2156 57486 2158 57538
rect 2210 57486 2212 57538
rect 1932 56980 1988 56990
rect 2156 56980 2212 57486
rect 1932 56978 2212 56980
rect 1932 56926 1934 56978
rect 1986 56926 2212 56978
rect 1932 56924 2212 56926
rect 1932 56914 1988 56924
rect 2156 56308 2212 56924
rect 2156 56242 2212 56252
rect 2268 57484 2548 57540
rect 2604 57538 2884 57540
rect 2604 57486 2830 57538
rect 2882 57486 2884 57538
rect 2604 57484 2884 57486
rect 1932 56084 1988 56094
rect 2268 56084 2324 57484
rect 2380 57316 2436 57326
rect 2380 56978 2436 57260
rect 2380 56926 2382 56978
rect 2434 56926 2436 56978
rect 2380 56914 2436 56926
rect 1932 56082 2324 56084
rect 1932 56030 1934 56082
rect 1986 56030 2324 56082
rect 1932 56028 2324 56030
rect 1932 56018 1988 56028
rect 2380 55970 2436 55982
rect 2380 55918 2382 55970
rect 2434 55918 2436 55970
rect 2380 55860 2436 55918
rect 2380 55794 2436 55804
rect 2380 55636 2436 55646
rect 2268 55524 2324 55534
rect 1820 55356 1988 55412
rect 1708 55188 1764 55356
rect 1820 55188 1876 55198
rect 1708 55186 1876 55188
rect 1708 55134 1822 55186
rect 1874 55134 1876 55186
rect 1708 55132 1876 55134
rect 1708 51154 1764 55132
rect 1820 55122 1876 55132
rect 1820 54628 1876 54638
rect 1820 54534 1876 54572
rect 1932 53956 1988 55356
rect 1932 53890 1988 53900
rect 2156 55074 2212 55086
rect 2156 55022 2158 55074
rect 2210 55022 2212 55074
rect 2156 54290 2212 55022
rect 2268 54738 2324 55468
rect 2268 54686 2270 54738
rect 2322 54686 2324 54738
rect 2268 54674 2324 54686
rect 2156 54238 2158 54290
rect 2210 54238 2212 54290
rect 2044 53620 2100 53630
rect 2044 53526 2100 53564
rect 2156 53396 2212 54238
rect 2044 53340 2212 53396
rect 2380 53730 2436 55580
rect 2604 55300 2660 57484
rect 2828 57474 2884 57484
rect 2828 56642 2884 56654
rect 2828 56590 2830 56642
rect 2882 56590 2884 56642
rect 2716 56308 2772 56318
rect 2716 56214 2772 56252
rect 2828 56308 2884 56590
rect 2940 56308 2996 56318
rect 2828 56252 2940 56308
rect 2828 55412 2884 56252
rect 2940 56242 2996 56252
rect 3052 55636 3108 57820
rect 3164 57810 3220 57820
rect 3164 57652 3220 57662
rect 3948 57652 4004 58158
rect 4060 57876 4116 57886
rect 4060 57782 4116 57820
rect 4172 57652 4228 59054
rect 4844 59108 4900 59118
rect 4476 58828 4740 58838
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4476 58762 4740 58772
rect 3948 57596 4228 57652
rect 3164 55972 3220 57596
rect 3724 57540 3780 57550
rect 3780 57484 3892 57540
rect 3724 57446 3780 57484
rect 3500 56644 3556 56654
rect 3500 56550 3556 56588
rect 3164 55878 3220 55916
rect 3612 55972 3668 55982
rect 3612 55970 3780 55972
rect 3612 55918 3614 55970
rect 3666 55918 3780 55970
rect 3612 55916 3780 55918
rect 3612 55906 3668 55916
rect 3052 55570 3108 55580
rect 3388 55860 3444 55870
rect 2604 55234 2660 55244
rect 2716 55356 2884 55412
rect 2604 55076 2660 55086
rect 2716 55076 2772 55356
rect 2492 55074 2772 55076
rect 2492 55022 2606 55074
rect 2658 55022 2772 55074
rect 2492 55020 2772 55022
rect 2828 55188 2884 55198
rect 2492 54290 2548 55020
rect 2604 55010 2660 55020
rect 2492 54238 2494 54290
rect 2546 54238 2548 54290
rect 2492 54226 2548 54238
rect 2604 54852 2660 54862
rect 2380 53678 2382 53730
rect 2434 53678 2436 53730
rect 1820 52834 1876 52846
rect 1820 52782 1822 52834
rect 1874 52782 1876 52834
rect 1820 52500 1876 52782
rect 1820 52444 1988 52500
rect 1820 52276 1876 52286
rect 1820 52182 1876 52220
rect 1932 51940 1988 52444
rect 1932 51874 1988 51884
rect 1932 51268 1988 51278
rect 2044 51268 2100 53340
rect 2380 53060 2436 53678
rect 2380 52994 2436 53004
rect 2268 52946 2324 52958
rect 2268 52894 2270 52946
rect 2322 52894 2324 52946
rect 2268 52836 2324 52894
rect 2268 52780 2548 52836
rect 2156 52724 2212 52734
rect 2156 52276 2212 52668
rect 2492 52386 2548 52780
rect 2492 52334 2494 52386
rect 2546 52334 2548 52386
rect 2268 52276 2324 52286
rect 2156 52274 2436 52276
rect 2156 52222 2270 52274
rect 2322 52222 2436 52274
rect 2156 52220 2436 52222
rect 2268 52210 2324 52220
rect 2268 51940 2324 51950
rect 2268 51602 2324 51884
rect 2268 51550 2270 51602
rect 2322 51550 2324 51602
rect 2268 51538 2324 51550
rect 1988 51212 2100 51268
rect 1932 51174 1988 51212
rect 1708 51102 1710 51154
rect 1762 51102 1764 51154
rect 1708 51090 1764 51102
rect 2156 50596 2212 50634
rect 2156 50530 2212 50540
rect 1820 50484 1876 50494
rect 2380 50428 2436 52220
rect 1484 48178 1540 48188
rect 1596 49252 1652 49262
rect 1596 47908 1652 49196
rect 1372 42802 1428 42812
rect 1484 47852 1652 47908
rect 1372 38836 1428 38846
rect 1372 36372 1428 38780
rect 1484 38164 1540 47852
rect 1596 47684 1652 47694
rect 1596 40292 1652 47628
rect 1820 47236 1876 50428
rect 2156 50372 2436 50428
rect 2044 49698 2100 49710
rect 2044 49646 2046 49698
rect 2098 49646 2100 49698
rect 2044 49586 2100 49646
rect 2044 49534 2046 49586
rect 2098 49534 2100 49586
rect 1932 49250 1988 49262
rect 1932 49198 1934 49250
rect 1986 49198 1988 49250
rect 1932 49138 1988 49198
rect 1932 49086 1934 49138
rect 1986 49086 1988 49138
rect 1932 49074 1988 49086
rect 2044 48916 2100 49534
rect 1708 47234 1876 47236
rect 1708 47182 1822 47234
rect 1874 47182 1876 47234
rect 1708 47180 1876 47182
rect 1708 41858 1764 47180
rect 1820 47170 1876 47180
rect 1932 48860 2100 48916
rect 1932 46900 1988 48860
rect 2044 48692 2100 48702
rect 2044 48466 2100 48636
rect 2044 48414 2046 48466
rect 2098 48414 2100 48466
rect 2044 48402 2100 48414
rect 1820 46844 1988 46900
rect 1820 46452 1876 46844
rect 2156 46788 2212 50372
rect 2380 49812 2436 49822
rect 2380 49718 2436 49756
rect 2380 48802 2436 48814
rect 2380 48750 2382 48802
rect 2434 48750 2436 48802
rect 2268 48468 2324 48478
rect 2268 48132 2324 48412
rect 2380 48356 2436 48750
rect 2380 48290 2436 48300
rect 2380 48132 2436 48142
rect 2268 48130 2436 48132
rect 2268 48078 2382 48130
rect 2434 48078 2436 48130
rect 2268 48076 2436 48078
rect 2380 48066 2436 48076
rect 2268 47348 2324 47358
rect 2268 47234 2324 47292
rect 2268 47182 2270 47234
rect 2322 47182 2324 47234
rect 2268 47170 2324 47182
rect 2380 47012 2436 47022
rect 2380 46898 2436 46956
rect 2380 46846 2382 46898
rect 2434 46846 2436 46898
rect 2380 46834 2436 46846
rect 2156 46722 2212 46732
rect 1932 46564 1988 46574
rect 1932 46562 2100 46564
rect 1932 46510 1934 46562
rect 1986 46510 2100 46562
rect 1932 46508 2100 46510
rect 1932 46498 1988 46508
rect 1820 46386 1876 46396
rect 1932 46116 1988 46126
rect 1932 46002 1988 46060
rect 1932 45950 1934 46002
rect 1986 45950 1988 46002
rect 1932 45938 1988 45950
rect 2044 46004 2100 46508
rect 2492 46004 2548 52334
rect 2604 52164 2660 54796
rect 2716 54740 2772 54750
rect 2716 54646 2772 54684
rect 2828 53732 2884 55132
rect 3052 55076 3108 55086
rect 2716 53676 2884 53732
rect 2940 55074 3108 55076
rect 2940 55022 3054 55074
rect 3106 55022 3108 55074
rect 2940 55020 3108 55022
rect 2716 53172 2772 53676
rect 2716 53106 2772 53116
rect 2828 53506 2884 53518
rect 2828 53454 2830 53506
rect 2882 53454 2884 53506
rect 2828 52948 2884 53454
rect 2940 53396 2996 55020
rect 3052 55010 3108 55020
rect 3164 54402 3220 54414
rect 3164 54350 3166 54402
rect 3218 54350 3220 54402
rect 3164 53732 3220 54350
rect 3388 54404 3444 55804
rect 3612 55636 3668 55646
rect 3612 55410 3668 55580
rect 3612 55358 3614 55410
rect 3666 55358 3668 55410
rect 3612 55346 3668 55358
rect 3724 55076 3780 55916
rect 3724 55010 3780 55020
rect 3500 54404 3556 54414
rect 3388 54402 3556 54404
rect 3388 54350 3502 54402
rect 3554 54350 3556 54402
rect 3388 54348 3556 54350
rect 3276 53844 3332 53854
rect 3276 53750 3332 53788
rect 3164 53666 3220 53676
rect 2940 53330 2996 53340
rect 3052 53508 3108 53518
rect 2828 52882 2884 52892
rect 2940 53172 2996 53182
rect 2716 52834 2772 52846
rect 2716 52782 2718 52834
rect 2770 52782 2772 52834
rect 2716 52386 2772 52782
rect 2716 52334 2718 52386
rect 2770 52334 2772 52386
rect 2716 52322 2772 52334
rect 2604 52108 2772 52164
rect 2604 51940 2660 51950
rect 2604 51846 2660 51884
rect 2716 51716 2772 52108
rect 2604 51660 2772 51716
rect 2604 50932 2660 51660
rect 2716 51266 2772 51278
rect 2716 51214 2718 51266
rect 2770 51214 2772 51266
rect 2716 51156 2772 51214
rect 2716 51154 2884 51156
rect 2716 51102 2718 51154
rect 2770 51102 2884 51154
rect 2716 51100 2884 51102
rect 2716 51090 2772 51100
rect 2604 50876 2772 50932
rect 2604 50708 2660 50718
rect 2604 50614 2660 50652
rect 2716 50428 2772 50876
rect 2604 50372 2772 50428
rect 2604 49250 2660 50372
rect 2604 49198 2606 49250
rect 2658 49198 2660 49250
rect 2604 49186 2660 49198
rect 2828 49028 2884 51100
rect 2940 50706 2996 53116
rect 3052 53170 3108 53452
rect 3052 53118 3054 53170
rect 3106 53118 3108 53170
rect 3052 53106 3108 53118
rect 3164 53396 3220 53406
rect 3052 52836 3108 52846
rect 3052 52274 3108 52780
rect 3052 52222 3054 52274
rect 3106 52222 3108 52274
rect 3052 52164 3108 52222
rect 3164 52276 3220 53340
rect 3164 52210 3220 52220
rect 3276 52948 3332 52958
rect 3052 52098 3108 52108
rect 2940 50654 2942 50706
rect 2994 50654 2996 50706
rect 2940 50148 2996 50654
rect 2940 50082 2996 50092
rect 3164 51604 3220 51614
rect 3276 51604 3332 52892
rect 3164 51602 3332 51604
rect 3164 51550 3166 51602
rect 3218 51550 3332 51602
rect 3164 51548 3332 51550
rect 2940 49700 2996 49710
rect 2940 49606 2996 49644
rect 3164 49586 3220 51548
rect 3388 51492 3444 54348
rect 3500 54338 3556 54348
rect 3836 53956 3892 57484
rect 3948 56642 4004 56654
rect 3948 56590 3950 56642
rect 4002 56590 4004 56642
rect 3948 55076 4004 56590
rect 4060 56084 4116 56094
rect 4060 55970 4116 56028
rect 4060 55918 4062 55970
rect 4114 55918 4116 55970
rect 4060 55636 4116 55918
rect 4060 55570 4116 55580
rect 3948 55010 4004 55020
rect 4172 54964 4228 57596
rect 4508 58210 4564 58222
rect 4508 58158 4510 58210
rect 4562 58158 4564 58210
rect 4508 57988 4564 58158
rect 4508 57428 4564 57932
rect 4620 57540 4676 57550
rect 4620 57446 4676 57484
rect 4508 57362 4564 57372
rect 4476 57260 4740 57270
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4476 57194 4740 57204
rect 4844 56868 4900 59052
rect 4956 58210 5012 59948
rect 9772 60004 9828 60014
rect 11340 60004 11396 60014
rect 9772 59910 9828 59948
rect 11004 60002 11396 60004
rect 11004 59950 11342 60002
rect 11394 59950 11396 60002
rect 11004 59948 11396 59950
rect 5068 59892 5124 59902
rect 5068 59798 5124 59836
rect 5852 59892 5908 59902
rect 5852 59778 5908 59836
rect 6300 59892 6356 59902
rect 6300 59798 6356 59836
rect 7644 59892 7700 59902
rect 5852 59726 5854 59778
rect 5906 59726 5908 59778
rect 5740 59444 5796 59454
rect 5068 59332 5124 59342
rect 5068 59238 5124 59276
rect 5404 59108 5460 59118
rect 5404 59106 5684 59108
rect 5404 59054 5406 59106
rect 5458 59054 5684 59106
rect 5404 59052 5684 59054
rect 5404 59042 5460 59052
rect 4956 58158 4958 58210
rect 5010 58158 5012 58210
rect 4956 57876 5012 58158
rect 4956 57810 5012 57820
rect 5068 57540 5124 57550
rect 5068 57446 5124 57484
rect 5516 57538 5572 57550
rect 5516 57486 5518 57538
rect 5570 57486 5572 57538
rect 4732 56812 4900 56868
rect 4284 56644 4340 56654
rect 4284 56550 4340 56588
rect 4620 55972 4676 55982
rect 4620 55878 4676 55916
rect 4732 55860 4788 56812
rect 4732 55794 4788 55804
rect 4844 56642 4900 56654
rect 4844 56590 4846 56642
rect 4898 56590 4900 56642
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 4844 55300 4900 56590
rect 5180 56644 5236 56654
rect 5068 55970 5124 55982
rect 5068 55918 5070 55970
rect 5122 55918 5124 55970
rect 5068 55860 5124 55918
rect 5068 55524 5124 55804
rect 5068 55458 5124 55468
rect 4844 55234 4900 55244
rect 4172 54898 4228 54908
rect 4396 55074 4452 55086
rect 4396 55022 4398 55074
rect 4450 55022 4452 55074
rect 4396 54964 4452 55022
rect 4844 55076 4900 55086
rect 4844 54982 4900 55020
rect 4396 54898 4452 54908
rect 4396 54516 4452 54526
rect 4396 54422 4452 54460
rect 4956 54516 5012 54526
rect 4956 54422 5012 54460
rect 3948 54404 4004 54414
rect 3948 54310 4004 54348
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 3724 53900 3892 53956
rect 4508 53956 4564 53966
rect 3724 53842 3780 53900
rect 3724 53790 3726 53842
rect 3778 53790 3780 53842
rect 3724 53284 3780 53790
rect 4284 53844 4340 53854
rect 3724 53218 3780 53228
rect 3836 53732 3892 53742
rect 3500 52836 3556 52846
rect 3500 52742 3556 52780
rect 3276 51436 3444 51492
rect 3276 49812 3332 51436
rect 3612 51380 3668 51390
rect 3612 51286 3668 51324
rect 3836 51156 3892 53676
rect 4172 53732 4228 53742
rect 4172 53638 4228 53676
rect 4172 52834 4228 52846
rect 4172 52782 4174 52834
rect 4226 52782 4228 52834
rect 3836 51090 3892 51100
rect 3948 51938 4004 51950
rect 3948 51886 3950 51938
rect 4002 51886 4004 51938
rect 3836 50708 3892 50718
rect 3388 50596 3444 50606
rect 3388 50260 3444 50540
rect 3724 50596 3780 50606
rect 3388 50034 3444 50204
rect 3388 49982 3390 50034
rect 3442 49982 3444 50034
rect 3388 49970 3444 49982
rect 3500 50372 3556 50382
rect 3500 50036 3556 50316
rect 3500 49970 3556 49980
rect 3612 50148 3668 50158
rect 3276 49746 3332 49756
rect 3164 49534 3166 49586
rect 3218 49534 3220 49586
rect 3164 49522 3220 49534
rect 2716 48972 2884 49028
rect 3052 49250 3108 49262
rect 3052 49198 3054 49250
rect 3106 49198 3108 49250
rect 2604 47460 2660 47470
rect 2604 47366 2660 47404
rect 2044 45938 2100 45948
rect 2268 45948 2548 46004
rect 2604 46452 2660 46462
rect 2156 45220 2212 45230
rect 1932 45164 2156 45220
rect 1708 41806 1710 41858
rect 1762 41806 1764 41858
rect 1708 41794 1764 41806
rect 1820 45108 1876 45118
rect 1596 40226 1652 40236
rect 1708 41636 1764 41646
rect 1484 38098 1540 38108
rect 1596 40068 1652 40078
rect 1596 37492 1652 40012
rect 1596 37426 1652 37436
rect 1708 36484 1764 41580
rect 1820 40514 1876 45052
rect 1932 43988 1988 45164
rect 2156 45126 2212 45164
rect 1932 43762 1988 43932
rect 1932 43710 1934 43762
rect 1986 43710 1988 43762
rect 1932 43698 1988 43710
rect 2156 44212 2212 44222
rect 2156 42866 2212 44156
rect 2156 42814 2158 42866
rect 2210 42814 2212 42866
rect 2156 42802 2212 42814
rect 1820 40462 1822 40514
rect 1874 40462 1876 40514
rect 1820 40450 1876 40462
rect 1932 41860 1988 41870
rect 1820 38948 1876 38958
rect 1820 37492 1876 38892
rect 1932 38724 1988 41804
rect 2044 41860 2100 41870
rect 2044 41858 2212 41860
rect 2044 41806 2046 41858
rect 2098 41806 2212 41858
rect 2044 41804 2212 41806
rect 2044 41794 2100 41804
rect 2044 40962 2100 40974
rect 2044 40910 2046 40962
rect 2098 40910 2100 40962
rect 2044 40180 2100 40910
rect 2044 40114 2100 40124
rect 2156 39508 2212 41804
rect 2156 39442 2212 39452
rect 2268 41410 2324 45948
rect 2492 45778 2548 45790
rect 2492 45726 2494 45778
rect 2546 45726 2548 45778
rect 2492 45444 2548 45726
rect 2492 45108 2548 45388
rect 2492 45042 2548 45052
rect 2380 44996 2436 45006
rect 2380 44902 2436 44940
rect 2604 44100 2660 46396
rect 2716 45892 2772 48972
rect 2828 48802 2884 48814
rect 2828 48750 2830 48802
rect 2882 48750 2884 48802
rect 2828 48466 2884 48750
rect 2828 48414 2830 48466
rect 2882 48414 2884 48466
rect 2828 48020 2884 48414
rect 2828 47954 2884 47964
rect 2828 47684 2884 47694
rect 2828 47570 2884 47628
rect 2828 47518 2830 47570
rect 2882 47518 2884 47570
rect 2828 47506 2884 47518
rect 2940 46788 2996 46798
rect 2828 46676 2884 46686
rect 2828 46582 2884 46620
rect 2828 45892 2884 45902
rect 2716 45890 2884 45892
rect 2716 45838 2830 45890
rect 2882 45838 2884 45890
rect 2716 45836 2884 45838
rect 2828 45220 2884 45836
rect 2828 45154 2884 45164
rect 2940 45108 2996 46732
rect 2940 45042 2996 45052
rect 3052 45330 3108 49198
rect 3276 49028 3332 49038
rect 3276 48804 3332 48972
rect 3276 48802 3444 48804
rect 3276 48750 3278 48802
rect 3330 48750 3444 48802
rect 3276 48748 3444 48750
rect 3276 48738 3332 48748
rect 3388 48466 3444 48748
rect 3388 48414 3390 48466
rect 3442 48414 3444 48466
rect 3388 48402 3444 48414
rect 3500 48132 3556 48142
rect 3500 47570 3556 48076
rect 3612 47796 3668 50092
rect 3724 48020 3780 50540
rect 3836 49138 3892 50652
rect 3948 50484 4004 51886
rect 4172 51604 4228 52782
rect 4284 52388 4340 53788
rect 4508 53170 4564 53900
rect 4956 53732 5012 53742
rect 4956 53638 5012 53676
rect 4508 53118 4510 53170
rect 4562 53118 4564 53170
rect 4508 53106 4564 53118
rect 5068 53396 5124 53406
rect 5068 53170 5124 53340
rect 5068 53118 5070 53170
rect 5122 53118 5124 53170
rect 5068 53106 5124 53118
rect 5180 52836 5236 56588
rect 5404 56308 5460 56318
rect 5404 56214 5460 56252
rect 5292 54402 5348 54414
rect 5292 54350 5294 54402
rect 5346 54350 5348 54402
rect 5292 54068 5348 54350
rect 5292 54002 5348 54012
rect 5404 53732 5460 53742
rect 5404 53508 5460 53676
rect 5404 53442 5460 53452
rect 5516 53172 5572 57486
rect 5628 53732 5684 59052
rect 5740 55412 5796 59388
rect 5852 59220 5908 59726
rect 6748 59778 6804 59790
rect 6748 59726 6750 59778
rect 6802 59726 6804 59778
rect 6748 59444 6804 59726
rect 6748 59378 6804 59388
rect 7196 59778 7252 59790
rect 7196 59726 7198 59778
rect 7250 59726 7252 59778
rect 6412 59332 6468 59342
rect 6412 59238 6468 59276
rect 5852 59154 5908 59164
rect 7196 59220 7252 59726
rect 7196 59154 7252 59164
rect 7644 59778 7700 59836
rect 7644 59726 7646 59778
rect 7698 59726 7700 59778
rect 5964 59108 6020 59118
rect 5964 59014 6020 59052
rect 6860 59108 6916 59118
rect 7308 59108 7364 59118
rect 7644 59108 7700 59726
rect 8092 59778 8148 59790
rect 8092 59726 8094 59778
rect 8146 59726 8148 59778
rect 8092 59444 8148 59726
rect 8540 59780 8596 59790
rect 8540 59778 8932 59780
rect 8540 59726 8542 59778
rect 8594 59726 8932 59778
rect 8540 59724 8932 59726
rect 8540 59714 8596 59724
rect 8092 59378 8148 59388
rect 8876 59444 8932 59724
rect 8988 59778 9044 59790
rect 8988 59726 8990 59778
rect 9042 59726 9044 59778
rect 8988 59668 9044 59726
rect 10668 59780 10724 59790
rect 8988 59602 9044 59612
rect 10108 59668 10164 59678
rect 9884 59556 9940 59566
rect 8988 59444 9044 59454
rect 8876 59442 9044 59444
rect 8876 59390 8990 59442
rect 9042 59390 9044 59442
rect 8876 59388 9044 59390
rect 8652 59332 8708 59342
rect 8652 59238 8708 59276
rect 6860 59106 7028 59108
rect 6860 59054 6862 59106
rect 6914 59054 7028 59106
rect 6860 59052 7028 59054
rect 6860 59042 6916 59052
rect 5852 58996 5908 59006
rect 5852 57540 5908 58940
rect 6300 58772 6356 58782
rect 5964 58212 6020 58222
rect 6300 58212 6356 58716
rect 5964 58118 6020 58156
rect 6188 58210 6356 58212
rect 6188 58158 6302 58210
rect 6354 58158 6356 58210
rect 6188 58156 6356 58158
rect 5852 57538 6020 57540
rect 5852 57486 5854 57538
rect 5906 57486 6020 57538
rect 5852 57484 6020 57486
rect 5852 57474 5908 57484
rect 5852 56756 5908 56766
rect 5852 56306 5908 56700
rect 5852 56254 5854 56306
rect 5906 56254 5908 56306
rect 5852 56242 5908 56254
rect 5964 55858 6020 57484
rect 5964 55806 5966 55858
rect 6018 55806 6020 55858
rect 5964 55794 6020 55806
rect 6076 56642 6132 56654
rect 6076 56590 6078 56642
rect 6130 56590 6132 56642
rect 5852 55412 5908 55422
rect 5740 55410 5908 55412
rect 5740 55358 5854 55410
rect 5906 55358 5908 55410
rect 5740 55356 5908 55358
rect 5740 54404 5796 54414
rect 5740 54310 5796 54348
rect 5852 53954 5908 55356
rect 5852 53902 5854 53954
rect 5906 53902 5908 53954
rect 5852 53890 5908 53902
rect 6076 54628 6132 56590
rect 6188 54740 6244 58156
rect 6300 58146 6356 58156
rect 6748 58212 6804 58222
rect 6748 58118 6804 58156
rect 6412 57540 6468 57550
rect 6860 57540 6916 57550
rect 6412 57538 6580 57540
rect 6412 57486 6414 57538
rect 6466 57486 6580 57538
rect 6412 57484 6580 57486
rect 6412 57474 6468 57484
rect 6412 56644 6468 56654
rect 6412 56550 6468 56588
rect 6188 54674 6244 54684
rect 6300 55970 6356 55982
rect 6300 55918 6302 55970
rect 6354 55918 6356 55970
rect 5628 53666 5684 53676
rect 5628 53506 5684 53518
rect 5628 53454 5630 53506
rect 5682 53454 5684 53506
rect 5628 53396 5684 53454
rect 6076 53508 6132 54572
rect 6300 54404 6356 55918
rect 6412 55074 6468 55086
rect 6412 55022 6414 55074
rect 6466 55022 6468 55074
rect 6412 54628 6468 55022
rect 6412 54562 6468 54572
rect 6300 54338 6356 54348
rect 6412 54402 6468 54414
rect 6412 54350 6414 54402
rect 6466 54350 6468 54402
rect 6300 53954 6356 53966
rect 6300 53902 6302 53954
rect 6354 53902 6356 53954
rect 6076 53414 6132 53452
rect 6188 53732 6244 53742
rect 5628 53340 6020 53396
rect 5852 53172 5908 53182
rect 5516 53170 5908 53172
rect 5516 53118 5854 53170
rect 5906 53118 5908 53170
rect 5516 53116 5908 53118
rect 5404 53060 5460 53070
rect 5404 52966 5460 53004
rect 5516 52948 5572 53116
rect 5852 53106 5908 53116
rect 5516 52882 5572 52892
rect 5180 52780 5460 52836
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 4284 52274 4340 52332
rect 4284 52222 4286 52274
rect 4338 52222 4340 52274
rect 4284 52210 4340 52222
rect 4396 52276 4452 52286
rect 4060 51266 4116 51278
rect 4060 51214 4062 51266
rect 4114 51214 4116 51266
rect 4060 51156 4116 51214
rect 4060 51090 4116 51100
rect 4060 50596 4116 50606
rect 4060 50502 4116 50540
rect 3948 50418 4004 50428
rect 3836 49086 3838 49138
rect 3890 49086 3892 49138
rect 3836 49074 3892 49086
rect 3948 49812 4004 49822
rect 3948 48356 4004 49756
rect 4172 48916 4228 51548
rect 4396 51156 4452 52220
rect 5292 52276 5348 52286
rect 4844 52164 4900 52174
rect 4844 52070 4900 52108
rect 4844 51604 4900 51614
rect 4844 51510 4900 51548
rect 5292 51602 5348 52220
rect 5404 51940 5460 52780
rect 5964 52722 6020 53340
rect 5964 52670 5966 52722
rect 6018 52670 6020 52722
rect 5964 52658 6020 52670
rect 6076 52276 6132 52286
rect 6188 52276 6244 53676
rect 6300 53396 6356 53902
rect 6412 53956 6468 54350
rect 6524 54068 6580 57484
rect 6972 57540 7028 59052
rect 7308 59106 7476 59108
rect 7308 59054 7310 59106
rect 7362 59054 7476 59106
rect 7308 59052 7476 59054
rect 7308 59042 7364 59052
rect 7308 58324 7364 58334
rect 7196 57540 7252 57550
rect 6972 57538 7252 57540
rect 6972 57486 7198 57538
rect 7250 57486 7252 57538
rect 6972 57484 7252 57486
rect 6860 57446 6916 57484
rect 6748 57426 6804 57438
rect 6748 57374 6750 57426
rect 6802 57374 6804 57426
rect 6748 56084 6804 57374
rect 6972 57090 7028 57102
rect 6972 57038 6974 57090
rect 7026 57038 7028 57090
rect 6972 56978 7028 57038
rect 6972 56926 6974 56978
rect 7026 56926 7028 56978
rect 6860 56308 6916 56318
rect 6860 56214 6916 56252
rect 6748 56028 6916 56084
rect 6524 54002 6580 54012
rect 6636 55972 6692 55982
rect 6412 53890 6468 53900
rect 6524 53732 6580 53742
rect 6524 53638 6580 53676
rect 6300 53340 6468 53396
rect 6300 53172 6356 53182
rect 6300 53078 6356 53116
rect 6412 52948 6468 53340
rect 6132 52220 6244 52276
rect 6300 52892 6468 52948
rect 5628 51940 5684 51950
rect 5404 51938 5684 51940
rect 5404 51886 5630 51938
rect 5682 51886 5684 51938
rect 5404 51884 5684 51886
rect 5292 51550 5294 51602
rect 5346 51550 5348 51602
rect 5292 51538 5348 51550
rect 5404 51604 5460 51614
rect 4396 51090 4452 51100
rect 5404 51268 5460 51548
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 4508 50708 4564 50718
rect 4508 50614 4564 50652
rect 4844 50596 4900 50606
rect 4732 49924 4788 49934
rect 4732 49830 4788 49868
rect 4844 49812 4900 50540
rect 5068 50482 5124 50494
rect 5068 50430 5070 50482
rect 5122 50430 5124 50482
rect 5068 50428 5124 50430
rect 5404 50428 5460 51212
rect 5068 50372 5236 50428
rect 4956 50260 5012 50270
rect 4956 50034 5012 50204
rect 4956 49982 4958 50034
rect 5010 49982 5012 50034
rect 4956 49970 5012 49982
rect 4844 49756 5012 49812
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 4172 48850 4228 48860
rect 4956 49138 5012 49756
rect 5180 49700 5236 50372
rect 5180 49634 5236 49644
rect 5292 50372 5460 50428
rect 5068 49588 5124 49598
rect 5068 49494 5124 49532
rect 4956 49086 4958 49138
rect 5010 49086 5012 49138
rect 4620 48804 4676 48814
rect 4620 48710 4676 48748
rect 3724 47954 3780 47964
rect 3836 48300 4004 48356
rect 3836 47908 3892 48300
rect 3948 48132 4004 48142
rect 3948 48130 4228 48132
rect 3948 48078 3950 48130
rect 4002 48078 4228 48130
rect 3948 48076 4228 48078
rect 3948 48066 4004 48076
rect 4060 47908 4116 47918
rect 3836 47852 4004 47908
rect 3612 47740 3892 47796
rect 3836 47682 3892 47740
rect 3836 47630 3838 47682
rect 3890 47630 3892 47682
rect 3836 47618 3892 47630
rect 3500 47518 3502 47570
rect 3554 47518 3556 47570
rect 3500 47506 3556 47518
rect 3388 47346 3444 47358
rect 3388 47294 3390 47346
rect 3442 47294 3444 47346
rect 3388 47012 3444 47294
rect 3612 47348 3668 47358
rect 3612 47254 3668 47292
rect 3164 46956 3444 47012
rect 3948 47012 4004 47852
rect 3164 46898 3220 46956
rect 3164 46846 3166 46898
rect 3218 46846 3220 46898
rect 3164 46834 3220 46846
rect 3388 46786 3444 46798
rect 3388 46734 3390 46786
rect 3442 46734 3444 46786
rect 3276 45890 3332 45902
rect 3276 45838 3278 45890
rect 3330 45838 3332 45890
rect 3276 45668 3332 45838
rect 3276 45602 3332 45612
rect 3052 45278 3054 45330
rect 3106 45278 3108 45330
rect 2716 44324 2772 44334
rect 2716 44230 2772 44268
rect 2940 44322 2996 44334
rect 2940 44270 2942 44322
rect 2994 44270 2996 44322
rect 2940 44100 2996 44270
rect 3052 44324 3108 45278
rect 3164 45332 3220 45342
rect 3164 44434 3220 45276
rect 3388 44548 3444 46734
rect 3500 46788 3556 46798
rect 3500 46694 3556 46732
rect 3612 46228 3668 46238
rect 3612 46114 3668 46172
rect 3612 46062 3614 46114
rect 3666 46062 3668 46114
rect 3612 45444 3668 46062
rect 3612 45378 3668 45388
rect 3612 45220 3668 45230
rect 3612 44996 3668 45164
rect 3612 44994 3780 44996
rect 3612 44942 3614 44994
rect 3666 44942 3780 44994
rect 3612 44940 3780 44942
rect 3612 44930 3668 44940
rect 3388 44482 3444 44492
rect 3164 44382 3166 44434
rect 3218 44382 3220 44434
rect 3164 44370 3220 44382
rect 3052 44258 3108 44268
rect 2604 44044 2772 44100
rect 2492 43426 2548 43438
rect 2492 43374 2494 43426
rect 2546 43374 2548 43426
rect 2492 43204 2548 43374
rect 2492 42308 2548 43148
rect 2604 42868 2660 42878
rect 2604 42774 2660 42812
rect 2492 42252 2660 42308
rect 2492 42084 2548 42094
rect 2492 41990 2548 42028
rect 2268 41358 2270 41410
rect 2322 41358 2324 41410
rect 2268 40402 2324 41358
rect 2268 40350 2270 40402
rect 2322 40350 2324 40402
rect 2044 39396 2100 39406
rect 2044 39302 2100 39340
rect 2044 38836 2100 38846
rect 2268 38836 2324 40350
rect 2380 41746 2436 41758
rect 2380 41694 2382 41746
rect 2434 41694 2436 41746
rect 2380 40180 2436 41694
rect 2604 41300 2660 42252
rect 2380 40114 2436 40124
rect 2492 41244 2660 41300
rect 2716 42082 2772 44044
rect 2940 44034 2996 44044
rect 3724 44100 3780 44940
rect 3724 44034 3780 44044
rect 3500 43988 3556 43998
rect 3388 43764 3444 43774
rect 3052 43652 3108 43662
rect 3388 43652 3444 43708
rect 2940 42868 2996 42878
rect 2940 42774 2996 42812
rect 2716 42030 2718 42082
rect 2770 42030 2772 42082
rect 2044 38742 2100 38780
rect 2156 38780 2324 38836
rect 2380 39956 2436 39966
rect 2380 39058 2436 39900
rect 2380 39006 2382 39058
rect 2434 39006 2436 39058
rect 1932 38658 1988 38668
rect 1932 37828 1988 37838
rect 1932 37826 2100 37828
rect 1932 37774 1934 37826
rect 1986 37774 2100 37826
rect 1932 37772 2100 37774
rect 1932 37762 1988 37772
rect 1932 37492 1988 37502
rect 1820 37490 1988 37492
rect 1820 37438 1934 37490
rect 1986 37438 1988 37490
rect 1820 37436 1988 37438
rect 1932 37426 1988 37436
rect 1820 36706 1876 36718
rect 1820 36654 1822 36706
rect 1874 36654 1876 36706
rect 1820 36594 1876 36654
rect 1820 36542 1822 36594
rect 1874 36542 1876 36594
rect 1820 36530 1876 36542
rect 1708 36418 1764 36428
rect 1484 36372 1540 36382
rect 1372 36316 1484 36372
rect 1484 32900 1540 36316
rect 2044 35812 2100 37772
rect 2156 36036 2212 38780
rect 2268 38668 2324 38678
rect 2268 37156 2324 38612
rect 2380 38388 2436 39006
rect 2492 39730 2548 41244
rect 2604 41076 2660 41086
rect 2604 40982 2660 41020
rect 2716 40740 2772 42030
rect 3052 42082 3108 43596
rect 3276 43596 3444 43652
rect 3052 42030 3054 42082
rect 3106 42030 3108 42082
rect 3052 42018 3108 42030
rect 3164 43538 3220 43550
rect 3164 43486 3166 43538
rect 3218 43486 3220 43538
rect 2940 41858 2996 41870
rect 2940 41806 2942 41858
rect 2994 41806 2996 41858
rect 2828 41410 2884 41422
rect 2828 41358 2830 41410
rect 2882 41358 2884 41410
rect 2828 41076 2884 41358
rect 2940 41412 2996 41806
rect 3052 41412 3108 41422
rect 2940 41410 3108 41412
rect 2940 41358 3054 41410
rect 3106 41358 3108 41410
rect 2940 41356 3108 41358
rect 3052 41346 3108 41356
rect 3164 41188 3220 43486
rect 3164 41122 3220 41132
rect 3276 43204 3332 43596
rect 3276 41186 3332 43148
rect 3500 43540 3556 43932
rect 3724 43540 3780 43550
rect 3500 43538 3780 43540
rect 3500 43486 3726 43538
rect 3778 43486 3780 43538
rect 3500 43484 3780 43486
rect 3500 42868 3556 43484
rect 3724 43474 3780 43484
rect 3276 41134 3278 41186
rect 3330 41134 3332 41186
rect 3276 41122 3332 41134
rect 3388 42812 3556 42868
rect 3612 42866 3668 42878
rect 3612 42814 3614 42866
rect 3666 42814 3668 42866
rect 2828 41020 2996 41076
rect 2716 40684 2884 40740
rect 2828 40516 2884 40684
rect 2940 40626 2996 41020
rect 2940 40574 2942 40626
rect 2994 40574 2996 40626
rect 2940 40562 2996 40574
rect 2828 40450 2884 40460
rect 2716 40404 2772 40414
rect 2492 39678 2494 39730
rect 2546 39678 2548 39730
rect 2492 39060 2548 39678
rect 2604 40180 2660 40190
rect 2604 39284 2660 40124
rect 2716 39842 2772 40348
rect 3388 39956 3444 42812
rect 3500 42530 3556 42542
rect 3500 42478 3502 42530
rect 3554 42478 3556 42530
rect 3500 42420 3556 42478
rect 3500 42354 3556 42364
rect 3612 42082 3668 42814
rect 3724 42532 3780 42542
rect 3724 42438 3780 42476
rect 3948 42420 4004 46956
rect 4060 45220 4116 47852
rect 4172 47796 4228 48076
rect 4844 47908 4900 47918
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 4172 47458 4228 47740
rect 4172 47406 4174 47458
rect 4226 47406 4228 47458
rect 4172 47394 4228 47406
rect 4284 47572 4340 47582
rect 4172 46564 4228 46574
rect 4172 46470 4228 46508
rect 4284 46004 4340 47516
rect 4844 47460 4900 47852
rect 4396 47404 4900 47460
rect 4956 47460 5012 49086
rect 5292 48468 5348 50372
rect 5516 49812 5572 51884
rect 5628 51874 5684 51884
rect 5740 51604 5796 51614
rect 5740 51510 5796 51548
rect 6076 50596 6132 52220
rect 6300 51940 6356 52892
rect 6524 52276 6580 52286
rect 6636 52276 6692 55916
rect 6748 55522 6804 55534
rect 6748 55470 6750 55522
rect 6802 55470 6804 55522
rect 6748 55410 6804 55470
rect 6748 55358 6750 55410
rect 6802 55358 6804 55410
rect 6748 55346 6804 55358
rect 6748 54402 6804 54414
rect 6748 54350 6750 54402
rect 6802 54350 6804 54402
rect 6748 54180 6804 54350
rect 6748 54114 6804 54124
rect 6860 53620 6916 56028
rect 6188 51378 6244 51390
rect 6188 51326 6190 51378
rect 6242 51326 6244 51378
rect 6188 51156 6244 51326
rect 6188 50708 6244 51100
rect 6188 50642 6244 50652
rect 6300 50818 6356 51884
rect 6300 50766 6302 50818
rect 6354 50766 6356 50818
rect 6076 50530 6132 50540
rect 5852 50484 5908 50494
rect 6300 50428 6356 50766
rect 5740 50372 5796 50382
rect 5740 50278 5796 50316
rect 5628 50036 5684 50046
rect 5628 49942 5684 49980
rect 5516 49756 5684 49812
rect 5628 49364 5684 49756
rect 5068 48412 5348 48468
rect 5516 49140 5572 49150
rect 5068 47572 5124 48412
rect 5404 48354 5460 48366
rect 5404 48302 5406 48354
rect 5458 48302 5460 48354
rect 5180 48244 5236 48254
rect 5180 48242 5348 48244
rect 5180 48190 5182 48242
rect 5234 48190 5348 48242
rect 5180 48188 5348 48190
rect 5180 48178 5236 48188
rect 5068 47516 5236 47572
rect 4956 47404 5124 47460
rect 4396 47124 4452 47404
rect 4396 47058 4452 47068
rect 4620 47292 5012 47348
rect 4620 47012 4676 47292
rect 4956 47234 5012 47292
rect 4956 47182 4958 47234
rect 5010 47182 5012 47234
rect 4956 47170 5012 47182
rect 4620 46946 4676 46956
rect 4732 47068 4900 47124
rect 4732 46788 4788 47068
rect 5068 47012 5124 47404
rect 4844 47002 4900 47012
rect 4956 46956 5124 47012
rect 4844 46900 4900 46910
rect 4844 46806 4900 46844
rect 4732 46656 4788 46732
rect 4956 46786 5012 46956
rect 4956 46734 4958 46786
rect 5010 46734 5012 46786
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 4284 45948 4564 46004
rect 4396 45780 4452 45790
rect 4284 45778 4452 45780
rect 4284 45726 4398 45778
rect 4450 45726 4452 45778
rect 4284 45724 4452 45726
rect 4284 45332 4340 45724
rect 4396 45714 4452 45724
rect 4508 45780 4564 45948
rect 4956 45892 5012 46734
rect 4956 45826 5012 45836
rect 4508 45648 4564 45724
rect 4732 45668 4788 45678
rect 4732 45666 5012 45668
rect 4732 45614 4734 45666
rect 4786 45614 5012 45666
rect 4732 45612 5012 45614
rect 4732 45602 4788 45612
rect 4284 45266 4340 45276
rect 4396 45556 4452 45566
rect 4396 45330 4452 45500
rect 4396 45278 4398 45330
rect 4450 45278 4452 45330
rect 4396 45266 4452 45278
rect 4844 45332 4900 45342
rect 4172 45220 4228 45230
rect 4060 45218 4228 45220
rect 4060 45166 4174 45218
rect 4226 45166 4228 45218
rect 4060 45164 4228 45166
rect 4060 44884 4116 45164
rect 4172 45154 4228 45164
rect 4508 44996 4564 45006
rect 4508 44902 4564 44940
rect 4060 44210 4116 44828
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 4396 44548 4452 44558
rect 4284 44436 4340 44446
rect 4284 44324 4340 44380
rect 4396 44434 4452 44492
rect 4396 44382 4398 44434
rect 4450 44382 4452 44434
rect 4396 44370 4452 44382
rect 4060 44158 4062 44210
rect 4114 44158 4116 44210
rect 4060 44146 4116 44158
rect 4172 44322 4340 44324
rect 4172 44270 4286 44322
rect 4338 44270 4340 44322
rect 4172 44268 4340 44270
rect 4172 43428 4228 44268
rect 4284 44258 4340 44268
rect 4844 43652 4900 45276
rect 4956 44548 5012 45612
rect 5180 45330 5236 47516
rect 5180 45278 5182 45330
rect 5234 45278 5236 45330
rect 5068 45106 5124 45118
rect 5068 45054 5070 45106
rect 5122 45054 5124 45106
rect 5068 44996 5124 45054
rect 5068 44930 5124 44940
rect 4956 44492 5124 44548
rect 4956 44212 5012 44222
rect 4956 44118 5012 44156
rect 4844 43586 4900 43596
rect 5068 43650 5124 44492
rect 5068 43598 5070 43650
rect 5122 43598 5124 43650
rect 5068 43586 5124 43598
rect 5180 43540 5236 45278
rect 5292 45332 5348 48188
rect 5404 46900 5460 48302
rect 5404 46834 5460 46844
rect 5404 45332 5460 45342
rect 5292 45330 5460 45332
rect 5292 45278 5406 45330
rect 5458 45278 5460 45330
rect 5292 45276 5460 45278
rect 5292 43762 5348 43774
rect 5292 43710 5294 43762
rect 5346 43710 5348 43762
rect 5292 43652 5348 43710
rect 5292 43586 5348 43596
rect 5404 43650 5460 45276
rect 5404 43598 5406 43650
rect 5458 43598 5460 43650
rect 5404 43586 5460 43598
rect 5180 43474 5236 43484
rect 5516 43538 5572 49084
rect 5628 47572 5684 49308
rect 5852 49588 5908 50428
rect 6188 50372 6356 50428
rect 6412 52274 6692 52276
rect 6412 52222 6526 52274
rect 6578 52222 6692 52274
rect 6412 52220 6692 52222
rect 6748 53284 6804 53294
rect 6860 53284 6916 53564
rect 6972 55522 7028 56926
rect 6972 55470 6974 55522
rect 7026 55470 7028 55522
rect 6972 53508 7028 55470
rect 7084 55524 7140 55534
rect 7084 53842 7140 55468
rect 7196 55300 7252 57484
rect 7308 56196 7364 58268
rect 7420 57540 7476 59052
rect 7644 59042 7700 59052
rect 7756 59108 7812 59118
rect 7756 59106 8036 59108
rect 7756 59054 7758 59106
rect 7810 59054 8036 59106
rect 7756 59052 8036 59054
rect 7756 59042 7812 59052
rect 7756 58212 7812 58222
rect 7756 58210 7924 58212
rect 7756 58158 7758 58210
rect 7810 58158 7924 58210
rect 7756 58156 7924 58158
rect 7756 58146 7812 58156
rect 7644 57540 7700 57550
rect 7420 57538 7812 57540
rect 7420 57486 7646 57538
rect 7698 57486 7812 57538
rect 7420 57484 7812 57486
rect 7644 57474 7700 57484
rect 7644 56756 7700 56766
rect 7420 56644 7476 56654
rect 7420 56550 7476 56588
rect 7644 56306 7700 56700
rect 7644 56254 7646 56306
rect 7698 56254 7700 56306
rect 7644 56242 7700 56254
rect 7308 56140 7476 56196
rect 7308 55972 7364 55982
rect 7308 55878 7364 55916
rect 7196 55234 7252 55244
rect 7196 55076 7252 55086
rect 7196 54982 7252 55020
rect 7420 54852 7476 56140
rect 7644 55522 7700 55534
rect 7644 55470 7646 55522
rect 7698 55470 7700 55522
rect 7644 55410 7700 55470
rect 7644 55358 7646 55410
rect 7698 55358 7700 55410
rect 7644 55346 7700 55358
rect 7420 54786 7476 54796
rect 7532 55188 7588 55198
rect 7532 54740 7588 55132
rect 7644 54740 7700 54750
rect 7532 54738 7700 54740
rect 7532 54686 7646 54738
rect 7698 54686 7700 54738
rect 7532 54684 7700 54686
rect 7644 54674 7700 54684
rect 7308 54404 7364 54414
rect 7308 54310 7364 54348
rect 7084 53790 7086 53842
rect 7138 53790 7140 53842
rect 7084 53732 7140 53790
rect 7084 53666 7140 53676
rect 7532 53732 7588 53742
rect 7532 53638 7588 53676
rect 7196 53620 7252 53630
rect 6972 53452 7140 53508
rect 6972 53284 7028 53294
rect 6860 53228 6972 53284
rect 6748 53170 6804 53228
rect 6972 53218 7028 53228
rect 6748 53118 6750 53170
rect 6802 53118 6804 53170
rect 5740 49252 5796 49262
rect 5852 49252 5908 49532
rect 5740 49250 5908 49252
rect 5740 49198 5742 49250
rect 5794 49198 5908 49250
rect 5740 49196 5908 49198
rect 6076 49700 6132 49710
rect 6188 49700 6244 50372
rect 6076 49698 6244 49700
rect 6076 49646 6078 49698
rect 6130 49646 6244 49698
rect 6076 49644 6244 49646
rect 6300 49700 6356 49710
rect 5740 49186 5796 49196
rect 6076 49140 6132 49644
rect 5852 48802 5908 48814
rect 5852 48750 5854 48802
rect 5906 48750 5908 48802
rect 5852 48244 5908 48750
rect 5964 48802 6020 48814
rect 5964 48750 5966 48802
rect 6018 48750 6020 48802
rect 5964 48692 6020 48750
rect 6076 48804 6132 49084
rect 6076 48738 6132 48748
rect 5964 48468 6020 48636
rect 5964 48402 6020 48412
rect 5852 48178 5908 48188
rect 6188 48020 6244 48030
rect 5628 47506 5684 47516
rect 6076 47572 6132 47582
rect 6076 47458 6132 47516
rect 6076 47406 6078 47458
rect 6130 47406 6132 47458
rect 6076 47394 6132 47406
rect 5964 47348 6020 47358
rect 5628 46562 5684 46574
rect 5628 46510 5630 46562
rect 5682 46510 5684 46562
rect 5628 46340 5684 46510
rect 5628 46274 5684 46284
rect 5852 45668 5908 45678
rect 5964 45668 6020 47292
rect 5516 43486 5518 43538
rect 5570 43486 5572 43538
rect 4172 43426 4340 43428
rect 4172 43374 4174 43426
rect 4226 43374 4340 43426
rect 4172 43372 4340 43374
rect 4172 43362 4228 43372
rect 4060 43316 4116 43326
rect 4060 43222 4116 43260
rect 4060 42756 4116 42766
rect 4060 42662 4116 42700
rect 3948 42354 4004 42364
rect 3724 42196 3780 42206
rect 3724 42102 3780 42140
rect 3612 42030 3614 42082
rect 3666 42030 3668 42082
rect 3612 42018 3668 42030
rect 3948 41970 4004 41982
rect 3948 41918 3950 41970
rect 4002 41918 4004 41970
rect 3612 41412 3668 41422
rect 3612 41318 3668 41356
rect 3836 41300 3892 41310
rect 3388 39890 3444 39900
rect 3500 40516 3556 40526
rect 3500 40290 3556 40460
rect 3500 40238 3502 40290
rect 3554 40238 3556 40290
rect 2716 39790 2718 39842
rect 2770 39790 2772 39842
rect 2716 39778 2772 39790
rect 3500 39842 3556 40238
rect 3500 39790 3502 39842
rect 3554 39790 3556 39842
rect 3500 39778 3556 39790
rect 3612 39844 3668 39854
rect 3388 39732 3444 39742
rect 3388 39620 3444 39676
rect 3612 39730 3668 39788
rect 3612 39678 3614 39730
rect 3666 39678 3668 39730
rect 3612 39666 3668 39678
rect 3388 39564 3556 39620
rect 2604 39218 2660 39228
rect 3052 39394 3108 39406
rect 3052 39342 3054 39394
rect 3106 39342 3108 39394
rect 2492 39004 2772 39060
rect 2604 38834 2660 38846
rect 2604 38782 2606 38834
rect 2658 38782 2660 38834
rect 2492 38724 2548 38762
rect 2492 38658 2548 38668
rect 2380 38332 2548 38388
rect 2380 38164 2436 38174
rect 2380 38070 2436 38108
rect 2492 37268 2548 38332
rect 2604 38164 2660 38782
rect 2604 38098 2660 38108
rect 2716 37828 2772 39004
rect 3052 38836 3108 39342
rect 3276 39396 3332 39406
rect 3164 38836 3220 38846
rect 3052 38834 3220 38836
rect 3052 38782 3166 38834
rect 3218 38782 3220 38834
rect 3052 38780 3220 38782
rect 3164 38770 3220 38780
rect 2940 38724 2996 38734
rect 2940 38050 2996 38668
rect 3276 38052 3332 39340
rect 3388 38724 3444 38762
rect 3388 38658 3444 38668
rect 2940 37998 2942 38050
rect 2994 37998 2996 38050
rect 2940 37986 2996 37998
rect 3164 37996 3332 38052
rect 3500 38050 3556 39564
rect 3500 37998 3502 38050
rect 3554 37998 3556 38050
rect 3052 37938 3108 37950
rect 3052 37886 3054 37938
rect 3106 37886 3108 37938
rect 3052 37828 3108 37886
rect 2716 37772 3108 37828
rect 3164 37268 3220 37996
rect 3500 37986 3556 37998
rect 3612 39284 3668 39294
rect 3612 38946 3668 39228
rect 3836 39284 3892 41244
rect 3948 40962 4004 41918
rect 4172 41972 4228 41982
rect 4172 41878 4228 41916
rect 4284 41748 4340 43372
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4620 42530 4676 42542
rect 4620 42478 4622 42530
rect 4674 42478 4676 42530
rect 4620 42084 4676 42478
rect 4620 42018 4676 42028
rect 5068 42530 5124 42542
rect 5068 42478 5070 42530
rect 5122 42478 5124 42530
rect 4956 41860 5012 41870
rect 4956 41766 5012 41804
rect 4172 41692 4340 41748
rect 3948 40910 3950 40962
rect 4002 40910 4004 40962
rect 3948 40898 4004 40910
rect 4060 41188 4116 41198
rect 4060 39956 4116 41132
rect 3836 39218 3892 39228
rect 3948 39900 4116 39956
rect 3724 39172 3780 39182
rect 3724 39058 3780 39116
rect 3724 39006 3726 39058
rect 3778 39006 3780 39058
rect 3724 38994 3780 39006
rect 3836 39060 3892 39070
rect 3836 38966 3892 39004
rect 3612 38894 3614 38946
rect 3666 38894 3668 38946
rect 3276 37828 3332 37838
rect 3276 37734 3332 37772
rect 3612 37716 3668 38894
rect 3948 38836 4004 39900
rect 4060 39732 4116 39742
rect 4060 39638 4116 39676
rect 3612 37650 3668 37660
rect 3724 38780 4004 38836
rect 4060 39172 4116 39182
rect 3724 37492 3780 38780
rect 3836 38500 3892 38510
rect 3836 37940 3892 38444
rect 4060 38276 4116 39116
rect 4172 38500 4228 41692
rect 5068 41636 5124 42478
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 5068 41570 5124 41580
rect 5180 42196 5236 42206
rect 4476 41514 4740 41524
rect 4844 41412 4900 41422
rect 4508 41188 4564 41198
rect 4508 41094 4564 41132
rect 4732 40740 4788 40750
rect 4284 40628 4340 40638
rect 4284 40534 4340 40572
rect 4732 40626 4788 40684
rect 4732 40574 4734 40626
rect 4786 40574 4788 40626
rect 4732 40562 4788 40574
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4732 39842 4788 39854
rect 4732 39790 4734 39842
rect 4786 39790 4788 39842
rect 4620 39508 4676 39518
rect 4620 39414 4676 39452
rect 4172 38434 4228 38444
rect 4284 38948 4340 38958
rect 4060 38210 4116 38220
rect 4284 38164 4340 38892
rect 4620 38948 4676 38958
rect 4732 38948 4788 39790
rect 4844 39396 4900 41356
rect 5068 40964 5124 40974
rect 5068 40870 5124 40908
rect 4956 40516 5012 40526
rect 4956 39730 5012 40460
rect 5068 40404 5124 40442
rect 5068 40338 5124 40348
rect 4956 39678 4958 39730
rect 5010 39678 5012 39730
rect 4956 39620 5012 39678
rect 5180 39732 5236 42140
rect 5516 42084 5572 43486
rect 5404 42028 5572 42084
rect 5628 45666 6020 45668
rect 5628 45614 5854 45666
rect 5906 45614 6020 45666
rect 5628 45612 6020 45614
rect 6076 46900 6132 46910
rect 5404 39732 5460 42028
rect 5628 41972 5684 45612
rect 5852 45602 5908 45612
rect 6076 45556 6132 46844
rect 6076 45490 6132 45500
rect 6188 45332 6244 47964
rect 5852 45276 6244 45332
rect 5740 44210 5796 44222
rect 5740 44158 5742 44210
rect 5794 44158 5796 44210
rect 5740 43988 5796 44158
rect 5740 43922 5796 43932
rect 5628 41906 5684 41916
rect 5740 42420 5796 42430
rect 5516 41860 5572 41870
rect 5516 41766 5572 41804
rect 5628 41186 5684 41198
rect 5628 41134 5630 41186
rect 5682 41134 5684 41186
rect 5516 40628 5572 40638
rect 5628 40628 5684 41134
rect 5740 41188 5796 42364
rect 5852 41412 5908 45276
rect 5964 45108 6020 45118
rect 5964 44548 6020 45052
rect 6076 44994 6132 45006
rect 6076 44942 6078 44994
rect 6130 44942 6132 44994
rect 6076 44772 6132 44942
rect 6076 44706 6132 44716
rect 5964 44492 6132 44548
rect 5964 44324 6020 44334
rect 5964 44230 6020 44268
rect 6076 42756 6132 44492
rect 6188 44546 6244 45276
rect 6188 44494 6190 44546
rect 6242 44494 6244 44546
rect 6188 44482 6244 44494
rect 6300 43652 6356 49644
rect 6412 47796 6468 52220
rect 6524 52210 6580 52220
rect 6636 51828 6692 51838
rect 6636 51380 6692 51772
rect 6748 51492 6804 53118
rect 7084 53060 7140 53452
rect 7196 53170 7252 53564
rect 7196 53118 7198 53170
rect 7250 53118 7252 53170
rect 7196 53106 7252 53118
rect 6972 53004 7140 53060
rect 6860 52724 6916 52734
rect 6860 51604 6916 52668
rect 6972 52388 7028 53004
rect 6972 52274 7028 52332
rect 6972 52222 6974 52274
rect 7026 52222 7028 52274
rect 6972 52210 7028 52222
rect 7196 52948 7252 52958
rect 6860 51538 6916 51548
rect 6748 51426 6804 51436
rect 7084 51492 7140 51502
rect 6524 51378 6692 51380
rect 6524 51326 6638 51378
rect 6690 51326 6692 51378
rect 6524 51324 6692 51326
rect 6524 50260 6580 51324
rect 6636 51314 6692 51324
rect 6860 51380 6916 51390
rect 6860 51286 6916 51324
rect 6748 51266 6804 51278
rect 6748 51214 6750 51266
rect 6802 51214 6804 51266
rect 6524 50194 6580 50204
rect 6636 50594 6692 50606
rect 6636 50542 6638 50594
rect 6690 50542 6692 50594
rect 6412 47740 6580 47796
rect 6524 45890 6580 47740
rect 6636 47236 6692 50542
rect 6748 50372 6804 51214
rect 6972 50932 7028 50942
rect 6860 50708 6916 50718
rect 6860 50614 6916 50652
rect 6972 50594 7028 50876
rect 6972 50542 6974 50594
rect 7026 50542 7028 50594
rect 6972 50530 7028 50542
rect 6748 50278 6804 50316
rect 6972 49812 7028 49822
rect 7084 49812 7140 51436
rect 6860 49810 7140 49812
rect 6860 49758 6974 49810
rect 7026 49758 7140 49810
rect 6860 49756 7140 49758
rect 6748 49588 6804 49598
rect 6748 48356 6804 49532
rect 6748 48242 6804 48300
rect 6748 48190 6750 48242
rect 6802 48190 6804 48242
rect 6748 47572 6804 48190
rect 6748 47506 6804 47516
rect 6860 49476 6916 49756
rect 6972 49746 7028 49756
rect 6860 47348 6916 49420
rect 6972 49140 7028 49150
rect 6972 48914 7028 49084
rect 6972 48862 6974 48914
rect 7026 48862 7028 48914
rect 6972 47796 7028 48862
rect 7196 48804 7252 52892
rect 7308 52836 7364 52846
rect 7308 50428 7364 52780
rect 7644 52834 7700 52846
rect 7644 52782 7646 52834
rect 7698 52782 7700 52834
rect 7644 52724 7700 52782
rect 7756 52836 7812 57484
rect 7868 57426 7924 58156
rect 7868 57374 7870 57426
rect 7922 57374 7924 57426
rect 7868 57362 7924 57374
rect 7868 56642 7924 56654
rect 7868 56590 7870 56642
rect 7922 56590 7924 56642
rect 7868 56532 7924 56590
rect 7868 56466 7924 56476
rect 7756 52770 7812 52780
rect 7868 55858 7924 55870
rect 7868 55806 7870 55858
rect 7922 55806 7924 55858
rect 7868 55076 7924 55806
rect 7980 55524 8036 59052
rect 8092 59106 8148 59118
rect 8092 59054 8094 59106
rect 8146 59054 8148 59106
rect 8092 58772 8148 59054
rect 8092 58706 8148 58716
rect 8204 58210 8260 58222
rect 8204 58158 8206 58210
rect 8258 58158 8260 58210
rect 8092 57538 8148 57550
rect 8092 57486 8094 57538
rect 8146 57486 8148 57538
rect 8092 57426 8148 57486
rect 8092 57374 8094 57426
rect 8146 57374 8148 57426
rect 8092 56868 8148 57374
rect 8204 57316 8260 58158
rect 8652 58210 8708 58222
rect 8652 58158 8654 58210
rect 8706 58158 8708 58210
rect 8652 57764 8708 58158
rect 8652 57698 8708 57708
rect 8764 57876 8820 57886
rect 8204 57250 8260 57260
rect 8428 57540 8484 57550
rect 8092 56802 8148 56812
rect 8204 57092 8260 57102
rect 8204 56978 8260 57036
rect 8204 56926 8206 56978
rect 8258 56926 8260 56978
rect 7980 55458 8036 55468
rect 8092 56644 8148 56654
rect 8092 56084 8148 56588
rect 8092 55300 8148 56028
rect 8204 55522 8260 56926
rect 8204 55470 8206 55522
rect 8258 55470 8260 55522
rect 8204 55458 8260 55470
rect 8092 55234 8148 55244
rect 7644 52658 7700 52668
rect 7644 51940 7700 51950
rect 7868 51940 7924 55020
rect 8092 55076 8148 55114
rect 8092 55010 8148 55020
rect 8092 54852 8148 54862
rect 7980 53508 8036 53518
rect 7980 53414 8036 53452
rect 8092 53060 8148 54796
rect 8428 54740 8484 57484
rect 8540 57538 8596 57550
rect 8540 57486 8542 57538
rect 8594 57486 8596 57538
rect 8540 57428 8596 57486
rect 8540 57296 8596 57372
rect 8764 56978 8820 57820
rect 8764 56926 8766 56978
rect 8818 56926 8820 56978
rect 8764 56756 8820 56926
rect 8764 56690 8820 56700
rect 8540 56420 8596 56430
rect 8540 56306 8596 56364
rect 8876 56420 8932 59388
rect 8988 59378 9044 59388
rect 9772 59332 9828 59342
rect 9324 59108 9380 59118
rect 9660 59108 9716 59118
rect 9380 59106 9716 59108
rect 9380 59054 9662 59106
rect 9714 59054 9716 59106
rect 9380 59052 9716 59054
rect 9100 58324 9156 58334
rect 9100 58230 9156 58268
rect 8876 56354 8932 56364
rect 8988 58100 9044 58110
rect 8988 57874 9044 58044
rect 8988 57822 8990 57874
rect 9042 57822 9044 57874
rect 8540 56254 8542 56306
rect 8594 56254 8596 56306
rect 8540 56242 8596 56254
rect 8988 56308 9044 57822
rect 8988 56242 9044 56252
rect 9212 56642 9268 56654
rect 9212 56590 9214 56642
rect 9266 56590 9268 56642
rect 9212 56196 9268 56590
rect 8540 56084 8596 56094
rect 8540 55410 8596 56028
rect 8988 55972 9044 55982
rect 8988 55970 9156 55972
rect 8988 55918 8990 55970
rect 9042 55918 9156 55970
rect 8988 55916 9156 55918
rect 8988 55906 9044 55916
rect 8540 55358 8542 55410
rect 8594 55358 8596 55410
rect 8540 55346 8596 55358
rect 8876 55522 8932 55534
rect 8876 55470 8878 55522
rect 8930 55470 8932 55522
rect 8764 55300 8820 55310
rect 8540 54740 8596 54750
rect 8428 54738 8708 54740
rect 8428 54686 8542 54738
rect 8594 54686 8708 54738
rect 8428 54684 8708 54686
rect 8540 54674 8596 54684
rect 8204 54404 8260 54414
rect 8204 54402 8372 54404
rect 8204 54350 8206 54402
rect 8258 54350 8372 54402
rect 8204 54348 8372 54350
rect 8204 54338 8260 54348
rect 8316 53506 8372 54348
rect 8316 53454 8318 53506
rect 8370 53454 8372 53506
rect 8092 53004 8260 53060
rect 7644 51938 7924 51940
rect 7644 51886 7646 51938
rect 7698 51886 7924 51938
rect 7644 51884 7924 51886
rect 8092 52836 8148 52846
rect 8092 52274 8148 52780
rect 8092 52222 8094 52274
rect 8146 52222 8148 52274
rect 7644 51828 7700 51884
rect 7644 51762 7700 51772
rect 7532 51378 7588 51390
rect 7532 51326 7534 51378
rect 7586 51326 7588 51378
rect 7308 50372 7476 50428
rect 7308 49700 7364 49710
rect 7308 49606 7364 49644
rect 7308 49140 7364 49150
rect 7308 49046 7364 49084
rect 6972 47730 7028 47740
rect 7084 48802 7252 48804
rect 7084 48750 7198 48802
rect 7250 48750 7252 48802
rect 7084 48748 7252 48750
rect 6860 47282 6916 47292
rect 7084 47458 7140 48748
rect 7196 48738 7252 48748
rect 7420 48802 7476 50372
rect 7420 48750 7422 48802
rect 7474 48750 7476 48802
rect 7420 48692 7476 48750
rect 7308 48636 7420 48692
rect 7308 47570 7364 48636
rect 7420 48626 7476 48636
rect 7532 48468 7588 51326
rect 7756 51378 7812 51390
rect 7756 51326 7758 51378
rect 7810 51326 7812 51378
rect 7756 51268 7812 51326
rect 7980 51378 8036 51390
rect 7980 51326 7982 51378
rect 8034 51326 8036 51378
rect 7756 51202 7812 51212
rect 7868 51266 7924 51278
rect 7868 51214 7870 51266
rect 7922 51214 7924 51266
rect 7644 50932 7700 50942
rect 7644 50708 7700 50876
rect 7868 50932 7924 51214
rect 7868 50866 7924 50876
rect 7756 50708 7812 50718
rect 7644 50706 7812 50708
rect 7644 50654 7758 50706
rect 7810 50654 7812 50706
rect 7644 50652 7812 50654
rect 7756 50642 7812 50652
rect 7980 50708 8036 51326
rect 7980 50642 8036 50652
rect 7868 50596 7924 50606
rect 7644 50484 7700 50522
rect 7644 50418 7700 50428
rect 7868 50482 7924 50540
rect 7868 50430 7870 50482
rect 7922 50430 7924 50482
rect 7868 50418 7924 50430
rect 7980 50372 8036 50382
rect 7980 49922 8036 50316
rect 7980 49870 7982 49922
rect 8034 49870 8036 49922
rect 7980 49858 8036 49870
rect 7868 48804 7924 48814
rect 7868 48710 7924 48748
rect 7308 47518 7310 47570
rect 7362 47518 7364 47570
rect 7308 47506 7364 47518
rect 7420 48412 7588 48468
rect 7084 47406 7086 47458
rect 7138 47406 7140 47458
rect 6636 47180 6804 47236
rect 6636 46788 6692 46798
rect 6636 46694 6692 46732
rect 6748 46002 6804 47180
rect 6748 45950 6750 46002
rect 6802 45950 6804 46002
rect 6748 45938 6804 45950
rect 6860 46898 6916 46910
rect 6860 46846 6862 46898
rect 6914 46846 6916 46898
rect 6524 45838 6526 45890
rect 6578 45838 6580 45890
rect 6412 44996 6468 45006
rect 6412 44322 6468 44940
rect 6412 44270 6414 44322
rect 6466 44270 6468 44322
rect 6412 43988 6468 44270
rect 6412 43922 6468 43932
rect 6524 43764 6580 45838
rect 6636 45892 6692 45902
rect 6860 45892 6916 46846
rect 6972 46674 7028 46686
rect 6972 46622 6974 46674
rect 7026 46622 7028 46674
rect 6972 46452 7028 46622
rect 6972 46386 7028 46396
rect 7084 46116 7140 47406
rect 7196 46676 7252 46686
rect 7196 46582 7252 46620
rect 7420 46452 7476 48412
rect 7532 48242 7588 48254
rect 7532 48190 7534 48242
rect 7586 48190 7588 48242
rect 7532 47570 7588 48190
rect 7868 48020 7924 48030
rect 7532 47518 7534 47570
rect 7586 47518 7588 47570
rect 7532 47506 7588 47518
rect 7756 47572 7812 47582
rect 7644 47460 7700 47470
rect 7644 47366 7700 47404
rect 7084 46050 7140 46060
rect 7196 46396 7476 46452
rect 7532 47012 7588 47022
rect 6860 45836 7028 45892
rect 6636 45798 6692 45836
rect 6748 45780 6804 45790
rect 6636 45108 6692 45118
rect 6636 45014 6692 45052
rect 6748 44660 6804 45724
rect 6860 45668 6916 45678
rect 6860 45574 6916 45612
rect 6972 45444 7028 45836
rect 7084 45778 7140 45790
rect 7084 45726 7086 45778
rect 7138 45726 7140 45778
rect 7084 45556 7140 45726
rect 7084 45490 7140 45500
rect 6860 45388 7028 45444
rect 6860 45106 6916 45388
rect 7196 45330 7252 46396
rect 7532 46340 7588 46956
rect 7644 46788 7700 46798
rect 7644 46694 7700 46732
rect 7308 46284 7588 46340
rect 7308 46004 7364 46284
rect 7756 46228 7812 47516
rect 7308 45938 7364 45948
rect 7420 46172 7812 46228
rect 7868 46676 7924 47964
rect 8092 47012 8148 52222
rect 8204 51828 8260 53004
rect 8316 52836 8372 53454
rect 8540 52836 8596 52846
rect 8316 52770 8372 52780
rect 8428 52834 8596 52836
rect 8428 52782 8542 52834
rect 8594 52782 8596 52834
rect 8428 52780 8596 52782
rect 8204 51380 8260 51772
rect 8204 51314 8260 51324
rect 8428 52722 8484 52780
rect 8540 52770 8596 52780
rect 8428 52670 8430 52722
rect 8482 52670 8484 52722
rect 8428 50372 8484 52670
rect 8540 52276 8596 52286
rect 8540 52182 8596 52220
rect 8652 51940 8708 54684
rect 8764 53842 8820 55244
rect 8764 53790 8766 53842
rect 8818 53790 8820 53842
rect 8764 53778 8820 53790
rect 8876 53732 8932 55470
rect 9100 55188 9156 55916
rect 8988 55076 9044 55086
rect 8988 54982 9044 55020
rect 8876 53666 8932 53676
rect 8988 54740 9044 54750
rect 9100 54740 9156 55132
rect 8988 54738 9156 54740
rect 8988 54686 8990 54738
rect 9042 54686 9156 54738
rect 8988 54684 9156 54686
rect 8988 53620 9044 54684
rect 9212 53956 9268 56140
rect 8988 53554 9044 53564
rect 9100 53900 9268 53956
rect 8988 53172 9044 53182
rect 9100 53172 9156 53900
rect 9212 53732 9268 53742
rect 9212 53638 9268 53676
rect 8988 53170 9100 53172
rect 8988 53118 8990 53170
rect 9042 53118 9100 53170
rect 8988 53116 9100 53118
rect 8988 53106 9044 53116
rect 9100 53040 9156 53116
rect 9100 52164 9156 52174
rect 9100 52070 9156 52108
rect 8652 51884 8820 51940
rect 8652 51380 8708 51390
rect 8652 51286 8708 51324
rect 8428 50306 8484 50316
rect 8652 50596 8708 50606
rect 8316 50036 8372 50046
rect 8652 50036 8708 50540
rect 8316 49942 8372 49980
rect 8428 49980 8708 50036
rect 8764 50482 8820 51884
rect 8876 51490 8932 51502
rect 8876 51438 8878 51490
rect 8930 51438 8932 51490
rect 8876 51268 8932 51438
rect 8876 51202 8932 51212
rect 8988 51378 9044 51390
rect 8988 51326 8990 51378
rect 9042 51326 9044 51378
rect 8988 50708 9044 51326
rect 9324 51268 9380 59052
rect 9660 59042 9716 59052
rect 9436 58324 9492 58334
rect 9436 58210 9492 58268
rect 9436 58158 9438 58210
rect 9490 58158 9492 58210
rect 9436 57428 9492 58158
rect 9436 57362 9492 57372
rect 9772 56868 9828 59276
rect 9884 58324 9940 59500
rect 10108 59442 10164 59612
rect 10108 59390 10110 59442
rect 10162 59390 10164 59442
rect 10108 59378 10164 59390
rect 10668 59332 10724 59724
rect 11004 59442 11060 59948
rect 11340 59938 11396 59948
rect 14588 60002 14644 60014
rect 14588 59950 14590 60002
rect 14642 59950 14644 60002
rect 14364 59892 14420 59902
rect 12348 59780 12404 59790
rect 12348 59686 12404 59724
rect 12908 59778 12964 59790
rect 12908 59726 12910 59778
rect 12962 59726 12964 59778
rect 12460 59668 12516 59678
rect 11004 59390 11006 59442
rect 11058 59390 11060 59442
rect 11004 59378 11060 59390
rect 11564 59444 11620 59454
rect 10668 59200 10724 59276
rect 11004 59220 11060 59230
rect 9884 58230 9940 58268
rect 10780 59108 10836 59118
rect 10444 58212 10500 58222
rect 10444 58210 10612 58212
rect 10444 58158 10446 58210
rect 10498 58158 10612 58210
rect 10444 58156 10612 58158
rect 10444 58146 10500 58156
rect 9996 57652 10052 57662
rect 9996 57558 10052 57596
rect 10444 57652 10500 57662
rect 10444 57558 10500 57596
rect 10332 57316 10388 57326
rect 9772 56812 9940 56868
rect 9772 56642 9828 56654
rect 9772 56590 9774 56642
rect 9826 56590 9828 56642
rect 9772 55188 9828 56590
rect 9772 55122 9828 55132
rect 9548 55074 9604 55086
rect 9548 55022 9550 55074
rect 9602 55022 9604 55074
rect 9548 53844 9604 55022
rect 9660 55076 9716 55086
rect 9660 54404 9716 55020
rect 9660 54402 9828 54404
rect 9660 54350 9662 54402
rect 9714 54350 9828 54402
rect 9660 54348 9828 54350
rect 9660 54338 9716 54348
rect 9772 54292 9828 54348
rect 9772 54226 9828 54236
rect 9548 53778 9604 53788
rect 9660 54180 9716 54190
rect 9884 54180 9940 56812
rect 10220 56642 10276 56654
rect 10220 56590 10222 56642
rect 10274 56590 10276 56642
rect 9996 56196 10052 56206
rect 9996 56102 10052 56140
rect 10108 55300 10164 55310
rect 9996 55188 10052 55198
rect 9996 55094 10052 55132
rect 10108 54964 10164 55244
rect 10220 55076 10276 56590
rect 10220 55010 10276 55020
rect 10108 54898 10164 54908
rect 10332 54740 10388 57260
rect 10556 57204 10612 58156
rect 10780 58210 10836 59052
rect 10780 58158 10782 58210
rect 10834 58158 10836 58210
rect 10780 58100 10836 58158
rect 10780 58034 10836 58044
rect 10892 57540 10948 57550
rect 10556 57138 10612 57148
rect 10780 57538 10948 57540
rect 10780 57486 10894 57538
rect 10946 57486 10948 57538
rect 10780 57484 10948 57486
rect 10668 56642 10724 56654
rect 10668 56590 10670 56642
rect 10722 56590 10724 56642
rect 10444 55970 10500 55982
rect 10444 55918 10446 55970
rect 10498 55918 10500 55970
rect 10444 55300 10500 55918
rect 10668 55522 10724 56590
rect 10780 56196 10836 57484
rect 10892 57474 10948 57484
rect 10780 56130 10836 56140
rect 10668 55470 10670 55522
rect 10722 55470 10724 55522
rect 10668 55412 10724 55470
rect 10668 55346 10724 55356
rect 11004 56082 11060 59164
rect 11228 58658 11284 58670
rect 11228 58606 11230 58658
rect 11282 58606 11284 58658
rect 11228 57538 11284 58606
rect 11340 58210 11396 58222
rect 11340 58158 11342 58210
rect 11394 58158 11396 58210
rect 11340 57764 11396 58158
rect 11340 57698 11396 57708
rect 11228 57486 11230 57538
rect 11282 57486 11284 57538
rect 11116 57090 11172 57102
rect 11116 57038 11118 57090
rect 11170 57038 11172 57090
rect 11116 56868 11172 57038
rect 11116 56774 11172 56812
rect 11228 56532 11284 57486
rect 11564 57428 11620 59388
rect 11900 59106 11956 59118
rect 11900 59054 11902 59106
rect 11954 59054 11956 59106
rect 11788 58772 11844 58782
rect 11564 57362 11620 57372
rect 11676 58212 11732 58222
rect 11676 57316 11732 58156
rect 11676 57250 11732 57260
rect 11564 56644 11620 56654
rect 11564 56550 11620 56588
rect 11116 56308 11172 56318
rect 11116 56214 11172 56252
rect 11004 56030 11006 56082
rect 11058 56030 11060 56082
rect 11004 55412 11060 56030
rect 11228 55412 11284 56476
rect 11340 56084 11396 56094
rect 11340 55990 11396 56028
rect 11788 55972 11844 58716
rect 11900 58658 11956 59054
rect 12348 59108 12404 59118
rect 12348 59014 12404 59052
rect 11900 58606 11902 58658
rect 11954 58606 11956 58658
rect 11900 58594 11956 58606
rect 12124 58996 12180 59006
rect 12124 58546 12180 58940
rect 12124 58494 12126 58546
rect 12178 58494 12180 58546
rect 12124 58482 12180 58494
rect 12012 57538 12068 57550
rect 12012 57486 12014 57538
rect 12066 57486 12068 57538
rect 12012 57092 12068 57486
rect 12348 57538 12404 57550
rect 12348 57486 12350 57538
rect 12402 57486 12404 57538
rect 12348 57204 12404 57486
rect 12348 57138 12404 57148
rect 12012 57026 12068 57036
rect 12348 56868 12404 56878
rect 12012 56866 12404 56868
rect 12012 56814 12350 56866
rect 12402 56814 12404 56866
rect 12012 56812 12404 56814
rect 11900 56642 11956 56654
rect 11900 56590 11902 56642
rect 11954 56590 11956 56642
rect 11900 56196 11956 56590
rect 11900 56130 11956 56140
rect 11788 55906 11844 55916
rect 11900 55972 11956 55982
rect 12012 55972 12068 56812
rect 12348 56802 12404 56812
rect 12124 56084 12180 56094
rect 12124 55990 12180 56028
rect 11900 55970 12068 55972
rect 11900 55918 11902 55970
rect 11954 55918 12068 55970
rect 11900 55916 12068 55918
rect 11004 55346 11060 55356
rect 11116 55356 11284 55412
rect 11452 55860 11508 55870
rect 10444 55234 10500 55244
rect 10444 55074 10500 55086
rect 10444 55022 10446 55074
rect 10498 55022 10500 55074
rect 10444 54964 10500 55022
rect 10892 55076 10948 55086
rect 11116 55076 11172 55356
rect 10892 55074 11172 55076
rect 10892 55022 10894 55074
rect 10946 55022 11172 55074
rect 10892 55020 11172 55022
rect 11228 55188 11284 55198
rect 11228 55076 11284 55132
rect 11340 55076 11396 55086
rect 11228 55074 11396 55076
rect 11228 55022 11342 55074
rect 11394 55022 11396 55074
rect 11228 55020 11396 55022
rect 10892 54964 10948 55020
rect 10444 54908 10948 54964
rect 10556 54740 10612 54750
rect 10388 54738 10612 54740
rect 10388 54686 10558 54738
rect 10610 54686 10612 54738
rect 10388 54684 10612 54686
rect 10108 54628 10164 54638
rect 10332 54608 10388 54684
rect 9884 54124 10052 54180
rect 9660 53842 9716 54124
rect 9660 53790 9662 53842
rect 9714 53790 9716 53842
rect 9660 53778 9716 53790
rect 9884 53172 9940 53182
rect 9884 53078 9940 53116
rect 9436 52724 9492 52734
rect 9436 52274 9492 52668
rect 9436 52222 9438 52274
rect 9490 52222 9492 52274
rect 9436 52210 9492 52222
rect 9996 52276 10052 54124
rect 10108 53730 10164 54572
rect 10220 54404 10276 54414
rect 10220 54310 10276 54348
rect 10556 54292 10612 54684
rect 10556 54226 10612 54236
rect 10892 54290 10948 54908
rect 10892 54238 10894 54290
rect 10946 54238 10948 54290
rect 10892 54226 10948 54238
rect 11116 54402 11172 54414
rect 11116 54350 11118 54402
rect 11170 54350 11172 54402
rect 10444 54068 10500 54078
rect 10108 53678 10110 53730
rect 10162 53678 10164 53730
rect 10108 53172 10164 53678
rect 10108 53106 10164 53116
rect 10332 53732 10388 53742
rect 10332 53170 10388 53676
rect 10332 53118 10334 53170
rect 10386 53118 10388 53170
rect 10332 53106 10388 53118
rect 9324 51202 9380 51212
rect 8988 50642 9044 50652
rect 9772 51156 9828 51166
rect 9100 50596 9156 50634
rect 9100 50530 9156 50540
rect 8764 50430 8766 50482
rect 8818 50430 8820 50482
rect 8316 49810 8372 49822
rect 8316 49758 8318 49810
rect 8370 49758 8372 49810
rect 8316 49700 8372 49758
rect 8316 49634 8372 49644
rect 8428 49140 8484 49980
rect 8092 46946 8148 46956
rect 8204 49084 8484 49140
rect 8540 49810 8596 49822
rect 8540 49758 8542 49810
rect 8594 49758 8596 49810
rect 8540 49140 8596 49758
rect 7196 45278 7198 45330
rect 7250 45278 7252 45330
rect 7196 45266 7252 45278
rect 7196 45108 7252 45118
rect 6860 45054 6862 45106
rect 6914 45054 6916 45106
rect 6860 45042 6916 45054
rect 6972 45106 7252 45108
rect 6972 45054 7198 45106
rect 7250 45054 7252 45106
rect 6972 45052 7252 45054
rect 6524 43698 6580 43708
rect 6636 44604 6804 44660
rect 6076 42624 6132 42700
rect 6188 43596 6356 43652
rect 5964 41858 6020 41870
rect 5964 41806 5966 41858
rect 6018 41806 6020 41858
rect 5964 41748 6020 41806
rect 5964 41682 6020 41692
rect 5852 41346 5908 41356
rect 5740 41132 6020 41188
rect 5516 40626 5684 40628
rect 5516 40574 5518 40626
rect 5570 40574 5684 40626
rect 5516 40572 5684 40574
rect 5516 40562 5572 40572
rect 5740 40514 5796 40526
rect 5740 40462 5742 40514
rect 5794 40462 5796 40514
rect 5740 39956 5796 40462
rect 5852 40402 5908 40414
rect 5852 40350 5854 40402
rect 5906 40350 5908 40402
rect 5852 40292 5908 40350
rect 5852 40226 5908 40236
rect 5964 40068 6020 41132
rect 6076 41076 6132 41086
rect 6076 40982 6132 41020
rect 5740 39890 5796 39900
rect 5852 40012 6020 40068
rect 5628 39732 5684 39742
rect 5404 39730 5684 39732
rect 5404 39678 5630 39730
rect 5682 39678 5684 39730
rect 5404 39676 5684 39678
rect 5180 39666 5236 39676
rect 4956 39554 5012 39564
rect 5180 39396 5236 39406
rect 4844 39340 5012 39396
rect 4844 38948 4900 38958
rect 4732 38892 4844 38948
rect 4620 38854 4676 38892
rect 4844 38854 4900 38892
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4620 38276 4676 38286
rect 4284 38108 4452 38164
rect 4060 38052 4116 38062
rect 4060 37958 4116 37996
rect 3948 37940 4004 37950
rect 3836 37938 4004 37940
rect 3836 37886 3950 37938
rect 4002 37886 4004 37938
rect 3836 37884 4004 37886
rect 3612 37436 3780 37492
rect 3276 37268 3332 37278
rect 2492 37212 2772 37268
rect 3164 37266 3332 37268
rect 3164 37214 3278 37266
rect 3330 37214 3332 37266
rect 3164 37212 3332 37214
rect 2268 37090 2324 37100
rect 2380 37154 2436 37166
rect 2380 37102 2382 37154
rect 2434 37102 2436 37154
rect 2380 36706 2436 37102
rect 2380 36654 2382 36706
rect 2434 36654 2436 36706
rect 2268 36260 2324 36270
rect 2268 36166 2324 36204
rect 2156 35980 2324 36036
rect 2044 35746 2100 35756
rect 2156 35588 2212 35598
rect 2044 35586 2212 35588
rect 2044 35534 2158 35586
rect 2210 35534 2212 35586
rect 2044 35532 2212 35534
rect 1820 35140 1876 35150
rect 1820 35026 1876 35084
rect 1820 34974 1822 35026
rect 1874 34974 1876 35026
rect 1820 34962 1876 34974
rect 1484 32834 1540 32844
rect 1596 34804 1652 34814
rect 1484 30772 1540 30782
rect 1484 23492 1540 30716
rect 1596 24052 1652 34748
rect 2044 34468 2100 35532
rect 2156 35522 2212 35532
rect 2268 35364 2324 35980
rect 2044 34402 2100 34412
rect 2156 35308 2324 35364
rect 1932 34020 1988 34030
rect 1932 33926 1988 33964
rect 2156 34020 2212 35308
rect 2380 35252 2436 36654
rect 2380 35186 2436 35196
rect 2492 37044 2548 37054
rect 2380 35028 2436 35038
rect 2492 35028 2548 36988
rect 2380 35026 2548 35028
rect 2380 34974 2382 35026
rect 2434 34974 2548 35026
rect 2380 34972 2548 34974
rect 2604 35586 2660 35598
rect 2604 35534 2606 35586
rect 2658 35534 2660 35586
rect 2380 34962 2436 34972
rect 2380 34692 2436 34702
rect 2156 33954 2212 33964
rect 2268 34244 2324 34254
rect 2268 33458 2324 34188
rect 2268 33406 2270 33458
rect 2322 33406 2324 33458
rect 2268 33394 2324 33406
rect 1932 32900 1988 32910
rect 1932 32786 1988 32844
rect 2380 32788 2436 34636
rect 1932 32734 1934 32786
rect 1986 32734 1988 32786
rect 1932 32722 1988 32734
rect 2044 32786 2436 32788
rect 2044 32734 2382 32786
rect 2434 32734 2436 32786
rect 2044 32732 2436 32734
rect 2044 32002 2100 32732
rect 2380 32722 2436 32732
rect 2492 34018 2548 34030
rect 2492 33966 2494 34018
rect 2546 33966 2548 34018
rect 2492 32788 2548 33966
rect 2492 32722 2548 32732
rect 2604 32452 2660 35534
rect 2044 31950 2046 32002
rect 2098 31950 2100 32002
rect 2044 31938 2100 31950
rect 2268 32396 2660 32452
rect 2716 32452 2772 37212
rect 3276 37202 3332 37212
rect 3052 37156 3108 37166
rect 3052 37062 3108 37100
rect 3500 37154 3556 37166
rect 3500 37102 3502 37154
rect 3554 37102 3556 37154
rect 2940 36596 2996 36606
rect 2828 36484 2884 36494
rect 2828 36390 2884 36428
rect 2828 34692 2884 34702
rect 2828 34598 2884 34636
rect 2940 34242 2996 36540
rect 2940 34190 2942 34242
rect 2994 34190 2996 34242
rect 2940 34178 2996 34190
rect 3276 36484 3332 36494
rect 3276 35924 3332 36428
rect 2828 33124 2884 33134
rect 3276 33124 3332 35868
rect 3388 36148 3444 36158
rect 3388 35698 3444 36092
rect 3388 35646 3390 35698
rect 3442 35646 3444 35698
rect 3388 35634 3444 35646
rect 3500 35586 3556 37102
rect 3612 36484 3668 37436
rect 3836 37380 3892 37390
rect 3836 37286 3892 37324
rect 3724 37266 3780 37278
rect 3724 37214 3726 37266
rect 3778 37214 3780 37266
rect 3724 37044 3780 37214
rect 3948 37268 4004 37884
rect 4284 37940 4340 37950
rect 4284 37846 4340 37884
rect 4172 37828 4228 37838
rect 3948 37202 4004 37212
rect 4060 37716 4116 37726
rect 3724 36978 3780 36988
rect 3612 36428 3780 36484
rect 3724 35700 3780 36428
rect 4060 36482 4116 37660
rect 4060 36430 4062 36482
rect 4114 36430 4116 36482
rect 3948 36372 4004 36382
rect 3948 36278 4004 36316
rect 3836 36258 3892 36270
rect 3836 36206 3838 36258
rect 3890 36206 3892 36258
rect 3836 36148 3892 36206
rect 3836 36082 3892 36092
rect 3724 35644 3892 35700
rect 3500 35534 3502 35586
rect 3554 35534 3556 35586
rect 3500 35522 3556 35534
rect 3724 35476 3780 35486
rect 3724 35382 3780 35420
rect 3500 35252 3556 35262
rect 3388 34916 3444 34926
rect 3388 34822 3444 34860
rect 3500 34914 3556 35196
rect 3500 34862 3502 34914
rect 3554 34862 3556 34914
rect 3500 34356 3556 34862
rect 3836 34802 3892 35644
rect 4060 35028 4116 36430
rect 4172 35698 4228 37772
rect 4396 37604 4452 38108
rect 4508 37938 4564 37950
rect 4508 37886 4510 37938
rect 4562 37886 4564 37938
rect 4508 37716 4564 37886
rect 4508 37650 4564 37660
rect 4284 37548 4452 37604
rect 4284 36708 4340 37548
rect 4396 37380 4452 37390
rect 4620 37380 4676 38220
rect 4396 37378 4676 37380
rect 4396 37326 4398 37378
rect 4450 37326 4676 37378
rect 4396 37324 4676 37326
rect 4396 37314 4452 37324
rect 4620 37156 4676 37324
rect 4732 37268 4788 37278
rect 4956 37268 5012 39340
rect 5180 38946 5236 39340
rect 5516 39172 5572 39676
rect 5628 39666 5684 39676
rect 5516 39106 5572 39116
rect 5180 38894 5182 38946
rect 5234 38894 5236 38946
rect 5180 38882 5236 38894
rect 5068 38722 5124 38734
rect 5628 38724 5684 38734
rect 5068 38670 5070 38722
rect 5122 38670 5124 38722
rect 5068 38388 5124 38670
rect 5068 38322 5124 38332
rect 5516 38668 5628 38724
rect 5068 38164 5124 38202
rect 5068 38098 5124 38108
rect 4732 37266 5012 37268
rect 4732 37214 4734 37266
rect 4786 37214 5012 37266
rect 4732 37212 5012 37214
rect 4732 37202 4788 37212
rect 4620 37090 4676 37100
rect 4732 37044 4788 37054
rect 4732 37042 4900 37044
rect 4732 36990 4734 37042
rect 4786 36990 4900 37042
rect 4732 36988 4900 36990
rect 4732 36978 4788 36988
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4284 36652 4564 36708
rect 4172 35646 4174 35698
rect 4226 35646 4228 35698
rect 4172 35634 4228 35646
rect 4508 36482 4564 36652
rect 4508 36430 4510 36482
rect 4562 36430 4564 36482
rect 4508 35476 4564 36430
rect 4844 36370 4900 36988
rect 4844 36318 4846 36370
rect 4898 36318 4900 36370
rect 4844 36306 4900 36318
rect 4732 35700 4788 35710
rect 4732 35606 4788 35644
rect 4508 35420 4900 35476
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 3836 34750 3838 34802
rect 3890 34750 3892 34802
rect 3500 34300 3780 34356
rect 3500 34130 3556 34142
rect 3500 34078 3502 34130
rect 3554 34078 3556 34130
rect 3388 33572 3444 33582
rect 3388 33346 3444 33516
rect 3388 33294 3390 33346
rect 3442 33294 3444 33346
rect 3388 33282 3444 33294
rect 3500 33348 3556 34078
rect 3724 34132 3780 34300
rect 3500 33282 3556 33292
rect 3612 33684 3668 33694
rect 3276 33068 3444 33124
rect 2828 33030 2884 33068
rect 2940 32452 2996 32462
rect 2716 32396 2940 32452
rect 2268 31892 2324 32396
rect 2940 32358 2996 32396
rect 3388 32450 3444 33068
rect 3388 32398 3390 32450
rect 3442 32398 3444 32450
rect 3388 32340 3444 32398
rect 3388 32274 3444 32284
rect 3612 32228 3668 33628
rect 3500 32172 3668 32228
rect 1932 31556 1988 31566
rect 1708 31554 1988 31556
rect 1708 31502 1934 31554
rect 1986 31502 1988 31554
rect 1708 31500 1988 31502
rect 1708 26516 1764 31500
rect 1932 31490 1988 31500
rect 2044 31556 2100 31566
rect 1932 30882 1988 30894
rect 1932 30830 1934 30882
rect 1986 30830 1988 30882
rect 1708 26450 1764 26460
rect 1820 29986 1876 29998
rect 1820 29934 1822 29986
rect 1874 29934 1876 29986
rect 1596 23986 1652 23996
rect 1820 25620 1876 29934
rect 1932 29876 1988 30830
rect 1932 29810 1988 29820
rect 2044 28754 2100 31500
rect 2268 31220 2324 31836
rect 2380 32004 2436 32014
rect 2380 31890 2436 31948
rect 2380 31838 2382 31890
rect 2434 31838 2436 31890
rect 2380 31826 2436 31838
rect 2492 32002 2548 32014
rect 2492 31950 2494 32002
rect 2546 31950 2548 32002
rect 2380 31220 2436 31230
rect 2268 31218 2436 31220
rect 2268 31166 2382 31218
rect 2434 31166 2436 31218
rect 2268 31164 2436 31166
rect 2380 31154 2436 31164
rect 2492 31220 2548 31950
rect 3500 32004 3556 32172
rect 3724 32116 3780 34076
rect 3836 33684 3892 34750
rect 3836 33618 3892 33628
rect 3948 34972 4116 35028
rect 4396 35028 4452 35038
rect 3948 33460 4004 34972
rect 4396 34934 4452 34972
rect 4060 34804 4116 34814
rect 4060 34802 4228 34804
rect 4060 34750 4062 34802
rect 4114 34750 4228 34802
rect 4060 34748 4228 34750
rect 4060 34738 4116 34748
rect 4172 34356 4228 34748
rect 4284 34802 4340 34814
rect 4284 34750 4286 34802
rect 4338 34750 4340 34802
rect 4284 34468 4340 34750
rect 4844 34804 4900 35420
rect 4956 35364 5012 37212
rect 5068 37940 5124 37950
rect 5068 36932 5124 37884
rect 5180 37156 5236 37166
rect 5404 37156 5460 37166
rect 5180 37154 5348 37156
rect 5180 37102 5182 37154
rect 5234 37102 5348 37154
rect 5180 37100 5348 37102
rect 5180 37090 5236 37100
rect 5292 37042 5348 37100
rect 5292 36990 5294 37042
rect 5346 36990 5348 37042
rect 5292 36978 5348 36990
rect 5068 36876 5236 36932
rect 4956 35298 5012 35308
rect 5068 36260 5124 36270
rect 5068 34916 5124 36204
rect 4844 34738 4900 34748
rect 4956 34860 5124 34916
rect 4284 34402 4340 34412
rect 4508 34692 4564 34702
rect 4060 34130 4116 34142
rect 4060 34078 4062 34130
rect 4114 34078 4116 34130
rect 4060 33572 4116 34078
rect 4172 34020 4228 34300
rect 4508 34354 4564 34636
rect 4508 34302 4510 34354
rect 4562 34302 4564 34354
rect 4508 34290 4564 34302
rect 4172 33954 4228 33964
rect 4284 34130 4340 34142
rect 4284 34078 4286 34130
rect 4338 34078 4340 34130
rect 4284 33908 4340 34078
rect 4284 33842 4340 33852
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4060 33460 4116 33516
rect 4060 33404 4228 33460
rect 3948 33348 4004 33404
rect 3948 33292 4116 33348
rect 3500 31938 3556 31948
rect 3612 32060 3780 32116
rect 3836 32564 3892 32574
rect 3388 31890 3444 31902
rect 3388 31838 3390 31890
rect 3442 31838 3444 31890
rect 2828 31668 2884 31678
rect 2828 31574 2884 31612
rect 3388 31332 3444 31838
rect 3388 31266 3444 31276
rect 2716 31220 2772 31230
rect 2492 31218 2772 31220
rect 2492 31166 2718 31218
rect 2770 31166 2772 31218
rect 2492 31164 2772 31166
rect 2380 30098 2436 30110
rect 2380 30046 2382 30098
rect 2434 30046 2436 30098
rect 2380 29876 2436 30046
rect 2380 29810 2436 29820
rect 2492 29652 2548 31164
rect 2716 31154 2772 31164
rect 3612 30770 3668 32060
rect 3612 30718 3614 30770
rect 3666 30718 3668 30770
rect 3388 30436 3444 30446
rect 2044 28702 2046 28754
rect 2098 28702 2100 28754
rect 2044 28690 2100 28702
rect 2380 29596 2548 29652
rect 2716 30212 2772 30222
rect 2044 27972 2100 27982
rect 1932 27748 1988 27758
rect 1932 27654 1988 27692
rect 1932 26852 1988 26862
rect 1932 26758 1988 26796
rect 1932 26516 1988 26526
rect 1932 26422 1988 26460
rect 1820 24050 1876 25564
rect 2044 25618 2100 27916
rect 2380 26852 2436 29596
rect 2716 29540 2772 30156
rect 2492 29538 2772 29540
rect 2492 29486 2718 29538
rect 2770 29486 2772 29538
rect 2492 29484 2772 29486
rect 2492 27858 2548 29484
rect 2716 29474 2772 29484
rect 3052 30210 3108 30222
rect 3052 30158 3054 30210
rect 3106 30158 3108 30210
rect 2716 29314 2772 29326
rect 2716 29262 2718 29314
rect 2770 29262 2772 29314
rect 2716 28868 2772 29262
rect 3052 28868 3108 30158
rect 3276 30212 3332 30222
rect 3276 30118 3332 30156
rect 3388 29428 3444 30380
rect 3500 29652 3556 29662
rect 3500 29558 3556 29596
rect 3388 29372 3556 29428
rect 2716 28812 3444 28868
rect 3164 28754 3220 28812
rect 3164 28702 3166 28754
rect 3218 28702 3220 28754
rect 3164 28690 3220 28702
rect 2492 27806 2494 27858
rect 2546 27806 2548 27858
rect 2492 26964 2548 27806
rect 3052 28642 3108 28654
rect 3052 28590 3054 28642
rect 3106 28590 3108 28642
rect 3052 27858 3108 28590
rect 3052 27806 3054 27858
rect 3106 27806 3108 27858
rect 2492 26898 2548 26908
rect 2604 27188 2660 27198
rect 2380 26628 2436 26796
rect 2380 26572 2548 26628
rect 2044 25566 2046 25618
rect 2098 25566 2100 25618
rect 2044 25554 2100 25566
rect 2268 26516 2324 26526
rect 2268 26292 2324 26460
rect 2380 26292 2436 26302
rect 2268 26290 2436 26292
rect 2268 26238 2382 26290
rect 2434 26238 2436 26290
rect 2268 26236 2436 26238
rect 2268 25508 2324 26236
rect 2380 26226 2436 26236
rect 2492 26180 2548 26572
rect 2492 26114 2548 26124
rect 2268 24946 2324 25452
rect 2380 25284 2436 25294
rect 2380 25190 2436 25228
rect 2268 24894 2270 24946
rect 2322 24894 2324 24946
rect 1820 23998 1822 24050
rect 1874 23998 1876 24050
rect 1820 23986 1876 23998
rect 1932 24610 1988 24622
rect 1932 24558 1934 24610
rect 1986 24558 1988 24610
rect 1484 23426 1540 23436
rect 1932 22930 1988 24558
rect 1932 22878 1934 22930
rect 1986 22878 1988 22930
rect 1932 22866 1988 22878
rect 2044 24498 2100 24510
rect 2044 24446 2046 24498
rect 2098 24446 2100 24498
rect 2044 23378 2100 24446
rect 2044 23326 2046 23378
rect 2098 23326 2100 23378
rect 1820 22146 1876 22158
rect 1820 22094 1822 22146
rect 1874 22094 1876 22146
rect 1820 22036 1876 22094
rect 1820 21970 1876 21980
rect 2044 21812 2100 23326
rect 2268 23268 2324 24894
rect 2380 24052 2436 24062
rect 2604 24052 2660 27132
rect 3052 27076 3108 27806
rect 3052 26944 3108 27020
rect 3388 27074 3444 28812
rect 3500 27748 3556 29372
rect 3500 27682 3556 27692
rect 3388 27022 3390 27074
rect 3442 27022 3444 27074
rect 2940 26516 2996 26526
rect 2940 26422 2996 26460
rect 3388 26292 3444 27022
rect 3388 26226 3444 26236
rect 3500 27188 3556 27198
rect 2828 26180 2884 26190
rect 2716 25172 2772 25182
rect 2716 24946 2772 25116
rect 2716 24894 2718 24946
rect 2770 24894 2772 24946
rect 2716 24882 2772 24894
rect 2380 24050 2660 24052
rect 2380 23998 2382 24050
rect 2434 23998 2660 24050
rect 2380 23996 2660 23998
rect 2716 24498 2772 24510
rect 2716 24446 2718 24498
rect 2770 24446 2772 24498
rect 2716 24050 2772 24446
rect 2716 23998 2718 24050
rect 2770 23998 2772 24050
rect 2380 23986 2436 23996
rect 2268 23202 2324 23212
rect 2380 23042 2436 23054
rect 2380 22990 2382 23042
rect 2434 22990 2436 23042
rect 2380 22930 2436 22990
rect 2380 22878 2382 22930
rect 2434 22878 2436 22930
rect 2380 22866 2436 22878
rect 2156 22484 2212 22494
rect 2156 22390 2212 22428
rect 2604 22484 2660 22494
rect 2716 22484 2772 23998
rect 2604 22482 2772 22484
rect 2604 22430 2606 22482
rect 2658 22430 2772 22482
rect 2604 22428 2772 22430
rect 2828 23378 2884 26124
rect 3276 26180 3332 26190
rect 3276 26086 3332 26124
rect 3500 26068 3556 27132
rect 3388 26012 3556 26068
rect 2940 25844 2996 25854
rect 2940 25618 2996 25788
rect 2940 25566 2942 25618
rect 2994 25566 2996 25618
rect 2940 25554 2996 25566
rect 3164 25284 3220 25294
rect 3164 24610 3220 25228
rect 3388 25172 3444 26012
rect 3164 24558 3166 24610
rect 3218 24558 3220 24610
rect 3164 24052 3220 24558
rect 3276 25116 3444 25172
rect 3500 25844 3556 25854
rect 3276 24498 3332 25116
rect 3276 24446 3278 24498
rect 3330 24446 3332 24498
rect 3276 24434 3332 24446
rect 3388 24162 3444 24174
rect 3388 24110 3390 24162
rect 3442 24110 3444 24162
rect 3276 24052 3332 24062
rect 3164 24050 3332 24052
rect 3164 23998 3278 24050
rect 3330 23998 3332 24050
rect 3164 23996 3332 23998
rect 3276 23986 3332 23996
rect 2828 23326 2830 23378
rect 2882 23326 2884 23378
rect 2828 22484 2884 23326
rect 3276 23042 3332 23054
rect 3276 22990 3278 23042
rect 3330 22990 3332 23042
rect 2604 22418 2660 22428
rect 2828 22418 2884 22428
rect 2940 22930 2996 22942
rect 2940 22878 2942 22930
rect 2994 22878 2996 22930
rect 2716 21924 2772 21934
rect 2156 21812 2212 21822
rect 2044 21810 2212 21812
rect 2044 21758 2158 21810
rect 2210 21758 2212 21810
rect 2044 21756 2212 21758
rect 1820 21700 1876 21710
rect 1820 21606 1876 21644
rect 2156 21588 2212 21756
rect 2156 21522 2212 21532
rect 2268 21812 2324 21822
rect 2716 21812 2772 21868
rect 2268 20914 2324 21756
rect 2268 20862 2270 20914
rect 2322 20862 2324 20914
rect 2268 20850 2324 20862
rect 2604 21810 2772 21812
rect 2604 21758 2718 21810
rect 2770 21758 2772 21810
rect 2604 21756 2772 21758
rect 1932 20578 1988 20590
rect 1932 20526 1934 20578
rect 1986 20526 1988 20578
rect 1932 20356 1988 20526
rect 1932 20290 1988 20300
rect 2604 20244 2660 21756
rect 2716 21746 2772 21756
rect 2940 21588 2996 22878
rect 3276 22930 3332 22990
rect 3276 22878 3278 22930
rect 3330 22878 3332 22930
rect 3276 22866 3332 22878
rect 3052 22146 3108 22158
rect 3052 22094 3054 22146
rect 3106 22094 3108 22146
rect 3052 21812 3108 22094
rect 3388 21812 3444 24110
rect 3500 24164 3556 25788
rect 3612 25284 3668 30718
rect 3724 31892 3780 31902
rect 3724 30994 3780 31836
rect 3724 30942 3726 30994
rect 3778 30942 3780 30994
rect 3724 28868 3780 30942
rect 3836 31554 3892 32508
rect 3836 31502 3838 31554
rect 3890 31502 3892 31554
rect 3836 30884 3892 31502
rect 3836 30818 3892 30828
rect 4060 32450 4116 33292
rect 4060 32398 4062 32450
rect 4114 32398 4116 32450
rect 3724 28802 3780 28812
rect 3948 29092 4004 29102
rect 3948 28866 4004 29036
rect 3948 28814 3950 28866
rect 4002 28814 4004 28866
rect 3948 28802 4004 28814
rect 3836 27748 3892 27758
rect 3724 26516 3780 26526
rect 3836 26516 3892 27692
rect 4060 26908 4116 32398
rect 4172 31332 4228 33404
rect 4284 33236 4340 33246
rect 4284 33142 4340 33180
rect 4844 33236 4900 33246
rect 4956 33236 5012 34860
rect 5068 34690 5124 34702
rect 5068 34638 5070 34690
rect 5122 34638 5124 34690
rect 5068 33684 5124 34638
rect 5180 34244 5236 36876
rect 5404 36036 5460 37100
rect 5292 35980 5460 36036
rect 5516 37044 5572 38668
rect 5628 38592 5684 38668
rect 5740 38388 5796 38398
rect 5740 38050 5796 38332
rect 5740 37998 5742 38050
rect 5794 37998 5796 38050
rect 5740 37986 5796 37998
rect 5628 37156 5684 37166
rect 5628 37062 5684 37100
rect 5292 34580 5348 35980
rect 5516 35810 5572 36988
rect 5740 36820 5796 36830
rect 5740 35924 5796 36764
rect 5852 36148 5908 40012
rect 6188 39844 6244 43596
rect 6300 43428 6356 43438
rect 6300 42196 6356 43372
rect 6636 42978 6692 44604
rect 6860 44548 6916 44558
rect 6972 44548 7028 45052
rect 7196 45042 7252 45052
rect 7084 44884 7140 44894
rect 7420 44884 7476 46172
rect 7532 46004 7588 46014
rect 7532 45890 7588 45948
rect 7532 45838 7534 45890
rect 7586 45838 7588 45890
rect 7532 45332 7588 45838
rect 7532 45266 7588 45276
rect 7756 45666 7812 45678
rect 7756 45614 7758 45666
rect 7810 45614 7812 45666
rect 7644 45108 7700 45118
rect 7756 45108 7812 45614
rect 7644 45106 7812 45108
rect 7644 45054 7646 45106
rect 7698 45054 7812 45106
rect 7644 45052 7812 45054
rect 7868 45108 7924 46620
rect 8092 46562 8148 46574
rect 8092 46510 8094 46562
rect 8146 46510 8148 46562
rect 7980 45892 8036 45902
rect 7980 45798 8036 45836
rect 8092 45668 8148 46510
rect 8204 46564 8260 49084
rect 8540 49074 8596 49084
rect 8204 46498 8260 46508
rect 8316 48916 8372 48926
rect 8204 45780 8260 45790
rect 8204 45686 8260 45724
rect 8092 45602 8148 45612
rect 8092 45108 8148 45118
rect 7868 45106 8148 45108
rect 7868 45054 8094 45106
rect 8146 45054 8148 45106
rect 7868 45052 8148 45054
rect 7644 45042 7700 45052
rect 7084 44882 7476 44884
rect 7084 44830 7086 44882
rect 7138 44830 7476 44882
rect 7084 44828 7476 44830
rect 7084 44660 7140 44828
rect 7084 44594 7140 44604
rect 6860 44546 7028 44548
rect 6860 44494 6862 44546
rect 6914 44494 7028 44546
rect 6860 44492 7028 44494
rect 6860 44482 6916 44492
rect 7196 44100 7252 44110
rect 7084 43652 7140 43662
rect 6748 43540 6804 43550
rect 6748 43446 6804 43484
rect 6636 42926 6638 42978
rect 6690 42926 6692 42978
rect 6412 42868 6468 42878
rect 6412 42754 6468 42812
rect 6412 42702 6414 42754
rect 6466 42702 6468 42754
rect 6412 42690 6468 42702
rect 6524 42530 6580 42542
rect 6524 42478 6526 42530
rect 6578 42478 6580 42530
rect 6524 42308 6580 42478
rect 6636 42532 6692 42926
rect 6860 42868 6916 42878
rect 6860 42754 6916 42812
rect 6860 42702 6862 42754
rect 6914 42702 6916 42754
rect 6860 42690 6916 42702
rect 6636 42466 6692 42476
rect 6524 42242 6580 42252
rect 6300 42130 6356 42140
rect 6636 42082 6692 42094
rect 6636 42030 6638 42082
rect 6690 42030 6692 42082
rect 6524 41970 6580 41982
rect 6524 41918 6526 41970
rect 6578 41918 6580 41970
rect 6524 41860 6580 41918
rect 6636 41972 6692 42030
rect 6636 41906 6692 41916
rect 6524 41794 6580 41804
rect 6972 41858 7028 41870
rect 6972 41806 6974 41858
rect 7026 41806 7028 41858
rect 6972 41410 7028 41806
rect 6972 41358 6974 41410
rect 7026 41358 7028 41410
rect 6972 41346 7028 41358
rect 7084 41298 7140 43596
rect 7196 43426 7252 44044
rect 7420 44098 7476 44110
rect 7420 44046 7422 44098
rect 7474 44046 7476 44098
rect 7420 43540 7476 44046
rect 7868 44098 7924 44110
rect 7868 44046 7870 44098
rect 7922 44046 7924 44098
rect 7868 43876 7924 44046
rect 7868 43810 7924 43820
rect 7868 43652 7924 43662
rect 7644 43540 7700 43550
rect 7476 43484 7588 43540
rect 7420 43474 7476 43484
rect 7196 43374 7198 43426
rect 7250 43374 7252 43426
rect 7196 43314 7252 43374
rect 7196 43262 7198 43314
rect 7250 43262 7252 43314
rect 7196 43250 7252 43262
rect 7420 41972 7476 41982
rect 7420 41878 7476 41916
rect 7084 41246 7086 41298
rect 7138 41246 7140 41298
rect 7084 41234 7140 41246
rect 7196 41858 7252 41870
rect 7196 41806 7198 41858
rect 7250 41806 7252 41858
rect 6748 40852 6804 40862
rect 6412 40628 6468 40638
rect 6412 40534 6468 40572
rect 6748 40292 6804 40796
rect 6972 40628 7028 40638
rect 6972 40534 7028 40572
rect 7196 40628 7252 41806
rect 7420 41188 7476 41198
rect 7420 41074 7476 41132
rect 7420 41022 7422 41074
rect 7474 41022 7476 41074
rect 7420 41010 7476 41022
rect 7532 40964 7588 43484
rect 7644 43446 7700 43484
rect 7756 42868 7812 42878
rect 7756 42644 7812 42812
rect 7532 40898 7588 40908
rect 7644 42642 7812 42644
rect 7644 42590 7758 42642
rect 7810 42590 7812 42642
rect 7644 42588 7812 42590
rect 7196 40562 7252 40572
rect 7644 40404 7700 42588
rect 7756 42578 7812 42588
rect 7868 42642 7924 43596
rect 7868 42590 7870 42642
rect 7922 42590 7924 42642
rect 7196 40348 7700 40404
rect 7756 40852 7812 40862
rect 7756 40402 7812 40796
rect 7868 40516 7924 42590
rect 7868 40450 7924 40460
rect 7980 40628 8036 45052
rect 8092 45042 8148 45052
rect 8204 43764 8260 43774
rect 8316 43764 8372 48860
rect 8428 48802 8484 48814
rect 8428 48750 8430 48802
rect 8482 48750 8484 48802
rect 8428 48692 8484 48750
rect 8764 48692 8820 50430
rect 9772 50484 9828 51100
rect 9884 50596 9940 50606
rect 9996 50596 10052 52220
rect 10332 52612 10388 52622
rect 9884 50594 10052 50596
rect 9884 50542 9886 50594
rect 9938 50542 10052 50594
rect 9884 50540 10052 50542
rect 9884 50530 9940 50540
rect 9772 50418 9828 50428
rect 8988 50372 9044 50382
rect 8988 49698 9044 50316
rect 9996 49924 10052 50540
rect 10220 50708 10276 50718
rect 10220 50034 10276 50652
rect 10220 49982 10222 50034
rect 10274 49982 10276 50034
rect 10220 49970 10276 49982
rect 10332 50036 10388 52556
rect 10444 52052 10500 54012
rect 11116 54068 11172 54350
rect 11116 54002 11172 54012
rect 10892 53508 10948 53518
rect 10892 53506 11060 53508
rect 10892 53454 10894 53506
rect 10946 53454 11060 53506
rect 10892 53452 11060 53454
rect 10892 53442 10948 53452
rect 10892 52834 10948 52846
rect 10892 52782 10894 52834
rect 10946 52782 10948 52834
rect 10892 52612 10948 52782
rect 10892 52546 10948 52556
rect 10556 52164 10612 52174
rect 11004 52164 11060 53452
rect 11228 52612 11284 55020
rect 11340 55010 11396 55020
rect 11452 54738 11508 55804
rect 11452 54686 11454 54738
rect 11506 54686 11508 54738
rect 11452 54674 11508 54686
rect 11676 55522 11732 55534
rect 11676 55470 11678 55522
rect 11730 55470 11732 55522
rect 11340 53506 11396 53518
rect 11340 53454 11342 53506
rect 11394 53454 11396 53506
rect 11340 53396 11396 53454
rect 11340 53340 11620 53396
rect 11228 52546 11284 52556
rect 11340 52834 11396 52846
rect 11340 52782 11342 52834
rect 11394 52782 11396 52834
rect 11340 52276 11396 52782
rect 11340 52210 11396 52220
rect 11116 52164 11172 52174
rect 10556 52162 10836 52164
rect 10556 52110 10558 52162
rect 10610 52110 10836 52162
rect 10556 52108 10836 52110
rect 11004 52162 11172 52164
rect 11004 52110 11118 52162
rect 11170 52110 11172 52162
rect 11004 52108 11172 52110
rect 10556 52098 10612 52108
rect 10444 51958 10500 51996
rect 10444 51378 10500 51390
rect 10444 51326 10446 51378
rect 10498 51326 10500 51378
rect 10444 51268 10500 51326
rect 10444 51202 10500 51212
rect 10668 51378 10724 51390
rect 10668 51326 10670 51378
rect 10722 51326 10724 51378
rect 10556 50372 10612 50382
rect 10332 49980 10500 50036
rect 8988 49646 8990 49698
rect 9042 49646 9044 49698
rect 8876 48804 8932 48814
rect 8876 48710 8932 48748
rect 8428 48626 8484 48636
rect 8540 48636 8820 48692
rect 8428 48244 8484 48254
rect 8428 48150 8484 48188
rect 8428 44436 8484 44446
rect 8428 44322 8484 44380
rect 8428 44270 8430 44322
rect 8482 44270 8484 44322
rect 8428 44258 8484 44270
rect 8540 44100 8596 48636
rect 8764 48466 8820 48478
rect 8764 48414 8766 48466
rect 8818 48414 8820 48466
rect 8652 48244 8708 48254
rect 8652 47570 8708 48188
rect 8764 47908 8820 48414
rect 8988 48468 9044 49646
rect 9548 49812 9604 49822
rect 9212 49476 9268 49486
rect 9212 49138 9268 49420
rect 9212 49086 9214 49138
rect 9266 49086 9268 49138
rect 9212 49074 9268 49086
rect 8988 48402 9044 48412
rect 8764 47842 8820 47852
rect 9324 47684 9380 47694
rect 8652 47518 8654 47570
rect 8706 47518 8708 47570
rect 8652 46004 8708 47518
rect 8988 47682 9380 47684
rect 8988 47630 9326 47682
rect 9378 47630 9380 47682
rect 8988 47628 9380 47630
rect 8764 47012 8820 47022
rect 8764 46898 8820 46956
rect 8764 46846 8766 46898
rect 8818 46846 8820 46898
rect 8764 46834 8820 46846
rect 8988 46786 9044 47628
rect 9324 47618 9380 47628
rect 9436 47572 9492 47582
rect 9436 47458 9492 47516
rect 9436 47406 9438 47458
rect 9490 47406 9492 47458
rect 9436 47394 9492 47406
rect 9212 47348 9268 47358
rect 9212 47254 9268 47292
rect 9548 47068 9604 49756
rect 9884 49026 9940 49038
rect 9884 48974 9886 49026
rect 9938 48974 9940 49026
rect 9884 48804 9940 48974
rect 9996 49026 10052 49868
rect 10108 49810 10164 49822
rect 10332 49812 10388 49822
rect 10108 49758 10110 49810
rect 10162 49758 10164 49810
rect 10108 49364 10164 49758
rect 10108 49298 10164 49308
rect 10220 49810 10388 49812
rect 10220 49758 10334 49810
rect 10386 49758 10388 49810
rect 10220 49756 10388 49758
rect 10444 49812 10500 49980
rect 10556 50034 10612 50316
rect 10556 49982 10558 50034
rect 10610 49982 10612 50034
rect 10556 49970 10612 49982
rect 10668 50036 10724 51326
rect 10780 50428 10836 52108
rect 10892 52052 10948 52062
rect 10892 52050 11060 52052
rect 10892 51998 10894 52050
rect 10946 51998 11060 52050
rect 10892 51996 11060 51998
rect 10892 51986 10948 51996
rect 11004 51604 11060 51996
rect 11116 51940 11172 52108
rect 11116 51874 11172 51884
rect 11564 51828 11620 53340
rect 11676 52388 11732 55470
rect 11788 54516 11844 54526
rect 11788 53170 11844 54460
rect 11900 53842 11956 55916
rect 12460 55860 12516 59612
rect 12796 59556 12852 59566
rect 12796 59442 12852 59500
rect 12796 59390 12798 59442
rect 12850 59390 12852 59442
rect 12796 59378 12852 59390
rect 12908 58884 12964 59726
rect 13580 59778 13636 59790
rect 13580 59726 13582 59778
rect 13634 59726 13636 59778
rect 13468 59668 13524 59678
rect 13580 59668 13636 59726
rect 13524 59612 13636 59668
rect 14028 59778 14084 59790
rect 14028 59726 14030 59778
rect 14082 59726 14084 59778
rect 12908 58818 12964 58828
rect 13020 59220 13076 59230
rect 12684 58436 12740 58446
rect 12684 58324 12740 58380
rect 13020 58434 13076 59164
rect 13244 59108 13300 59118
rect 13244 59014 13300 59052
rect 13020 58382 13022 58434
rect 13074 58382 13076 58434
rect 13020 58370 13076 58382
rect 13468 58996 13524 59612
rect 12236 55804 12516 55860
rect 12572 58322 12740 58324
rect 12572 58270 12686 58322
rect 12738 58270 12740 58322
rect 12572 58268 12740 58270
rect 12124 55412 12180 55450
rect 12124 55346 12180 55356
rect 12012 55300 12068 55310
rect 12012 54738 12068 55244
rect 12012 54686 12014 54738
rect 12066 54686 12068 54738
rect 12012 54674 12068 54686
rect 12124 55188 12180 55198
rect 12124 54516 12180 55132
rect 11900 53790 11902 53842
rect 11954 53790 11956 53842
rect 11900 53778 11956 53790
rect 12012 54460 12180 54516
rect 11788 53118 11790 53170
rect 11842 53118 11844 53170
rect 11788 52722 11844 53118
rect 11788 52670 11790 52722
rect 11842 52670 11844 52722
rect 11788 52658 11844 52670
rect 11900 53172 11956 53182
rect 11676 52322 11732 52332
rect 11564 51762 11620 51772
rect 11676 52162 11732 52174
rect 11676 52110 11678 52162
rect 11730 52110 11732 52162
rect 11004 51548 11396 51604
rect 10892 51380 10948 51390
rect 11116 51380 11172 51390
rect 10892 51378 11060 51380
rect 10892 51326 10894 51378
rect 10946 51326 11060 51378
rect 10892 51324 11060 51326
rect 10892 51314 10948 51324
rect 10892 50596 10948 50634
rect 10892 50530 10948 50540
rect 10780 50372 10948 50428
rect 10668 49970 10724 49980
rect 10892 50036 10948 50372
rect 11004 50370 11060 51324
rect 11116 51286 11172 51324
rect 11340 51378 11396 51548
rect 11340 51326 11342 51378
rect 11394 51326 11396 51378
rect 11340 51314 11396 51326
rect 11564 51156 11620 51166
rect 11564 51062 11620 51100
rect 11676 50708 11732 52110
rect 11676 50642 11732 50652
rect 11004 50318 11006 50370
rect 11058 50318 11060 50370
rect 11004 50306 11060 50318
rect 11340 50370 11396 50382
rect 11340 50318 11342 50370
rect 11394 50318 11396 50370
rect 10892 49970 10948 49980
rect 10444 49756 10836 49812
rect 9996 48974 9998 49026
rect 10050 48974 10052 49026
rect 9996 48962 10052 48974
rect 9884 48738 9940 48748
rect 10108 48802 10164 48814
rect 10108 48750 10110 48802
rect 10162 48750 10164 48802
rect 9772 48468 9828 48478
rect 9660 48466 9828 48468
rect 9660 48414 9774 48466
rect 9826 48414 9828 48466
rect 9660 48412 9828 48414
rect 9660 47684 9716 48412
rect 9772 48402 9828 48412
rect 9996 48468 10052 48478
rect 9772 48242 9828 48254
rect 9772 48190 9774 48242
rect 9826 48190 9828 48242
rect 9772 48020 9828 48190
rect 9996 48020 10052 48412
rect 10108 48242 10164 48750
rect 10220 48692 10276 49756
rect 10332 49746 10388 49756
rect 10332 49028 10388 49038
rect 10332 48934 10388 48972
rect 10668 49028 10724 49038
rect 10220 48468 10276 48636
rect 10220 48402 10276 48412
rect 10332 48804 10388 48814
rect 10108 48190 10110 48242
rect 10162 48190 10164 48242
rect 10108 48178 10164 48190
rect 10220 48244 10276 48254
rect 9996 47964 10164 48020
rect 9772 47954 9828 47964
rect 9772 47684 9828 47694
rect 9660 47682 9828 47684
rect 9660 47630 9774 47682
rect 9826 47630 9828 47682
rect 9660 47628 9828 47630
rect 9772 47618 9828 47628
rect 9996 47458 10052 47470
rect 9996 47406 9998 47458
rect 10050 47406 10052 47458
rect 9548 47012 9716 47068
rect 8988 46734 8990 46786
rect 9042 46734 9044 46786
rect 8988 46722 9044 46734
rect 9100 46676 9156 46686
rect 8652 45938 8708 45948
rect 8764 46564 8820 46574
rect 8764 45890 8820 46508
rect 8876 46562 8932 46574
rect 8876 46510 8878 46562
rect 8930 46510 8932 46562
rect 8876 46452 8932 46510
rect 8876 46386 8932 46396
rect 8764 45838 8766 45890
rect 8818 45838 8820 45890
rect 8652 44994 8708 45006
rect 8652 44942 8654 44994
rect 8706 44942 8708 44994
rect 8652 44436 8708 44942
rect 8652 44370 8708 44380
rect 8540 44034 8596 44044
rect 8204 43762 8372 43764
rect 8204 43710 8206 43762
rect 8258 43710 8372 43762
rect 8204 43708 8372 43710
rect 8540 43876 8596 43886
rect 8204 43698 8260 43708
rect 8540 43428 8596 43820
rect 8764 43652 8820 45838
rect 8876 46004 8932 46014
rect 8876 45668 8932 45948
rect 9100 45892 9156 46620
rect 9100 45760 9156 45836
rect 8876 45666 9044 45668
rect 8876 45614 8878 45666
rect 8930 45614 9044 45666
rect 8876 45612 9044 45614
rect 8876 45602 8932 45612
rect 8988 44210 9044 45612
rect 9660 44996 9716 47012
rect 9772 46564 9828 46574
rect 9772 46470 9828 46508
rect 9772 46228 9828 46238
rect 9772 46002 9828 46172
rect 9772 45950 9774 46002
rect 9826 45950 9828 46002
rect 9772 45938 9828 45950
rect 9660 44902 9716 44940
rect 8988 44158 8990 44210
rect 9042 44158 9044 44210
rect 8988 43988 9044 44158
rect 9212 44884 9268 44894
rect 9212 44210 9268 44828
rect 9212 44158 9214 44210
rect 9266 44158 9268 44210
rect 9212 44146 9268 44158
rect 9436 44212 9492 44222
rect 8988 43932 9380 43988
rect 8764 43586 8820 43596
rect 8876 43876 8932 43886
rect 8540 43426 8708 43428
rect 8540 43374 8542 43426
rect 8594 43374 8708 43426
rect 8540 43372 8708 43374
rect 8540 43362 8596 43372
rect 8092 43092 8148 43102
rect 8092 42754 8148 43036
rect 8092 42702 8094 42754
rect 8146 42702 8148 42754
rect 8092 42690 8148 42702
rect 8428 42868 8484 42878
rect 8428 42532 8484 42812
rect 8540 42756 8596 42766
rect 8540 42662 8596 42700
rect 8428 42476 8596 42532
rect 8428 42308 8484 42318
rect 8204 42084 8260 42094
rect 7756 40350 7758 40402
rect 7810 40350 7812 40402
rect 7196 40292 7252 40348
rect 7756 40338 7812 40350
rect 6636 40236 6804 40292
rect 7084 40236 7252 40292
rect 6188 39788 6468 39844
rect 6300 39620 6356 39630
rect 6188 39506 6244 39518
rect 6188 39454 6190 39506
rect 6242 39454 6244 39506
rect 6188 39396 6244 39454
rect 6076 38836 6132 38846
rect 6076 38742 6132 38780
rect 5964 37268 6020 37278
rect 5964 36932 6020 37212
rect 6076 37156 6132 37166
rect 6188 37156 6244 39340
rect 6300 39506 6356 39564
rect 6300 39454 6302 39506
rect 6354 39454 6356 39506
rect 6300 38948 6356 39454
rect 6300 38882 6356 38892
rect 6412 38834 6468 39788
rect 6636 39620 6692 40236
rect 6636 39554 6692 39564
rect 7084 40178 7140 40236
rect 7308 40180 7364 40190
rect 7868 40180 7924 40190
rect 7084 40126 7086 40178
rect 7138 40126 7140 40178
rect 7084 39844 7140 40126
rect 6524 39396 6580 39406
rect 6524 39394 6692 39396
rect 6524 39342 6526 39394
rect 6578 39342 6692 39394
rect 6524 39340 6692 39342
rect 6524 39330 6580 39340
rect 6412 38782 6414 38834
rect 6466 38782 6468 38834
rect 6412 38770 6468 38782
rect 6300 38724 6356 38762
rect 6300 38658 6356 38668
rect 6636 37940 6692 39340
rect 6860 39172 6916 39182
rect 6748 38834 6804 38846
rect 6748 38782 6750 38834
rect 6802 38782 6804 38834
rect 6748 38388 6804 38782
rect 6748 38322 6804 38332
rect 6636 37874 6692 37884
rect 6748 38052 6804 38062
rect 6748 37492 6804 37996
rect 6860 37938 6916 39116
rect 7084 38724 7140 39788
rect 7084 38658 7140 38668
rect 7196 40124 7308 40180
rect 7196 38668 7252 40124
rect 7308 40086 7364 40124
rect 7420 40178 7924 40180
rect 7420 40126 7870 40178
rect 7922 40126 7924 40178
rect 7420 40124 7924 40126
rect 7420 39506 7476 40124
rect 7868 40114 7924 40124
rect 7420 39454 7422 39506
rect 7474 39454 7476 39506
rect 7308 38948 7364 38958
rect 7308 38854 7364 38892
rect 7196 38612 7364 38668
rect 6860 37886 6862 37938
rect 6914 37886 6916 37938
rect 6860 37874 6916 37886
rect 7084 38052 7140 38062
rect 6748 37426 6804 37436
rect 6860 37268 6916 37278
rect 6188 37100 6356 37156
rect 6076 37062 6132 37100
rect 5964 36876 6132 36932
rect 5852 36082 5908 36092
rect 5964 36482 6020 36494
rect 5964 36430 5966 36482
rect 6018 36430 6020 36482
rect 5740 35868 5908 35924
rect 5516 35758 5518 35810
rect 5570 35758 5572 35810
rect 5404 35698 5460 35710
rect 5404 35646 5406 35698
rect 5458 35646 5460 35698
rect 5404 35028 5460 35646
rect 5516 35588 5572 35758
rect 5740 35700 5796 35710
rect 5740 35606 5796 35644
rect 5516 35522 5572 35532
rect 5404 34962 5460 34972
rect 5516 35364 5572 35374
rect 5516 34916 5572 35308
rect 5516 34850 5572 34860
rect 5292 34514 5348 34524
rect 5516 34580 5572 34590
rect 5404 34468 5460 34478
rect 5404 34354 5460 34412
rect 5404 34302 5406 34354
rect 5458 34302 5460 34354
rect 5404 34290 5460 34302
rect 5180 34178 5236 34188
rect 5292 34242 5348 34254
rect 5292 34190 5294 34242
rect 5346 34190 5348 34242
rect 5292 33908 5348 34190
rect 5516 34132 5572 34524
rect 5292 33842 5348 33852
rect 5404 34076 5572 34132
rect 5068 33618 5124 33628
rect 4900 33180 5012 33236
rect 5180 33348 5236 33358
rect 4284 32674 4340 32686
rect 4284 32622 4286 32674
rect 4338 32622 4340 32674
rect 4284 32564 4340 32622
rect 4284 32498 4340 32508
rect 4508 32564 4564 32574
rect 4508 32470 4564 32508
rect 4172 31266 4228 31276
rect 4284 32340 4340 32350
rect 4172 30996 4228 31006
rect 4172 29428 4228 30940
rect 4284 30436 4340 32284
rect 4844 32228 4900 33180
rect 5068 32564 5124 32574
rect 5180 32564 5236 33292
rect 5068 32562 5236 32564
rect 5068 32510 5070 32562
rect 5122 32510 5236 32562
rect 5068 32508 5236 32510
rect 5068 32498 5124 32508
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4844 32162 4900 32172
rect 4476 32106 4740 32116
rect 5068 31892 5124 31902
rect 5068 31798 5124 31836
rect 4620 31554 4676 31566
rect 4620 31502 4622 31554
rect 4674 31502 4676 31554
rect 4620 30772 4676 31502
rect 4844 30994 4900 31006
rect 4844 30942 4846 30994
rect 4898 30942 4900 30994
rect 4844 30884 4900 30942
rect 5180 30996 5236 32508
rect 5180 30902 5236 30940
rect 5292 33124 5348 33134
rect 4844 30818 4900 30828
rect 4620 30706 4676 30716
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4284 30380 4676 30436
rect 4620 30210 4676 30380
rect 5068 30324 5124 30334
rect 5068 30212 5124 30268
rect 4620 30158 4622 30210
rect 4674 30158 4676 30210
rect 4620 30146 4676 30158
rect 4956 30156 5124 30212
rect 4956 30154 5012 30156
rect 4956 30102 4958 30154
rect 5010 30102 5012 30154
rect 4956 30090 5012 30102
rect 4844 29988 4900 29998
rect 5292 29988 5348 33068
rect 5404 32788 5460 34076
rect 5516 33908 5572 33918
rect 5740 33908 5796 33918
rect 5516 33906 5796 33908
rect 5516 33854 5518 33906
rect 5570 33854 5742 33906
rect 5794 33854 5796 33906
rect 5516 33852 5796 33854
rect 5516 33012 5572 33852
rect 5740 33842 5796 33852
rect 5852 33684 5908 35868
rect 5964 35364 6020 36430
rect 6076 35924 6132 36876
rect 6188 36708 6244 36718
rect 6188 36594 6244 36652
rect 6188 36542 6190 36594
rect 6242 36542 6244 36594
rect 6188 36530 6244 36542
rect 6076 35868 6244 35924
rect 5964 35298 6020 35308
rect 6076 34804 6132 34814
rect 5964 34692 6020 34702
rect 5964 34598 6020 34636
rect 6076 34690 6132 34748
rect 6076 34638 6078 34690
rect 6130 34638 6132 34690
rect 5964 34244 6020 34254
rect 5964 34150 6020 34188
rect 6076 33796 6132 34638
rect 6188 34802 6244 35868
rect 6300 35586 6356 37100
rect 6524 37154 6580 37166
rect 6524 37102 6526 37154
rect 6578 37102 6580 37154
rect 6412 37042 6468 37054
rect 6412 36990 6414 37042
rect 6466 36990 6468 37042
rect 6412 36596 6468 36990
rect 6524 36820 6580 37102
rect 6524 36754 6580 36764
rect 6636 37156 6692 37166
rect 6412 36540 6580 36596
rect 6524 36482 6580 36540
rect 6524 36430 6526 36482
rect 6578 36430 6580 36482
rect 6412 36370 6468 36382
rect 6412 36318 6414 36370
rect 6466 36318 6468 36370
rect 6412 36260 6468 36318
rect 6412 36194 6468 36204
rect 6300 35534 6302 35586
rect 6354 35534 6356 35586
rect 6300 35522 6356 35534
rect 6524 35308 6580 36430
rect 6412 35252 6580 35308
rect 6188 34750 6190 34802
rect 6242 34750 6244 34802
rect 6188 33906 6244 34750
rect 6188 33854 6190 33906
rect 6242 33854 6244 33906
rect 6188 33842 6244 33854
rect 6300 34916 6356 34926
rect 5740 33628 5908 33684
rect 5964 33740 6132 33796
rect 5628 33348 5684 33358
rect 5628 33254 5684 33292
rect 5516 32956 5684 33012
rect 5516 32788 5572 32798
rect 5404 32732 5516 32788
rect 5516 32694 5572 32732
rect 5516 32228 5572 32238
rect 4844 29986 5348 29988
rect 4844 29934 4846 29986
rect 4898 29934 5348 29986
rect 4844 29932 5348 29934
rect 4844 29922 4900 29932
rect 4620 29876 4676 29886
rect 4284 29652 4340 29662
rect 4284 29558 4340 29596
rect 4620 29540 4676 29820
rect 4172 29372 4340 29428
rect 4172 28868 4228 28878
rect 4172 27970 4228 28812
rect 4172 27918 4174 27970
rect 4226 27918 4228 27970
rect 4172 27906 4228 27918
rect 4172 27636 4228 27646
rect 4172 27188 4228 27580
rect 4172 27056 4228 27132
rect 4060 26852 4228 26908
rect 3724 26514 3892 26516
rect 3724 26462 3726 26514
rect 3778 26462 3892 26514
rect 3724 26460 3892 26462
rect 3724 26450 3780 26460
rect 3612 25218 3668 25228
rect 3724 24948 3780 24958
rect 3724 24854 3780 24892
rect 3836 24948 3892 26460
rect 4060 26628 4116 26638
rect 4060 26292 4116 26572
rect 4172 26516 4228 26852
rect 4284 26628 4340 29372
rect 4620 29426 4676 29484
rect 4620 29374 4622 29426
rect 4674 29374 4676 29426
rect 4620 29362 4676 29374
rect 4844 29540 4900 29550
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4508 28756 4564 28766
rect 4508 28662 4564 28700
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4284 26562 4340 26572
rect 4732 26964 4788 26974
rect 4172 26450 4228 26460
rect 4172 26292 4228 26302
rect 4060 26290 4228 26292
rect 4060 26238 4174 26290
rect 4226 26238 4228 26290
rect 4060 26236 4228 26238
rect 4060 25844 4116 26236
rect 4172 26226 4228 26236
rect 4284 26292 4340 26302
rect 4060 25778 4116 25788
rect 4060 25620 4116 25630
rect 4284 25620 4340 26236
rect 4732 26068 4788 26908
rect 4844 26740 4900 29484
rect 5292 29538 5348 29932
rect 5292 29486 5294 29538
rect 5346 29486 5348 29538
rect 5292 29474 5348 29486
rect 5404 30996 5460 31006
rect 5404 30324 5460 30940
rect 5404 29426 5460 30268
rect 5516 29652 5572 32172
rect 5628 30436 5684 32956
rect 5740 31892 5796 33628
rect 5852 31892 5908 31902
rect 5740 31890 5908 31892
rect 5740 31838 5854 31890
rect 5906 31838 5908 31890
rect 5740 31836 5908 31838
rect 5628 30370 5684 30380
rect 5516 29586 5572 29596
rect 5404 29374 5406 29426
rect 5458 29374 5460 29426
rect 5180 28756 5236 28766
rect 4956 28642 5012 28654
rect 4956 28590 4958 28642
rect 5010 28590 5012 28642
rect 4956 27188 5012 28590
rect 4956 27122 5012 27132
rect 4956 26964 5012 27002
rect 4956 26898 5012 26908
rect 4844 26674 4900 26684
rect 5068 26852 5124 26862
rect 4844 26404 4900 26414
rect 4844 26310 4900 26348
rect 4956 26180 5012 26190
rect 4732 26012 4900 26068
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4060 25618 4340 25620
rect 4060 25566 4062 25618
rect 4114 25566 4340 25618
rect 4060 25564 4340 25566
rect 4060 25554 4116 25564
rect 4060 25396 4116 25406
rect 4060 25302 4116 25340
rect 3836 24892 4116 24948
rect 3500 22594 3556 24108
rect 3724 24052 3780 24062
rect 3724 23958 3780 23996
rect 3500 22542 3502 22594
rect 3554 22542 3556 22594
rect 3500 22482 3556 22542
rect 3500 22430 3502 22482
rect 3554 22430 3556 22482
rect 3500 22418 3556 22430
rect 3612 23604 3668 23614
rect 3500 21812 3556 21822
rect 3388 21810 3556 21812
rect 3388 21758 3502 21810
rect 3554 21758 3556 21810
rect 3388 21756 3556 21758
rect 3052 21746 3108 21756
rect 2716 21532 2996 21588
rect 3052 21588 3108 21598
rect 2716 20916 2772 21532
rect 3052 21494 3108 21532
rect 2716 20784 2772 20860
rect 3164 21476 3220 21486
rect 3164 20914 3220 21420
rect 3500 21362 3556 21756
rect 3500 21310 3502 21362
rect 3554 21310 3556 21362
rect 3500 21298 3556 21310
rect 3164 20862 3166 20914
rect 3218 20862 3220 20914
rect 3164 20850 3220 20862
rect 3612 20578 3668 23548
rect 3836 23378 3892 24892
rect 3836 23326 3838 23378
rect 3890 23326 3892 23378
rect 3836 23314 3892 23326
rect 3948 24724 4004 24734
rect 3724 22594 3780 22606
rect 3724 22542 3726 22594
rect 3778 22542 3780 22594
rect 3724 21476 3780 22542
rect 3948 21700 4004 24668
rect 4060 24050 4116 24892
rect 4060 23998 4062 24050
rect 4114 23998 4116 24050
rect 4060 23986 4116 23998
rect 4172 23042 4228 23054
rect 4172 22990 4174 23042
rect 4226 22990 4228 23042
rect 4060 22484 4116 22494
rect 4060 22390 4116 22428
rect 3724 21410 3780 21420
rect 3836 21644 3948 21700
rect 3612 20526 3614 20578
rect 3666 20526 3668 20578
rect 2716 20244 2772 20254
rect 2604 20242 2772 20244
rect 2604 20190 2718 20242
rect 2770 20190 2772 20242
rect 2604 20188 2772 20190
rect 2380 20132 2436 20142
rect 1820 19908 1876 19918
rect 1820 19814 1876 19852
rect 2268 19906 2324 19918
rect 2268 19854 2270 19906
rect 2322 19854 2324 19906
rect 1148 19730 1204 19740
rect 2268 17780 2324 19854
rect 2380 19346 2436 20076
rect 2380 19294 2382 19346
rect 2434 19294 2436 19346
rect 2380 19282 2436 19294
rect 2716 19012 2772 20188
rect 3052 20020 3108 20030
rect 3052 19926 3108 19964
rect 3500 20020 3556 20030
rect 3500 19926 3556 19964
rect 3612 19908 3668 20526
rect 3836 19908 3892 21644
rect 3948 21634 4004 21644
rect 4060 22260 4116 22270
rect 3948 21476 4004 21486
rect 3948 21382 4004 21420
rect 4060 21140 4116 22204
rect 4172 22148 4228 22990
rect 4172 22082 4228 22092
rect 3948 21084 4116 21140
rect 4172 21362 4228 21374
rect 4172 21310 4174 21362
rect 4226 21310 4228 21362
rect 3948 21026 4004 21084
rect 3948 20974 3950 21026
rect 4002 20974 4004 21026
rect 3948 20962 4004 20974
rect 4060 20916 4116 20926
rect 4060 20822 4116 20860
rect 3948 19908 4004 19918
rect 3836 19906 4116 19908
rect 3836 19854 3950 19906
rect 4002 19854 4116 19906
rect 3836 19852 4116 19854
rect 3612 19236 3668 19852
rect 3948 19842 4004 19852
rect 3612 19170 3668 19180
rect 3164 19012 3220 19022
rect 3612 19012 3668 19022
rect 2716 19010 3780 19012
rect 2716 18958 2718 19010
rect 2770 18958 3166 19010
rect 3218 18958 3614 19010
rect 3666 18958 3780 19010
rect 2716 18956 3780 18958
rect 2716 18946 2772 18956
rect 3164 18946 3220 18956
rect 3612 18946 3668 18956
rect 3724 18564 3780 18956
rect 3724 18470 3780 18508
rect 4060 19010 4116 19852
rect 4172 19460 4228 21310
rect 4172 19394 4228 19404
rect 4284 20020 4340 25564
rect 4844 25508 4900 26012
rect 4732 25452 4900 25508
rect 4732 24724 4788 25452
rect 4956 25396 5012 26124
rect 4844 25284 4900 25294
rect 4844 25190 4900 25228
rect 4732 24592 4788 24668
rect 4956 24610 5012 25340
rect 4956 24558 4958 24610
rect 5010 24558 5012 24610
rect 4956 24546 5012 24558
rect 5068 24388 5124 26796
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4844 24332 5124 24388
rect 4508 24162 4564 24174
rect 4508 24110 4510 24162
rect 4562 24110 4564 24162
rect 4508 24052 4564 24110
rect 4844 24052 4900 24332
rect 4508 24050 4900 24052
rect 4508 23998 4510 24050
rect 4562 23998 4900 24050
rect 4508 23996 4900 23998
rect 4508 23986 4564 23996
rect 4956 23828 5012 23838
rect 4620 23268 4676 23278
rect 4620 23174 4676 23212
rect 4956 22930 5012 23772
rect 5068 23268 5124 23278
rect 5068 23174 5124 23212
rect 4956 22878 4958 22930
rect 5010 22878 5012 22930
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4396 22594 4452 22606
rect 4396 22542 4398 22594
rect 4450 22542 4452 22594
rect 4396 22482 4452 22542
rect 4956 22594 5012 22878
rect 4956 22542 4958 22594
rect 5010 22542 5012 22594
rect 4956 22530 5012 22542
rect 4396 22430 4398 22482
rect 4450 22430 4452 22482
rect 4396 22418 4452 22430
rect 4844 22372 4900 22382
rect 4844 22278 4900 22316
rect 5068 22260 5124 22270
rect 5068 21924 5124 22204
rect 4956 21868 5124 21924
rect 4844 21588 4900 21598
rect 4844 21494 4900 21532
rect 4396 21476 4452 21486
rect 4396 21382 4452 21420
rect 4956 21252 5012 21868
rect 5180 21812 5236 28700
rect 5404 28532 5460 29374
rect 5852 29204 5908 31836
rect 5852 28754 5908 29148
rect 5852 28702 5854 28754
rect 5906 28702 5908 28754
rect 5852 28690 5908 28702
rect 5292 28084 5348 28094
rect 5404 28084 5460 28476
rect 5292 28082 5460 28084
rect 5292 28030 5294 28082
rect 5346 28030 5460 28082
rect 5292 28028 5460 28030
rect 5740 28532 5796 28542
rect 5292 28018 5348 28028
rect 5292 27300 5348 27310
rect 5292 26964 5348 27244
rect 5740 27186 5796 28476
rect 5740 27134 5742 27186
rect 5794 27134 5796 27186
rect 5740 27122 5796 27134
rect 5964 26908 6020 33740
rect 6300 33684 6356 34860
rect 6412 34132 6468 35252
rect 6636 35140 6692 37100
rect 6636 35074 6692 35084
rect 6748 35698 6804 35710
rect 6748 35646 6750 35698
rect 6802 35646 6804 35698
rect 6412 34066 6468 34076
rect 6524 34244 6580 34254
rect 6188 33628 6356 33684
rect 6412 33908 6468 33918
rect 6076 33572 6132 33582
rect 6076 33458 6132 33516
rect 6076 33406 6078 33458
rect 6130 33406 6132 33458
rect 6076 33394 6132 33406
rect 6188 33236 6244 33628
rect 6412 33346 6468 33852
rect 6412 33294 6414 33346
rect 6466 33294 6468 33346
rect 6412 33236 6468 33294
rect 6188 33180 6356 33236
rect 6076 33124 6132 33134
rect 6076 32674 6132 33068
rect 6076 32622 6078 32674
rect 6130 32622 6132 32674
rect 6076 32004 6132 32622
rect 6188 32676 6244 32686
rect 6188 32582 6244 32620
rect 6076 31938 6132 31948
rect 6300 31890 6356 33180
rect 6412 33170 6468 33180
rect 6412 32788 6468 32798
rect 6524 32788 6580 34188
rect 6748 34132 6804 35646
rect 6860 34914 6916 37212
rect 7084 37266 7140 37996
rect 7084 37214 7086 37266
rect 7138 37214 7140 37266
rect 7084 37044 7140 37214
rect 7084 36978 7140 36988
rect 7196 36932 7252 36942
rect 7196 35922 7252 36876
rect 7196 35870 7198 35922
rect 7250 35870 7252 35922
rect 7196 35858 7252 35870
rect 7308 36596 7364 38612
rect 7420 38500 7476 39454
rect 7644 39956 7700 39966
rect 7644 39618 7700 39900
rect 7756 39844 7812 39854
rect 7756 39730 7812 39788
rect 7756 39678 7758 39730
rect 7810 39678 7812 39730
rect 7756 39666 7812 39678
rect 7644 39566 7646 39618
rect 7698 39566 7700 39618
rect 7644 39396 7700 39566
rect 7644 39330 7700 39340
rect 7868 39620 7924 39630
rect 7756 39060 7812 39070
rect 7420 38434 7476 38444
rect 7644 38836 7700 38846
rect 7420 38162 7476 38174
rect 7420 38110 7422 38162
rect 7474 38110 7476 38162
rect 7420 37266 7476 38110
rect 7644 38050 7700 38780
rect 7756 38834 7812 39004
rect 7756 38782 7758 38834
rect 7810 38782 7812 38834
rect 7756 38770 7812 38782
rect 7644 37998 7646 38050
rect 7698 37998 7700 38050
rect 7644 37986 7700 37998
rect 7756 38612 7812 38622
rect 7532 37940 7588 37950
rect 7532 37846 7588 37884
rect 7756 37380 7812 38556
rect 7868 37492 7924 39564
rect 7980 39060 8036 40572
rect 7980 38994 8036 39004
rect 8092 40964 8148 40974
rect 8092 38948 8148 40908
rect 8204 39396 8260 42028
rect 8316 40962 8372 40974
rect 8316 40910 8318 40962
rect 8370 40910 8372 40962
rect 8316 40628 8372 40910
rect 8316 40562 8372 40572
rect 8316 40402 8372 40414
rect 8316 40350 8318 40402
rect 8370 40350 8372 40402
rect 8316 40292 8372 40350
rect 8428 40404 8484 42252
rect 8540 41970 8596 42476
rect 8540 41918 8542 41970
rect 8594 41918 8596 41970
rect 8540 41906 8596 41918
rect 8652 41076 8708 43372
rect 8876 43314 8932 43820
rect 8988 43428 9044 43438
rect 8988 43334 9044 43372
rect 8876 43262 8878 43314
rect 8930 43262 8932 43314
rect 8876 43250 8932 43262
rect 9100 43204 9156 43214
rect 8764 43092 8820 43102
rect 8764 42754 8820 43036
rect 8764 42702 8766 42754
rect 8818 42702 8820 42754
rect 8764 42690 8820 42702
rect 8988 42756 9044 42766
rect 8988 42662 9044 42700
rect 8876 42530 8932 42542
rect 8876 42478 8878 42530
rect 8930 42478 8932 42530
rect 8652 41010 8708 41020
rect 8764 42308 8820 42318
rect 8764 42082 8820 42252
rect 8764 42030 8766 42082
rect 8818 42030 8820 42082
rect 8652 40404 8708 40414
rect 8428 40348 8596 40404
rect 8316 40236 8484 40292
rect 8316 39396 8372 39406
rect 8204 39394 8372 39396
rect 8204 39342 8318 39394
rect 8370 39342 8372 39394
rect 8204 39340 8372 39342
rect 8316 39172 8372 39340
rect 8316 39106 8372 39116
rect 8204 38948 8260 38958
rect 8092 38946 8260 38948
rect 8092 38894 8206 38946
rect 8258 38894 8260 38946
rect 8092 38892 8260 38894
rect 8204 38882 8260 38892
rect 8316 38948 8372 38958
rect 7980 38724 8036 38762
rect 7980 38658 8036 38668
rect 8092 38722 8148 38734
rect 8092 38670 8094 38722
rect 8146 38670 8148 38722
rect 8092 38276 8148 38670
rect 8316 38668 8372 38892
rect 8428 38836 8484 40236
rect 8428 38770 8484 38780
rect 8316 38612 8484 38668
rect 8092 38210 8148 38220
rect 8204 38500 8260 38510
rect 7868 37436 8148 37492
rect 7756 37324 7924 37380
rect 7420 37214 7422 37266
rect 7474 37214 7476 37266
rect 7420 37202 7476 37214
rect 7756 37044 7812 37054
rect 7756 36708 7812 36988
rect 7868 36932 7924 37324
rect 7980 37156 8036 37166
rect 7980 37062 8036 37100
rect 7868 36876 8036 36932
rect 7308 35924 7364 36540
rect 7532 36652 7812 36708
rect 7532 36482 7588 36652
rect 7868 36596 7924 36606
rect 7868 36502 7924 36540
rect 7532 36430 7534 36482
rect 7586 36430 7588 36482
rect 7532 36418 7588 36430
rect 7980 36482 8036 36876
rect 7980 36430 7982 36482
rect 8034 36430 8036 36482
rect 7980 36418 8036 36430
rect 7308 35858 7364 35868
rect 7420 36372 7476 36382
rect 6860 34862 6862 34914
rect 6914 34862 6916 34914
rect 6860 34244 6916 34862
rect 6860 34178 6916 34188
rect 6972 35252 7028 35262
rect 6972 34690 7028 35196
rect 7196 35140 7252 35150
rect 7196 35026 7252 35084
rect 7196 34974 7198 35026
rect 7250 34974 7252 35026
rect 7196 34962 7252 34974
rect 7308 34916 7364 34926
rect 7308 34822 7364 34860
rect 6972 34638 6974 34690
rect 7026 34638 7028 34690
rect 6412 32786 6580 32788
rect 6412 32734 6414 32786
rect 6466 32734 6580 32786
rect 6412 32732 6580 32734
rect 6636 33460 6692 33470
rect 6748 33460 6804 34076
rect 6636 33458 6804 33460
rect 6636 33406 6638 33458
rect 6690 33406 6804 33458
rect 6636 33404 6804 33406
rect 6972 33460 7028 34638
rect 7196 34692 7252 34702
rect 7196 34598 7252 34636
rect 7420 34468 7476 36316
rect 7644 36370 7700 36382
rect 7644 36318 7646 36370
rect 7698 36318 7700 36370
rect 7644 36148 7700 36318
rect 7700 36092 7812 36148
rect 7644 36082 7700 36092
rect 7644 35588 7700 35598
rect 7644 35494 7700 35532
rect 7196 34412 7476 34468
rect 6412 32722 6468 32732
rect 6300 31838 6302 31890
rect 6354 31838 6356 31890
rect 6188 31780 6244 31790
rect 6188 31444 6244 31724
rect 6300 31556 6356 31838
rect 6300 31490 6356 31500
rect 6076 29652 6132 29662
rect 6076 29558 6132 29596
rect 6076 28084 6132 28094
rect 6188 28084 6244 31388
rect 6076 28082 6244 28084
rect 6076 28030 6078 28082
rect 6130 28030 6244 28082
rect 6076 28028 6244 28030
rect 6076 28018 6132 28028
rect 6188 26908 6244 28028
rect 6300 31332 6356 31342
rect 6300 30098 6356 31276
rect 6636 31332 6692 33404
rect 6972 33394 7028 33404
rect 7084 34244 7140 34254
rect 6972 32788 7028 32798
rect 6972 32338 7028 32732
rect 6972 32286 6974 32338
rect 7026 32286 7028 32338
rect 6972 32228 7028 32286
rect 6972 32162 7028 32172
rect 7084 32004 7140 34188
rect 7196 32228 7252 34412
rect 7308 34244 7364 34254
rect 7308 34242 7476 34244
rect 7308 34190 7310 34242
rect 7362 34190 7476 34242
rect 7308 34188 7476 34190
rect 7308 34178 7364 34188
rect 7420 32564 7476 34188
rect 7532 34242 7588 34254
rect 7532 34190 7534 34242
rect 7586 34190 7588 34242
rect 7532 33348 7588 34190
rect 7532 33282 7588 33292
rect 7756 33348 7812 36092
rect 8092 35924 8148 37436
rect 8204 37268 8260 38444
rect 8428 37604 8484 38612
rect 8540 38050 8596 40348
rect 8652 39732 8708 40348
rect 8764 40402 8820 42030
rect 8876 42084 8932 42478
rect 8876 42018 8932 42028
rect 8876 41860 8932 41870
rect 8876 41766 8932 41804
rect 8876 41412 8932 41422
rect 9100 41412 9156 43148
rect 9212 42756 9268 42766
rect 9212 42662 9268 42700
rect 9324 42308 9380 43932
rect 9324 42242 9380 42252
rect 8876 41410 9156 41412
rect 8876 41358 8878 41410
rect 8930 41358 9156 41410
rect 8876 41356 9156 41358
rect 8876 41346 8932 41356
rect 8988 41186 9044 41198
rect 8988 41134 8990 41186
rect 9042 41134 9044 41186
rect 8876 40628 8932 40638
rect 8988 40628 9044 41134
rect 9100 40852 9156 41356
rect 9212 41076 9268 41086
rect 9212 40982 9268 41020
rect 9436 41076 9492 44156
rect 9660 44100 9716 44110
rect 9660 43428 9716 44044
rect 9884 43764 9940 43774
rect 9996 43764 10052 47406
rect 10108 44660 10164 47964
rect 10220 47684 10276 48188
rect 10220 47618 10276 47628
rect 10332 46786 10388 48748
rect 10332 46734 10334 46786
rect 10386 46734 10388 46786
rect 10332 46116 10388 46734
rect 10444 48468 10500 48478
rect 10444 48244 10500 48412
rect 10556 48244 10612 48254
rect 10444 48242 10612 48244
rect 10444 48190 10558 48242
rect 10610 48190 10612 48242
rect 10444 48188 10612 48190
rect 10444 46340 10500 48188
rect 10556 48178 10612 48188
rect 10556 47684 10612 47694
rect 10556 47348 10612 47628
rect 10556 47282 10612 47292
rect 10668 47458 10724 48972
rect 10668 47406 10670 47458
rect 10722 47406 10724 47458
rect 10668 46898 10724 47406
rect 10668 46846 10670 46898
rect 10722 46846 10724 46898
rect 10668 46834 10724 46846
rect 10556 46788 10612 46798
rect 10556 46694 10612 46732
rect 10780 46674 10836 49756
rect 10892 49588 10948 49598
rect 10892 49494 10948 49532
rect 11004 49586 11060 49598
rect 11004 49534 11006 49586
rect 11058 49534 11060 49586
rect 11004 49028 11060 49534
rect 11004 48962 11060 48972
rect 11116 49140 11172 49150
rect 11004 48804 11060 48814
rect 11004 48710 11060 48748
rect 11004 48468 11060 48478
rect 10892 48132 10948 48142
rect 10892 47346 10948 48076
rect 10892 47294 10894 47346
rect 10946 47294 10948 47346
rect 10892 47282 10948 47294
rect 11004 47346 11060 48412
rect 11116 47572 11172 49084
rect 11340 48468 11396 50318
rect 11452 50036 11508 50046
rect 11452 49942 11508 49980
rect 11676 50036 11732 50074
rect 11676 49970 11732 49980
rect 11452 49812 11508 49822
rect 11452 49364 11508 49756
rect 11788 49810 11844 49822
rect 11788 49758 11790 49810
rect 11842 49758 11844 49810
rect 11788 49476 11844 49758
rect 11788 49410 11844 49420
rect 11452 49138 11508 49308
rect 11452 49086 11454 49138
rect 11506 49086 11508 49138
rect 11452 49074 11508 49086
rect 11676 49252 11732 49262
rect 11340 48412 11620 48468
rect 11340 48244 11396 48254
rect 11340 48150 11396 48188
rect 11452 47684 11508 47694
rect 11116 47516 11284 47572
rect 11004 47294 11006 47346
rect 11058 47294 11060 47346
rect 11004 47124 11060 47294
rect 11116 47346 11172 47358
rect 11116 47294 11118 47346
rect 11170 47294 11172 47346
rect 11116 47236 11172 47294
rect 11228 47348 11284 47516
rect 11452 47570 11508 47628
rect 11452 47518 11454 47570
rect 11506 47518 11508 47570
rect 11452 47506 11508 47518
rect 11228 47292 11508 47348
rect 11116 47170 11172 47180
rect 11004 47058 11060 47068
rect 10780 46622 10782 46674
rect 10834 46622 10836 46674
rect 10780 46340 10836 46622
rect 10444 46284 10612 46340
rect 10332 46060 10500 46116
rect 10332 45890 10388 45902
rect 10332 45838 10334 45890
rect 10386 45838 10388 45890
rect 10108 44594 10164 44604
rect 10220 44994 10276 45006
rect 10220 44942 10222 44994
rect 10274 44942 10276 44994
rect 10220 44436 10276 44942
rect 10332 44996 10388 45838
rect 10444 45108 10500 46060
rect 10444 45042 10500 45052
rect 10332 44930 10388 44940
rect 10220 44370 10276 44380
rect 10332 44324 10388 44334
rect 9884 43762 10052 43764
rect 9884 43710 9886 43762
rect 9938 43710 10052 43762
rect 9884 43708 10052 43710
rect 10220 44212 10276 44222
rect 9884 43698 9940 43708
rect 9772 43652 9828 43662
rect 9772 43558 9828 43596
rect 10220 43540 10276 44156
rect 10332 43764 10388 44268
rect 10444 44212 10500 44222
rect 10444 44118 10500 44156
rect 10332 43698 10388 43708
rect 10444 43652 10500 43662
rect 10444 43558 10500 43596
rect 10220 43484 10388 43540
rect 9996 43428 10052 43438
rect 9660 43426 10052 43428
rect 9660 43374 9998 43426
rect 10050 43374 10052 43426
rect 9660 43372 10052 43374
rect 9996 43362 10052 43372
rect 10220 43316 10276 43326
rect 10220 43222 10276 43260
rect 9660 42868 9716 42878
rect 9660 41970 9716 42812
rect 10332 42866 10388 43484
rect 10332 42814 10334 42866
rect 10386 42814 10388 42866
rect 9884 42644 9940 42654
rect 9884 42196 9940 42588
rect 10332 42532 10388 42814
rect 10332 42466 10388 42476
rect 10556 42308 10612 46284
rect 10780 45780 10836 46284
rect 11004 46900 11060 46910
rect 10892 45780 10948 45790
rect 10780 45778 10948 45780
rect 10780 45726 10894 45778
rect 10946 45726 10948 45778
rect 10780 45724 10948 45726
rect 10892 45714 10948 45724
rect 11004 45556 11060 46844
rect 11452 46898 11508 47292
rect 11564 47012 11620 48412
rect 11564 46946 11620 46956
rect 11452 46846 11454 46898
rect 11506 46846 11508 46898
rect 11452 46834 11508 46846
rect 10892 45500 11060 45556
rect 11340 46788 11396 46798
rect 10780 45332 10836 45342
rect 10780 45238 10836 45276
rect 10780 45108 10836 45118
rect 10780 45014 10836 45052
rect 10668 44434 10724 44446
rect 10668 44382 10670 44434
rect 10722 44382 10724 44434
rect 10668 43538 10724 44382
rect 10668 43486 10670 43538
rect 10722 43486 10724 43538
rect 10668 42756 10724 43486
rect 10668 42690 10724 42700
rect 10332 42252 10612 42308
rect 10668 42420 10724 42430
rect 10108 42196 10164 42206
rect 9884 42194 10164 42196
rect 9884 42142 10110 42194
rect 10162 42142 10164 42194
rect 9884 42140 10164 42142
rect 9660 41918 9662 41970
rect 9714 41918 9716 41970
rect 9660 41906 9716 41918
rect 10108 41524 10164 42140
rect 10108 41458 10164 41468
rect 9548 41300 9604 41310
rect 9548 41186 9604 41244
rect 9884 41300 9940 41310
rect 9884 41298 10052 41300
rect 9884 41246 9886 41298
rect 9938 41246 10052 41298
rect 9884 41244 10052 41246
rect 9884 41234 9940 41244
rect 9548 41134 9550 41186
rect 9602 41134 9604 41186
rect 9548 41122 9604 41134
rect 9100 40796 9380 40852
rect 8876 40626 9044 40628
rect 8876 40574 8878 40626
rect 8930 40574 9044 40626
rect 8876 40572 9044 40574
rect 8876 40562 8932 40572
rect 8764 40350 8766 40402
rect 8818 40350 8820 40402
rect 8764 40180 8820 40350
rect 8988 40402 9044 40414
rect 8988 40350 8990 40402
rect 9042 40350 9044 40402
rect 8988 40292 9044 40350
rect 8988 40236 9268 40292
rect 8764 40124 9156 40180
rect 8764 39732 8820 39742
rect 8652 39730 8820 39732
rect 8652 39678 8766 39730
rect 8818 39678 8820 39730
rect 8652 39676 8820 39678
rect 8652 38388 8708 38398
rect 8652 38162 8708 38332
rect 8652 38110 8654 38162
rect 8706 38110 8708 38162
rect 8652 38098 8708 38110
rect 8764 38164 8820 39676
rect 8988 39060 9044 39070
rect 8988 38966 9044 39004
rect 9100 38668 9156 40124
rect 8764 38098 8820 38108
rect 8876 38612 9156 38668
rect 9212 39730 9268 40236
rect 9212 39678 9214 39730
rect 9266 39678 9268 39730
rect 9212 38724 9268 39678
rect 9212 38658 9268 38668
rect 9324 38612 9380 40796
rect 9436 40404 9492 41020
rect 9772 41074 9828 41086
rect 9772 41022 9774 41074
rect 9826 41022 9828 41074
rect 9772 40964 9828 41022
rect 9828 40908 9940 40964
rect 9772 40898 9828 40908
rect 9436 40348 9604 40404
rect 8540 37998 8542 38050
rect 8594 37998 8596 38050
rect 8540 37986 8596 37998
rect 8764 37938 8820 37950
rect 8764 37886 8766 37938
rect 8818 37886 8820 37938
rect 8428 37548 8596 37604
rect 8428 37378 8484 37390
rect 8428 37326 8430 37378
rect 8482 37326 8484 37378
rect 8204 37266 8372 37268
rect 8204 37214 8206 37266
rect 8258 37214 8372 37266
rect 8204 37212 8372 37214
rect 8204 37202 8260 37212
rect 7980 35868 8148 35924
rect 7756 33282 7812 33292
rect 7868 35474 7924 35486
rect 7868 35422 7870 35474
rect 7922 35422 7924 35474
rect 7868 33236 7924 35422
rect 7980 34804 8036 35868
rect 8204 35586 8260 35598
rect 8204 35534 8206 35586
rect 8258 35534 8260 35586
rect 8204 35474 8260 35534
rect 8204 35422 8206 35474
rect 8258 35422 8260 35474
rect 8204 35410 8260 35422
rect 7980 34710 8036 34748
rect 8316 34802 8372 37212
rect 8428 36596 8484 37326
rect 8428 36530 8484 36540
rect 8540 36148 8596 37548
rect 8764 37268 8820 37886
rect 8764 37202 8820 37212
rect 8652 36932 8708 36942
rect 8652 36708 8708 36876
rect 8652 36642 8708 36652
rect 8764 36484 8820 36494
rect 8540 36082 8596 36092
rect 8652 36482 8820 36484
rect 8652 36430 8766 36482
rect 8818 36430 8820 36482
rect 8652 36428 8820 36430
rect 8540 35924 8596 35934
rect 8540 35830 8596 35868
rect 8316 34750 8318 34802
rect 8370 34750 8372 34802
rect 8092 34692 8148 34702
rect 8092 34598 8148 34636
rect 8204 34690 8260 34702
rect 8204 34638 8206 34690
rect 8258 34638 8260 34690
rect 8204 34468 8260 34638
rect 7868 32900 7924 33180
rect 7644 32676 7700 32686
rect 7420 32562 7588 32564
rect 7420 32510 7422 32562
rect 7474 32510 7588 32562
rect 7420 32508 7588 32510
rect 7420 32498 7476 32508
rect 7196 32172 7364 32228
rect 6860 31948 7140 32004
rect 7196 32004 7252 32014
rect 6636 31266 6692 31276
rect 6748 31778 6804 31790
rect 6748 31726 6750 31778
rect 6802 31726 6804 31778
rect 6636 30994 6692 31006
rect 6636 30942 6638 30994
rect 6690 30942 6692 30994
rect 6636 30548 6692 30942
rect 6300 30046 6302 30098
rect 6354 30046 6356 30098
rect 6300 27188 6356 30046
rect 6524 30098 6580 30110
rect 6524 30046 6526 30098
rect 6578 30046 6580 30098
rect 6412 28756 6468 28766
rect 6412 28662 6468 28700
rect 6524 27972 6580 30046
rect 6524 27906 6580 27916
rect 6300 27122 6356 27132
rect 5292 26898 5348 26908
rect 5852 26852 6020 26908
rect 6076 26852 6244 26908
rect 6524 26964 6580 26974
rect 6636 26964 6692 30492
rect 6748 30884 6804 31726
rect 6748 29426 6804 30828
rect 6860 30434 6916 31948
rect 7084 31778 7140 31790
rect 7084 31726 7086 31778
rect 7138 31726 7140 31778
rect 7084 30996 7140 31726
rect 7084 30864 7140 30940
rect 7196 31106 7252 31948
rect 7196 31054 7198 31106
rect 7250 31054 7252 31106
rect 7196 30436 7252 31054
rect 7308 30884 7364 32172
rect 7532 31556 7588 32508
rect 7644 32562 7700 32620
rect 7644 32510 7646 32562
rect 7698 32510 7700 32562
rect 7644 32498 7700 32510
rect 7756 31780 7812 31790
rect 7756 31686 7812 31724
rect 7868 31778 7924 32844
rect 7868 31726 7870 31778
rect 7922 31726 7924 31778
rect 7644 31556 7700 31566
rect 7532 31500 7644 31556
rect 7644 31462 7700 31500
rect 7308 30752 7364 30828
rect 6860 30382 6862 30434
rect 6914 30382 6916 30434
rect 6860 29540 6916 30382
rect 6860 29474 6916 29484
rect 6972 30380 7252 30436
rect 6748 29374 6750 29426
rect 6802 29374 6804 29426
rect 6748 29362 6804 29374
rect 6972 27858 7028 30380
rect 7196 30212 7252 30222
rect 7196 30118 7252 30156
rect 7868 29988 7924 31726
rect 7980 34412 8260 34468
rect 7980 33908 8036 34412
rect 8092 34244 8148 34254
rect 8092 34130 8148 34188
rect 8204 34244 8260 34254
rect 8316 34244 8372 34750
rect 8204 34242 8372 34244
rect 8204 34190 8206 34242
rect 8258 34190 8372 34242
rect 8204 34188 8372 34190
rect 8428 34804 8484 34814
rect 8652 34804 8708 36428
rect 8764 36418 8820 36428
rect 8428 34802 8708 34804
rect 8428 34750 8430 34802
rect 8482 34750 8708 34802
rect 8428 34748 8708 34750
rect 8764 35028 8820 35038
rect 8204 34178 8260 34188
rect 8092 34078 8094 34130
rect 8146 34078 8148 34130
rect 8092 34066 8148 34078
rect 7980 31668 8036 33852
rect 8428 33796 8484 34748
rect 8540 34468 8596 34478
rect 8540 34354 8596 34412
rect 8540 34302 8542 34354
rect 8594 34302 8596 34354
rect 8540 34290 8596 34302
rect 8428 33730 8484 33740
rect 8092 33460 8148 33470
rect 8092 33366 8148 33404
rect 8540 33122 8596 33134
rect 8540 33070 8542 33122
rect 8594 33070 8596 33122
rect 8540 32900 8596 33070
rect 8540 32834 8596 32844
rect 8428 32788 8484 32798
rect 8428 32676 8484 32732
rect 8540 32676 8596 32686
rect 8428 32674 8596 32676
rect 8428 32622 8542 32674
rect 8594 32622 8596 32674
rect 8428 32620 8596 32622
rect 8540 32610 8596 32620
rect 8092 32452 8148 32462
rect 8148 32396 8260 32452
rect 8092 32358 8148 32396
rect 7980 31602 8036 31612
rect 8092 31554 8148 31566
rect 8092 31502 8094 31554
rect 8146 31502 8148 31554
rect 8092 31332 8148 31502
rect 8092 31266 8148 31276
rect 7980 30212 8036 30222
rect 7980 30118 8036 30156
rect 7756 29932 7924 29988
rect 7084 28532 7140 28542
rect 7084 28438 7140 28476
rect 6972 27806 6974 27858
rect 7026 27806 7028 27858
rect 6972 27636 7028 27806
rect 6972 27570 7028 27580
rect 7532 27972 7588 27982
rect 6748 27076 6804 27086
rect 6748 26982 6804 27020
rect 7084 27076 7140 27086
rect 6580 26908 6692 26964
rect 5292 26740 5348 26750
rect 5292 22260 5348 26684
rect 5404 26292 5460 26302
rect 5404 26198 5460 26236
rect 5852 25618 5908 26852
rect 5964 26290 6020 26302
rect 5964 26238 5966 26290
rect 6018 26238 6020 26290
rect 5964 26180 6020 26238
rect 5964 26114 6020 26124
rect 5852 25566 5854 25618
rect 5906 25566 5908 25618
rect 5852 25554 5908 25566
rect 5740 25172 5796 25182
rect 5740 24834 5796 25116
rect 5740 24782 5742 24834
rect 5794 24782 5796 24834
rect 5740 24052 5796 24782
rect 5628 23380 5684 23390
rect 5628 23286 5684 23324
rect 5292 22194 5348 22204
rect 5516 23268 5572 23278
rect 5404 21812 5460 21822
rect 5180 21810 5460 21812
rect 5180 21758 5406 21810
rect 5458 21758 5460 21810
rect 5180 21756 5460 21758
rect 5404 21746 5460 21756
rect 5516 21588 5572 23212
rect 5740 22484 5796 23996
rect 5740 22418 5796 22428
rect 5964 23380 6020 23390
rect 6076 23380 6132 26852
rect 6300 25732 6356 25742
rect 6300 23940 6356 25676
rect 6412 25508 6468 25518
rect 6524 25508 6580 26908
rect 6748 26068 6804 26078
rect 6748 25618 6804 26012
rect 6748 25566 6750 25618
rect 6802 25566 6804 25618
rect 6748 25554 6804 25566
rect 6412 25506 6580 25508
rect 6412 25454 6414 25506
rect 6466 25454 6580 25506
rect 6412 25452 6580 25454
rect 6412 25442 6468 25452
rect 6524 24164 6580 25452
rect 6972 24724 7028 24734
rect 6972 24630 7028 24668
rect 7084 24722 7140 27020
rect 7308 27074 7364 27086
rect 7308 27022 7310 27074
rect 7362 27022 7364 27074
rect 7308 26180 7364 27022
rect 7308 26114 7364 26124
rect 7532 26178 7588 27916
rect 7756 26908 7812 29932
rect 7868 29426 7924 29438
rect 7868 29374 7870 29426
rect 7922 29374 7924 29426
rect 7868 28980 7924 29374
rect 7868 28914 7924 28924
rect 7980 28532 8036 28542
rect 7980 28418 8036 28476
rect 7980 28366 7982 28418
rect 8034 28366 8036 28418
rect 7980 27524 8036 28366
rect 8092 28308 8148 28318
rect 8092 27860 8148 28252
rect 8092 27746 8148 27804
rect 8092 27694 8094 27746
rect 8146 27694 8148 27746
rect 8092 27682 8148 27694
rect 7980 27458 8036 27468
rect 8204 26908 8260 32396
rect 8652 31668 8708 31678
rect 8652 31574 8708 31612
rect 8540 31220 8596 31230
rect 8428 30996 8484 31006
rect 8428 30436 8484 30940
rect 8540 30994 8596 31164
rect 8764 30996 8820 34972
rect 8876 33460 8932 38612
rect 9324 38546 9380 38556
rect 9436 40180 9492 40190
rect 8988 38276 9044 38286
rect 8988 38182 9044 38220
rect 9100 38052 9156 38062
rect 9100 37958 9156 37996
rect 9212 37940 9268 37950
rect 9212 37716 9268 37884
rect 9212 36484 9268 37660
rect 9436 36820 9492 40124
rect 9548 37044 9604 40348
rect 9772 40290 9828 40302
rect 9772 40238 9774 40290
rect 9826 40238 9828 40290
rect 9772 40180 9828 40238
rect 9772 40114 9828 40124
rect 9772 39844 9828 39854
rect 9884 39844 9940 40908
rect 9772 39842 9940 39844
rect 9772 39790 9774 39842
rect 9826 39790 9940 39842
rect 9772 39788 9940 39790
rect 9772 39778 9828 39788
rect 9884 39620 9940 39630
rect 9884 39526 9940 39564
rect 9996 38948 10052 41244
rect 10220 40178 10276 40190
rect 10220 40126 10222 40178
rect 10274 40126 10276 40178
rect 10108 39732 10164 39742
rect 10108 39506 10164 39676
rect 10108 39454 10110 39506
rect 10162 39454 10164 39506
rect 10108 39442 10164 39454
rect 10220 39620 10276 40126
rect 10220 39284 10276 39564
rect 10332 39396 10388 42252
rect 10668 42194 10724 42364
rect 10668 42142 10670 42194
rect 10722 42142 10724 42194
rect 10668 42130 10724 42142
rect 10556 41410 10612 41422
rect 10556 41358 10558 41410
rect 10610 41358 10612 41410
rect 10556 40404 10612 41358
rect 10668 41188 10724 41198
rect 10668 41094 10724 41132
rect 10556 40338 10612 40348
rect 10556 40180 10612 40218
rect 10612 40124 10724 40180
rect 10556 40114 10612 40124
rect 10444 40068 10500 40078
rect 10444 39618 10500 40012
rect 10444 39566 10446 39618
rect 10498 39566 10500 39618
rect 10444 39554 10500 39566
rect 10668 39618 10724 40124
rect 10892 39956 10948 45500
rect 11340 45218 11396 46732
rect 11452 46450 11508 46462
rect 11452 46398 11454 46450
rect 11506 46398 11508 46450
rect 11452 46340 11508 46398
rect 11452 46274 11508 46284
rect 11564 46452 11620 46462
rect 11676 46452 11732 49196
rect 11788 48468 11844 48478
rect 11788 48374 11844 48412
rect 11788 46788 11844 46798
rect 11788 46674 11844 46732
rect 11788 46622 11790 46674
rect 11842 46622 11844 46674
rect 11788 46610 11844 46622
rect 11564 46450 11732 46452
rect 11564 46398 11566 46450
rect 11618 46398 11732 46450
rect 11564 46396 11732 46398
rect 11340 45166 11342 45218
rect 11394 45166 11396 45218
rect 11340 44772 11396 45166
rect 11116 44716 11396 44772
rect 11452 45780 11508 45790
rect 11452 45108 11508 45724
rect 11116 44212 11172 44716
rect 11228 44324 11284 44334
rect 11452 44324 11508 45052
rect 11228 44322 11508 44324
rect 11228 44270 11230 44322
rect 11282 44270 11508 44322
rect 11228 44268 11508 44270
rect 11564 44324 11620 46396
rect 11676 46228 11732 46238
rect 11676 45220 11732 46172
rect 11676 45108 11732 45164
rect 11676 45106 11844 45108
rect 11676 45054 11678 45106
rect 11730 45054 11844 45106
rect 11676 45052 11844 45054
rect 11676 45042 11732 45052
rect 11788 44324 11844 45052
rect 11228 44258 11284 44268
rect 11564 44258 11620 44268
rect 11676 44322 11844 44324
rect 11676 44270 11790 44322
rect 11842 44270 11844 44322
rect 11676 44268 11844 44270
rect 11116 42642 11172 44156
rect 11564 43764 11620 43774
rect 11452 43652 11508 43662
rect 11452 43558 11508 43596
rect 11116 42590 11118 42642
rect 11170 42590 11172 42642
rect 11116 41410 11172 42590
rect 11228 42868 11284 42878
rect 11564 42868 11620 43708
rect 11228 42084 11284 42812
rect 11452 42812 11620 42868
rect 11452 42196 11508 42812
rect 11564 42644 11620 42654
rect 11676 42644 11732 44268
rect 11788 44258 11844 44268
rect 11900 44098 11956 53116
rect 12012 48132 12068 54460
rect 12236 54292 12292 55804
rect 12572 55468 12628 58268
rect 12684 58258 12740 58268
rect 12796 58212 12852 58222
rect 12796 58118 12852 58156
rect 12796 57540 12852 57550
rect 12796 57446 12852 57484
rect 13132 57428 13188 57438
rect 12684 56642 12740 56654
rect 12684 56590 12686 56642
rect 12738 56590 12740 56642
rect 12684 55636 12740 56590
rect 12908 56642 12964 56654
rect 12908 56590 12910 56642
rect 12962 56590 12964 56642
rect 12908 56308 12964 56590
rect 13020 56642 13076 56654
rect 13020 56590 13022 56642
rect 13074 56590 13076 56642
rect 13020 56532 13076 56590
rect 13020 56466 13076 56476
rect 12796 56196 12852 56206
rect 12796 56102 12852 56140
rect 12908 55636 12964 56252
rect 12908 55580 13076 55636
rect 12684 55570 12740 55580
rect 12572 55412 12852 55468
rect 12908 55412 12964 55422
rect 12796 55410 12964 55412
rect 12796 55358 12910 55410
rect 12962 55358 12964 55410
rect 12796 55356 12964 55358
rect 12908 55346 12964 55356
rect 12460 55298 12516 55310
rect 12460 55246 12462 55298
rect 12514 55246 12516 55298
rect 12236 53842 12292 54236
rect 12236 53790 12238 53842
rect 12290 53790 12292 53842
rect 12236 53778 12292 53790
rect 12348 54402 12404 54414
rect 12348 54350 12350 54402
rect 12402 54350 12404 54402
rect 12348 54290 12404 54350
rect 12460 54404 12516 55246
rect 13020 55188 13076 55580
rect 12908 55132 13076 55188
rect 12908 54404 12964 55132
rect 12460 54402 12964 54404
rect 12460 54350 12910 54402
rect 12962 54350 12964 54402
rect 12460 54348 12964 54350
rect 12908 54338 12964 54348
rect 13020 54740 13076 54750
rect 13132 54740 13188 57372
rect 13468 56756 13524 58940
rect 13692 59106 13748 59118
rect 13692 59054 13694 59106
rect 13746 59054 13748 59106
rect 13692 57540 13748 59054
rect 13916 59108 13972 59118
rect 13804 58436 13860 58446
rect 13804 58342 13860 58380
rect 13692 57474 13748 57484
rect 13804 57650 13860 57662
rect 13804 57598 13806 57650
rect 13858 57598 13860 57650
rect 13692 57316 13748 57326
rect 13580 57092 13636 57102
rect 13580 56978 13636 57036
rect 13580 56926 13582 56978
rect 13634 56926 13636 56978
rect 13580 56914 13636 56926
rect 13468 56700 13636 56756
rect 13468 56532 13524 56542
rect 13020 54738 13188 54740
rect 13020 54686 13022 54738
rect 13074 54686 13188 54738
rect 13020 54684 13188 54686
rect 13244 56420 13300 56430
rect 12348 54238 12350 54290
rect 12402 54238 12404 54290
rect 12348 52948 12404 54238
rect 12348 52882 12404 52892
rect 12460 54068 12516 54078
rect 12236 52834 12292 52846
rect 12236 52782 12238 52834
rect 12290 52782 12292 52834
rect 12124 52722 12180 52734
rect 12124 52670 12126 52722
rect 12178 52670 12180 52722
rect 12124 51154 12180 52670
rect 12236 52612 12292 52782
rect 12236 52546 12292 52556
rect 12460 52164 12516 54012
rect 12572 53732 12628 53742
rect 12572 53638 12628 53676
rect 13020 53508 13076 54684
rect 13244 54626 13300 56364
rect 13468 56194 13524 56476
rect 13468 56142 13470 56194
rect 13522 56142 13524 56194
rect 13468 56130 13524 56142
rect 13580 55972 13636 56700
rect 13468 55916 13636 55972
rect 13692 56194 13748 57260
rect 13692 56142 13694 56194
rect 13746 56142 13748 56194
rect 13244 54574 13246 54626
rect 13298 54574 13300 54626
rect 13244 53956 13300 54574
rect 13356 55412 13412 55422
rect 13356 54516 13412 55356
rect 13356 54450 13412 54460
rect 13244 53890 13300 53900
rect 12908 53452 13076 53508
rect 13468 53508 13524 55916
rect 13692 55188 13748 56142
rect 13804 55410 13860 57598
rect 13804 55358 13806 55410
rect 13858 55358 13860 55410
rect 13804 55346 13860 55358
rect 13916 55300 13972 59052
rect 14028 58884 14084 59726
rect 14364 59220 14420 59836
rect 14364 59126 14420 59164
rect 14588 59218 14644 59950
rect 14700 59892 14756 59902
rect 14700 59798 14756 59836
rect 15036 59890 15092 59902
rect 15036 59838 15038 59890
rect 15090 59838 15092 59890
rect 14924 59780 14980 59790
rect 14924 59686 14980 59724
rect 14588 59166 14590 59218
rect 14642 59166 14644 59218
rect 14588 58884 14644 59166
rect 14700 59220 14756 59230
rect 15036 59220 15092 59838
rect 15708 59778 15764 59790
rect 15708 59726 15710 59778
rect 15762 59726 15764 59778
rect 15708 59668 15764 59726
rect 15708 59602 15764 59612
rect 15932 59780 15988 59790
rect 14700 59218 15092 59220
rect 14700 59166 14702 59218
rect 14754 59166 15092 59218
rect 14700 59164 15092 59166
rect 15932 59442 15988 59724
rect 15932 59390 15934 59442
rect 15986 59390 15988 59442
rect 14700 59154 14756 59164
rect 14028 58818 14084 58828
rect 14364 58828 14644 58884
rect 14028 58434 14084 58446
rect 14028 58382 14030 58434
rect 14082 58382 14084 58434
rect 14028 58212 14084 58382
rect 14028 56644 14084 58156
rect 14364 57762 14420 58828
rect 14812 58436 14868 59164
rect 15148 58996 15204 59006
rect 15708 58996 15764 59006
rect 15148 58994 15764 58996
rect 15148 58942 15150 58994
rect 15202 58942 15710 58994
rect 15762 58942 15764 58994
rect 15148 58940 15764 58942
rect 15148 58930 15204 58940
rect 15708 58930 15764 58940
rect 15932 58884 15988 59390
rect 16156 59778 16212 59790
rect 16604 59780 16660 59790
rect 16156 59726 16158 59778
rect 16210 59726 16212 59778
rect 16044 59108 16100 59118
rect 16044 59014 16100 59052
rect 16156 58828 16212 59726
rect 15932 58818 15988 58828
rect 16044 58772 16212 58828
rect 16380 59778 16660 59780
rect 16380 59726 16606 59778
rect 16658 59726 16660 59778
rect 16380 59724 16660 59726
rect 15148 58436 15204 58446
rect 14812 58434 15204 58436
rect 14812 58382 15150 58434
rect 15202 58382 15204 58434
rect 14812 58380 15204 58382
rect 15148 58370 15204 58380
rect 14700 58324 14756 58334
rect 14700 58230 14756 58268
rect 15484 58324 15540 58334
rect 15484 58230 15540 58268
rect 15372 58210 15428 58222
rect 15372 58158 15374 58210
rect 15426 58158 15428 58210
rect 14364 57710 14366 57762
rect 14418 57710 14420 57762
rect 14364 57698 14420 57710
rect 14924 57876 14980 57886
rect 14252 57650 14308 57662
rect 14252 57598 14254 57650
rect 14306 57598 14308 57650
rect 14140 56868 14196 56878
rect 14140 56774 14196 56812
rect 14028 56588 14196 56644
rect 14028 55972 14084 55982
rect 14028 55524 14084 55916
rect 14140 55860 14196 56588
rect 14252 56196 14308 57598
rect 14924 57540 14980 57820
rect 14924 57446 14980 57484
rect 15260 57764 15316 57774
rect 15372 57764 15428 58158
rect 15372 57708 15540 57764
rect 14812 56980 14868 56990
rect 14364 56868 14420 56878
rect 14364 56306 14420 56812
rect 14588 56644 14644 56654
rect 14588 56550 14644 56588
rect 14364 56254 14366 56306
rect 14418 56254 14420 56306
rect 14364 56242 14420 56254
rect 14252 56082 14308 56140
rect 14252 56030 14254 56082
rect 14306 56030 14308 56082
rect 14252 56018 14308 56030
rect 14140 55804 14308 55860
rect 14140 55524 14196 55534
rect 14028 55522 14196 55524
rect 14028 55470 14142 55522
rect 14194 55470 14196 55522
rect 14028 55468 14196 55470
rect 13916 55244 14084 55300
rect 13804 55188 13860 55198
rect 13692 55132 13804 55188
rect 13860 55132 13972 55188
rect 13804 55056 13860 55132
rect 13916 55074 13972 55132
rect 13916 55022 13918 55074
rect 13970 55022 13972 55074
rect 13916 55010 13972 55022
rect 14028 54852 14084 55244
rect 13916 54796 14084 54852
rect 13804 54514 13860 54526
rect 13804 54462 13806 54514
rect 13858 54462 13860 54514
rect 13692 53842 13748 53854
rect 13692 53790 13694 53842
rect 13746 53790 13748 53842
rect 13692 53732 13748 53790
rect 13692 53666 13748 53676
rect 13468 53452 13748 53508
rect 12908 53396 12964 53452
rect 12684 53172 12740 53182
rect 12684 53078 12740 53116
rect 12460 52070 12516 52108
rect 12460 51940 12516 51950
rect 12124 51102 12126 51154
rect 12178 51102 12180 51154
rect 12124 50818 12180 51102
rect 12124 50766 12126 50818
rect 12178 50766 12180 50818
rect 12124 50754 12180 50766
rect 12348 51828 12404 51838
rect 12236 50708 12292 50718
rect 12236 50614 12292 50652
rect 12348 50482 12404 51772
rect 12348 50430 12350 50482
rect 12402 50430 12404 50482
rect 12348 50428 12404 50430
rect 12124 50372 12404 50428
rect 12460 51602 12516 51884
rect 12460 51550 12462 51602
rect 12514 51550 12516 51602
rect 12124 49252 12180 50372
rect 12460 50148 12516 51550
rect 12908 51492 12964 53340
rect 13132 52836 13188 52846
rect 13132 52742 13188 52780
rect 13468 52836 13524 52846
rect 13132 52500 13188 52510
rect 13020 52164 13076 52174
rect 13020 52070 13076 52108
rect 13020 51492 13076 51502
rect 12908 51490 13076 51492
rect 12908 51438 13022 51490
rect 13074 51438 13076 51490
rect 12908 51436 13076 51438
rect 13020 51426 13076 51436
rect 12796 51156 12852 51166
rect 12796 51154 12964 51156
rect 12796 51102 12798 51154
rect 12850 51102 12964 51154
rect 12796 51100 12964 51102
rect 12796 51090 12852 51100
rect 12236 50092 12516 50148
rect 12572 51044 12628 51054
rect 12236 49588 12292 50092
rect 12460 49924 12516 49934
rect 12572 49924 12628 50988
rect 12908 50706 12964 51100
rect 12908 50654 12910 50706
rect 12962 50654 12964 50706
rect 12684 50596 12740 50606
rect 12684 50034 12740 50540
rect 12684 49982 12686 50034
rect 12738 49982 12740 50034
rect 12684 49970 12740 49982
rect 12516 49868 12628 49924
rect 12460 49830 12516 49868
rect 12348 49812 12404 49822
rect 12348 49718 12404 49756
rect 12796 49588 12852 49598
rect 12236 49532 12516 49588
rect 12124 49196 12292 49252
rect 12124 49026 12180 49038
rect 12124 48974 12126 49026
rect 12178 48974 12180 49026
rect 12124 48804 12180 48974
rect 12124 48738 12180 48748
rect 12236 48692 12292 49196
rect 12348 49140 12404 49150
rect 12348 49046 12404 49084
rect 12236 48466 12292 48636
rect 12236 48414 12238 48466
rect 12290 48414 12292 48466
rect 12236 48402 12292 48414
rect 12012 48066 12068 48076
rect 12012 47682 12068 47694
rect 12012 47630 12014 47682
rect 12066 47630 12068 47682
rect 12012 47570 12068 47630
rect 12012 47518 12014 47570
rect 12066 47518 12068 47570
rect 12012 47506 12068 47518
rect 12460 47460 12516 49532
rect 12572 49028 12628 49038
rect 12572 48802 12628 48972
rect 12796 49026 12852 49532
rect 12796 48974 12798 49026
rect 12850 48974 12852 49026
rect 12796 48962 12852 48974
rect 12572 48750 12574 48802
rect 12626 48750 12628 48802
rect 12572 48244 12628 48750
rect 12684 48804 12740 48814
rect 12684 48710 12740 48748
rect 12908 48468 12964 50654
rect 13132 50428 13188 52444
rect 12572 48178 12628 48188
rect 12684 48412 12964 48468
rect 13020 50372 13188 50428
rect 12348 47404 12516 47460
rect 12236 47012 12292 47022
rect 12236 46676 12292 46956
rect 12348 46900 12404 47404
rect 12460 47236 12516 47246
rect 12460 47234 12628 47236
rect 12460 47182 12462 47234
rect 12514 47182 12628 47234
rect 12460 47180 12628 47182
rect 12460 47170 12516 47180
rect 12348 46844 12516 46900
rect 12348 46676 12404 46686
rect 12236 46674 12404 46676
rect 12236 46622 12350 46674
rect 12402 46622 12404 46674
rect 12236 46620 12404 46622
rect 12124 46004 12180 46014
rect 12124 45910 12180 45948
rect 12348 44884 12404 46620
rect 12348 44818 12404 44828
rect 12012 44324 12068 44334
rect 12012 44230 12068 44268
rect 12236 44324 12292 44334
rect 11900 44046 11902 44098
rect 11954 44046 11956 44098
rect 11788 43876 11844 43886
rect 11788 42980 11844 43820
rect 11900 43540 11956 44046
rect 12236 43650 12292 44268
rect 12236 43598 12238 43650
rect 12290 43598 12292 43650
rect 12236 43586 12292 43598
rect 12348 43988 12404 43998
rect 12348 43650 12404 43932
rect 12460 43764 12516 46844
rect 12572 45780 12628 47180
rect 12684 46228 12740 48412
rect 12796 48242 12852 48254
rect 12796 48190 12798 48242
rect 12850 48190 12852 48242
rect 12796 46900 12852 48190
rect 12908 48244 12964 48254
rect 12908 48150 12964 48188
rect 12908 47682 12964 47694
rect 12908 47630 12910 47682
rect 12962 47630 12964 47682
rect 12908 47348 12964 47630
rect 13020 47572 13076 50372
rect 13132 49810 13188 49822
rect 13132 49758 13134 49810
rect 13186 49758 13188 49810
rect 13132 49588 13188 49758
rect 13356 49810 13412 49822
rect 13356 49758 13358 49810
rect 13410 49758 13412 49810
rect 13244 49700 13300 49710
rect 13244 49606 13300 49644
rect 13132 49522 13188 49532
rect 13356 49028 13412 49758
rect 13356 48962 13412 48972
rect 13132 48244 13188 48254
rect 13132 48242 13300 48244
rect 13132 48190 13134 48242
rect 13186 48190 13300 48242
rect 13132 48188 13300 48190
rect 13132 48178 13188 48188
rect 13020 47570 13188 47572
rect 13020 47518 13022 47570
rect 13074 47518 13188 47570
rect 13020 47516 13188 47518
rect 13020 47506 13076 47516
rect 12908 47292 13076 47348
rect 12908 46900 12964 46910
rect 12796 46898 12964 46900
rect 12796 46846 12910 46898
rect 12962 46846 12964 46898
rect 12796 46844 12964 46846
rect 12908 46834 12964 46844
rect 12684 46162 12740 46172
rect 12796 46674 12852 46686
rect 12796 46622 12798 46674
rect 12850 46622 12852 46674
rect 12684 46004 12740 46014
rect 12684 45910 12740 45948
rect 12796 45892 12852 46622
rect 12796 45826 12852 45836
rect 13020 46674 13076 47292
rect 13020 46622 13022 46674
rect 13074 46622 13076 46674
rect 12572 45724 12740 45780
rect 12684 45332 12740 45724
rect 12572 45106 12628 45118
rect 12572 45054 12574 45106
rect 12626 45054 12628 45106
rect 12572 44884 12628 45054
rect 12572 44818 12628 44828
rect 12684 44100 12740 45276
rect 12796 45220 12852 45230
rect 12796 45126 12852 45164
rect 12684 44034 12740 44044
rect 13020 43876 13076 46622
rect 13132 44212 13188 47516
rect 13244 45668 13300 48188
rect 13356 48242 13412 48254
rect 13356 48190 13358 48242
rect 13410 48190 13412 48242
rect 13356 48132 13412 48190
rect 13356 48066 13412 48076
rect 13468 45780 13524 52780
rect 13692 51492 13748 53452
rect 13804 53506 13860 54462
rect 13804 53454 13806 53506
rect 13858 53454 13860 53506
rect 13804 53284 13860 53454
rect 13916 53508 13972 54796
rect 14140 54740 14196 55468
rect 14028 54628 14084 54638
rect 14028 54534 14084 54572
rect 14140 54626 14196 54684
rect 14140 54574 14142 54626
rect 14194 54574 14196 54626
rect 14140 54562 14196 54574
rect 14252 54628 14308 55804
rect 14252 54562 14308 54572
rect 14476 55522 14532 55534
rect 14476 55470 14478 55522
rect 14530 55470 14532 55522
rect 14028 54180 14084 54190
rect 14028 53956 14084 54124
rect 14028 53862 14084 53900
rect 13916 53452 14084 53508
rect 13804 52612 13860 53228
rect 13916 52834 13972 52846
rect 13916 52782 13918 52834
rect 13970 52782 13972 52834
rect 13916 52722 13972 52782
rect 13916 52670 13918 52722
rect 13970 52670 13972 52722
rect 13916 52658 13972 52670
rect 13804 52546 13860 52556
rect 13804 52276 13860 52286
rect 14028 52276 14084 53452
rect 14364 52836 14420 52846
rect 14364 52742 14420 52780
rect 14476 52722 14532 55470
rect 14588 55074 14644 55086
rect 14588 55022 14590 55074
rect 14642 55022 14644 55074
rect 14588 54964 14644 55022
rect 14588 54898 14644 54908
rect 14588 54292 14644 54302
rect 14588 53730 14644 54236
rect 14588 53678 14590 53730
rect 14642 53678 14644 53730
rect 14588 53172 14644 53678
rect 14700 53732 14756 53742
rect 14700 53618 14756 53676
rect 14700 53566 14702 53618
rect 14754 53566 14756 53618
rect 14700 53554 14756 53566
rect 14812 53396 14868 56924
rect 15036 56642 15092 56654
rect 15036 56590 15038 56642
rect 15090 56590 15092 56642
rect 14924 55970 14980 55982
rect 14924 55918 14926 55970
rect 14978 55918 14980 55970
rect 14924 55522 14980 55918
rect 14924 55470 14926 55522
rect 14978 55470 14980 55522
rect 14924 55458 14980 55470
rect 15036 55468 15092 56590
rect 15260 56306 15316 57708
rect 15372 57540 15428 57550
rect 15372 57446 15428 57484
rect 15484 56980 15540 57708
rect 16044 57092 16100 58772
rect 16380 58660 16436 59724
rect 16604 59714 16660 59724
rect 17612 59778 17668 59790
rect 17612 59726 17614 59778
rect 17666 59726 17668 59778
rect 17612 59556 17668 59726
rect 17612 59490 17668 59500
rect 18060 59778 18116 59790
rect 18060 59726 18062 59778
rect 18114 59726 18116 59778
rect 18060 59556 18116 59726
rect 18732 59778 18788 59790
rect 18732 59726 18734 59778
rect 18786 59726 18788 59778
rect 18060 59490 18116 59500
rect 18508 59556 18564 59566
rect 17948 59444 18004 59454
rect 17948 59350 18004 59388
rect 18396 59332 18452 59342
rect 16604 59106 16660 59118
rect 16604 59054 16606 59106
rect 16658 59054 16660 59106
rect 16604 58996 16660 59054
rect 16604 58930 16660 58940
rect 17052 59106 17108 59118
rect 17052 59054 17054 59106
rect 17106 59054 17108 59106
rect 15484 56914 15540 56924
rect 15932 57036 16100 57092
rect 16156 58604 16436 58660
rect 16492 58884 16548 58894
rect 15932 56644 15988 57036
rect 16044 56868 16100 56878
rect 16044 56774 16100 56812
rect 15932 56588 16100 56644
rect 15260 56254 15262 56306
rect 15314 56254 15316 56306
rect 15260 56242 15316 56254
rect 15932 56308 15988 56318
rect 15036 55412 15204 55468
rect 15148 55280 15204 55356
rect 15820 55188 15876 55198
rect 15708 55076 15764 55086
rect 15708 54982 15764 55020
rect 15036 54626 15092 54638
rect 15036 54574 15038 54626
rect 15090 54574 15092 54626
rect 15036 53956 15092 54574
rect 15596 54514 15652 54526
rect 15596 54462 15598 54514
rect 15650 54462 15652 54514
rect 15596 54068 15652 54462
rect 15820 54180 15876 55132
rect 15596 54002 15652 54012
rect 15708 54124 15876 54180
rect 14924 53732 14980 53742
rect 15036 53732 15092 53900
rect 14924 53730 15092 53732
rect 14924 53678 14926 53730
rect 14978 53678 15092 53730
rect 14924 53676 15092 53678
rect 15708 53732 15764 54124
rect 15820 53956 15876 53966
rect 15820 53862 15876 53900
rect 15932 53954 15988 56252
rect 15932 53902 15934 53954
rect 15986 53902 15988 53954
rect 15932 53890 15988 53902
rect 16044 55970 16100 56588
rect 16156 56308 16212 58604
rect 16492 58548 16548 58828
rect 16940 58772 16996 58782
rect 16380 58492 16548 58548
rect 16604 58548 16660 58558
rect 16268 58436 16324 58446
rect 16268 57538 16324 58380
rect 16380 57874 16436 58492
rect 16604 58454 16660 58492
rect 16380 57822 16382 57874
rect 16434 57822 16436 57874
rect 16380 57810 16436 57822
rect 16492 58210 16548 58222
rect 16492 58158 16494 58210
rect 16546 58158 16548 58210
rect 16268 57486 16270 57538
rect 16322 57486 16324 57538
rect 16268 57474 16324 57486
rect 16492 57092 16548 58158
rect 16492 57026 16548 57036
rect 16604 57426 16660 57438
rect 16604 57374 16606 57426
rect 16658 57374 16660 57426
rect 16604 56980 16660 57374
rect 16716 56980 16772 56990
rect 16604 56978 16772 56980
rect 16604 56926 16718 56978
rect 16770 56926 16772 56978
rect 16604 56924 16772 56926
rect 16716 56914 16772 56924
rect 16492 56866 16548 56878
rect 16492 56814 16494 56866
rect 16546 56814 16548 56866
rect 16492 56756 16548 56814
rect 16492 56690 16548 56700
rect 16828 56756 16884 56766
rect 16492 56308 16548 56318
rect 16156 56306 16548 56308
rect 16156 56254 16494 56306
rect 16546 56254 16548 56306
rect 16156 56252 16548 56254
rect 16044 55918 16046 55970
rect 16098 55918 16100 55970
rect 15932 53732 15988 53742
rect 15708 53730 15988 53732
rect 15708 53678 15934 53730
rect 15986 53678 15988 53730
rect 15708 53676 15988 53678
rect 14924 53666 14980 53676
rect 14588 53106 14644 53116
rect 14700 53340 14868 53396
rect 14924 53508 14980 53518
rect 14476 52670 14478 52722
rect 14530 52670 14532 52722
rect 13804 52182 13860 52220
rect 13916 52220 14084 52276
rect 14252 52388 14308 52398
rect 14252 52274 14308 52332
rect 14252 52222 14254 52274
rect 14306 52222 14308 52274
rect 13916 51492 13972 52220
rect 14252 52210 14308 52222
rect 13692 51426 13748 51436
rect 13804 51436 13972 51492
rect 14028 52052 14084 52062
rect 13804 51268 13860 51436
rect 13580 51212 13860 51268
rect 13916 51266 13972 51278
rect 13916 51214 13918 51266
rect 13970 51214 13972 51266
rect 13580 49812 13636 51212
rect 13916 50706 13972 51214
rect 13916 50654 13918 50706
rect 13970 50654 13972 50706
rect 13916 50642 13972 50654
rect 14028 50596 14084 51996
rect 14476 51940 14532 52670
rect 14700 52052 14756 53340
rect 14812 52948 14868 52958
rect 14812 52854 14868 52892
rect 14924 52724 14980 53452
rect 15372 53508 15428 53518
rect 15372 53414 15428 53452
rect 14476 51874 14532 51884
rect 14588 51996 14756 52052
rect 14812 52052 14868 52062
rect 13804 50484 13860 50522
rect 14028 50464 14084 50540
rect 14140 51492 14196 51502
rect 14140 50820 14196 51436
rect 14252 51380 14308 51390
rect 14252 51286 14308 51324
rect 14588 51268 14644 51996
rect 14812 51958 14868 51996
rect 14924 52050 14980 52668
rect 15260 52836 15316 52846
rect 15148 52164 15204 52174
rect 15148 52070 15204 52108
rect 14924 51998 14926 52050
rect 14978 51998 14980 52050
rect 14924 51986 14980 51998
rect 14140 50594 14196 50764
rect 14364 51212 14644 51268
rect 14364 50596 14420 51212
rect 14700 50708 14756 50718
rect 14140 50542 14142 50594
rect 14194 50542 14196 50594
rect 14140 50530 14196 50542
rect 14252 50540 14420 50596
rect 14476 50594 14532 50606
rect 14476 50542 14478 50594
rect 14530 50542 14532 50594
rect 14252 50428 14308 50540
rect 14476 50428 14532 50542
rect 14700 50596 14756 50652
rect 14700 50594 14868 50596
rect 14700 50542 14702 50594
rect 14754 50542 14868 50594
rect 14700 50540 14868 50542
rect 14700 50530 14756 50540
rect 13804 50418 13860 50428
rect 14140 50372 14308 50428
rect 14364 50372 14532 50428
rect 13804 49812 13860 49822
rect 13580 49756 13804 49812
rect 13804 49718 13860 49756
rect 13916 49250 13972 49262
rect 13916 49198 13918 49250
rect 13970 49198 13972 49250
rect 13916 49140 13972 49198
rect 13468 45714 13524 45724
rect 13580 49138 13972 49140
rect 13580 49086 13918 49138
rect 13970 49086 13972 49138
rect 13580 49084 13972 49086
rect 13244 45602 13300 45612
rect 13132 44146 13188 44156
rect 13020 43810 13076 43820
rect 12572 43764 12628 43774
rect 13580 43764 13636 49084
rect 13916 49074 13972 49084
rect 14140 48692 14196 50372
rect 14252 50036 14308 50046
rect 14364 50036 14420 50372
rect 14252 50034 14420 50036
rect 14252 49982 14254 50034
rect 14306 49982 14420 50034
rect 14252 49980 14420 49982
rect 14700 50260 14756 50270
rect 14252 49970 14308 49980
rect 14476 49924 14532 49934
rect 14476 49250 14532 49868
rect 14476 49198 14478 49250
rect 14530 49198 14532 49250
rect 14476 49186 14532 49198
rect 14588 49586 14644 49598
rect 14588 49534 14590 49586
rect 14642 49534 14644 49586
rect 14364 49140 14420 49150
rect 14364 49046 14420 49084
rect 14588 49028 14644 49534
rect 14588 48962 14644 48972
rect 14140 48626 14196 48636
rect 14588 48804 14644 48814
rect 14588 48466 14644 48748
rect 14588 48414 14590 48466
rect 14642 48414 14644 48466
rect 14588 48402 14644 48414
rect 14140 48244 14196 48254
rect 14140 48150 14196 48188
rect 14364 48244 14420 48254
rect 14700 48244 14756 50204
rect 14812 50148 14868 50540
rect 14812 50082 14868 50092
rect 15148 50594 15204 50606
rect 15148 50542 15150 50594
rect 15202 50542 15204 50594
rect 14812 49700 14868 49710
rect 14812 49606 14868 49644
rect 14924 49252 14980 49262
rect 14924 49026 14980 49196
rect 14924 48974 14926 49026
rect 14978 48974 14980 49026
rect 14924 48916 14980 48974
rect 14924 48850 14980 48860
rect 15036 48802 15092 48814
rect 15036 48750 15038 48802
rect 15090 48750 15092 48802
rect 14924 48692 14980 48702
rect 15036 48692 15092 48750
rect 15148 48804 15204 50542
rect 15260 49700 15316 52780
rect 15372 52834 15428 52846
rect 15372 52782 15374 52834
rect 15426 52782 15428 52834
rect 15372 52500 15428 52782
rect 15372 52434 15428 52444
rect 15932 52500 15988 53676
rect 16044 53060 16100 55918
rect 16156 55074 16212 55086
rect 16156 55022 16158 55074
rect 16210 55022 16212 55074
rect 16156 53284 16212 55022
rect 16380 54180 16436 54190
rect 16380 53954 16436 54124
rect 16380 53902 16382 53954
rect 16434 53902 16436 53954
rect 16380 53890 16436 53902
rect 16156 53218 16212 53228
rect 16492 53060 16548 56252
rect 16604 55410 16660 55422
rect 16604 55358 16606 55410
rect 16658 55358 16660 55410
rect 16604 54626 16660 55358
rect 16716 55188 16772 55198
rect 16716 55094 16772 55132
rect 16828 54738 16884 56700
rect 16940 56308 16996 58716
rect 17052 57540 17108 59054
rect 18172 58660 18228 58670
rect 18172 58546 18228 58604
rect 18172 58494 18174 58546
rect 18226 58494 18228 58546
rect 18172 58482 18228 58494
rect 17500 58436 17556 58446
rect 17500 58342 17556 58380
rect 18060 58436 18116 58446
rect 18060 58342 18116 58380
rect 17052 57474 17108 57484
rect 17612 57540 17668 57550
rect 17500 56868 17556 56878
rect 17500 56774 17556 56812
rect 17276 56756 17332 56766
rect 17276 56662 17332 56700
rect 16940 56306 17108 56308
rect 16940 56254 16942 56306
rect 16994 56254 17108 56306
rect 16940 56252 17108 56254
rect 16940 56242 16996 56252
rect 16828 54686 16830 54738
rect 16882 54686 16884 54738
rect 16828 54674 16884 54686
rect 16940 55186 16996 55198
rect 16940 55134 16942 55186
rect 16994 55134 16996 55186
rect 16604 54574 16606 54626
rect 16658 54574 16660 54626
rect 16604 54562 16660 54574
rect 16940 54180 16996 55134
rect 16940 54114 16996 54124
rect 16604 53956 16660 53966
rect 16604 53862 16660 53900
rect 17052 53060 17108 56252
rect 17612 56196 17668 57484
rect 18172 57540 18228 57550
rect 18172 57446 18228 57484
rect 17724 57092 17780 57102
rect 17724 56998 17780 57036
rect 17836 56866 17892 56878
rect 17836 56814 17838 56866
rect 17890 56814 17892 56866
rect 17836 56308 17892 56814
rect 18396 56868 18452 59276
rect 18396 56802 18452 56812
rect 18060 56756 18116 56766
rect 18060 56642 18116 56700
rect 18060 56590 18062 56642
rect 18114 56590 18116 56642
rect 18060 56578 18116 56590
rect 17836 56242 17892 56252
rect 18508 56308 18564 59500
rect 18620 59108 18676 59118
rect 18620 59014 18676 59052
rect 18732 57764 18788 59726
rect 19180 59780 19236 59790
rect 19740 59780 19796 59790
rect 19180 59778 19460 59780
rect 19180 59726 19182 59778
rect 19234 59726 19460 59778
rect 19180 59724 19460 59726
rect 19180 59714 19236 59724
rect 19068 59220 19124 59230
rect 19068 59218 19348 59220
rect 19068 59166 19070 59218
rect 19122 59166 19348 59218
rect 19068 59164 19348 59166
rect 19068 59154 19124 59164
rect 19068 58546 19124 58558
rect 19068 58494 19070 58546
rect 19122 58494 19124 58546
rect 18620 57708 18788 57764
rect 18956 58324 19012 58334
rect 18620 57092 18676 57708
rect 18956 57650 19012 58268
rect 18956 57598 18958 57650
rect 19010 57598 19012 57650
rect 18956 57586 19012 57598
rect 18732 57538 18788 57550
rect 18732 57486 18734 57538
rect 18786 57486 18788 57538
rect 18732 57092 18788 57486
rect 18732 57036 19012 57092
rect 18620 57026 18676 57036
rect 18956 56754 19012 57036
rect 19068 56978 19124 58494
rect 19180 58434 19236 58446
rect 19180 58382 19182 58434
rect 19234 58382 19236 58434
rect 19180 58324 19236 58382
rect 19180 58258 19236 58268
rect 19292 57874 19348 59164
rect 19292 57822 19294 57874
rect 19346 57822 19348 57874
rect 19292 57652 19348 57822
rect 19292 57586 19348 57596
rect 19404 57316 19460 59724
rect 19628 59778 19796 59780
rect 19628 59726 19742 59778
rect 19794 59726 19796 59778
rect 19628 59724 19796 59726
rect 19516 59332 19572 59342
rect 19516 59238 19572 59276
rect 19404 57250 19460 57260
rect 19628 57316 19684 59724
rect 19740 59714 19796 59724
rect 20188 59778 20244 59790
rect 20188 59726 20190 59778
rect 20242 59726 20244 59778
rect 19836 59612 20100 59622
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 19836 59546 20100 59556
rect 20188 59444 20244 59726
rect 20636 59778 20692 59790
rect 21420 59780 21476 59790
rect 20636 59726 20638 59778
rect 20690 59726 20692 59778
rect 20636 59556 20692 59726
rect 21308 59778 21476 59780
rect 21308 59726 21422 59778
rect 21474 59726 21476 59778
rect 21308 59724 21476 59726
rect 20636 59500 21252 59556
rect 20188 59388 20692 59444
rect 20076 59332 20132 59342
rect 20076 59238 20132 59276
rect 20300 59218 20356 59230
rect 20300 59166 20302 59218
rect 20354 59166 20356 59218
rect 20076 59108 20132 59118
rect 19852 58324 19908 58334
rect 19852 58230 19908 58268
rect 20076 58212 20132 59052
rect 20188 59106 20244 59118
rect 20188 59054 20190 59106
rect 20242 59054 20244 59106
rect 20188 58436 20244 59054
rect 20300 58548 20356 59166
rect 20300 58482 20356 58492
rect 20524 59218 20580 59230
rect 20524 59166 20526 59218
rect 20578 59166 20580 59218
rect 20524 58436 20580 59166
rect 20188 58370 20244 58380
rect 20412 58380 20580 58436
rect 20076 58156 20244 58212
rect 19836 58044 20100 58054
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 19836 57978 20100 57988
rect 20188 57876 20244 58156
rect 20076 57820 20244 57876
rect 20412 57874 20468 58380
rect 20412 57822 20414 57874
rect 20466 57822 20468 57874
rect 19852 57652 19908 57662
rect 19852 57558 19908 57596
rect 20076 57650 20132 57820
rect 20412 57810 20468 57822
rect 20524 58210 20580 58222
rect 20524 58158 20526 58210
rect 20578 58158 20580 58210
rect 20076 57598 20078 57650
rect 20130 57598 20132 57650
rect 20076 57586 20132 57598
rect 19404 57092 19460 57102
rect 19068 56926 19070 56978
rect 19122 56926 19124 56978
rect 19068 56914 19124 56926
rect 19180 56980 19236 56990
rect 18956 56702 18958 56754
rect 19010 56702 19012 56754
rect 18620 56308 18676 56318
rect 18508 56306 18676 56308
rect 18508 56254 18622 56306
rect 18674 56254 18676 56306
rect 18508 56252 18676 56254
rect 17500 56140 17668 56196
rect 17388 55074 17444 55086
rect 17388 55022 17390 55074
rect 17442 55022 17444 55074
rect 17388 53844 17444 55022
rect 17388 53778 17444 53788
rect 17276 53732 17332 53742
rect 17164 53508 17220 53518
rect 17276 53508 17332 53676
rect 17164 53506 17332 53508
rect 17164 53454 17166 53506
rect 17218 53454 17332 53506
rect 17164 53452 17332 53454
rect 17164 53442 17220 53452
rect 16044 53004 16212 53060
rect 16492 53004 16772 53060
rect 16044 52836 16100 52846
rect 16044 52742 16100 52780
rect 15932 52434 15988 52444
rect 16044 52388 16100 52398
rect 15708 52162 15764 52174
rect 15708 52110 15710 52162
rect 15762 52110 15764 52162
rect 15260 49634 15316 49644
rect 15372 52052 15428 52062
rect 15260 49364 15316 49374
rect 15260 49028 15316 49308
rect 15260 48896 15316 48972
rect 15148 48738 15204 48748
rect 14980 48636 15092 48692
rect 14812 48244 14868 48254
rect 14700 48242 14868 48244
rect 14700 48190 14814 48242
rect 14866 48190 14868 48242
rect 14700 48188 14868 48190
rect 14364 48150 14420 48188
rect 14476 48130 14532 48142
rect 14476 48078 14478 48130
rect 14530 48078 14532 48130
rect 14364 47572 14420 47582
rect 13692 47236 13748 47246
rect 14364 47236 14420 47516
rect 14476 47460 14532 48078
rect 14476 47394 14532 47404
rect 14476 47236 14532 47246
rect 14364 47234 14532 47236
rect 14364 47182 14478 47234
rect 14530 47182 14532 47234
rect 14364 47180 14532 47182
rect 13692 47142 13748 47180
rect 14476 47124 14532 47180
rect 14812 47236 14868 48188
rect 14924 48020 14980 48636
rect 14924 47954 14980 47964
rect 15148 47572 15204 47582
rect 15148 47478 15204 47516
rect 14812 47170 14868 47180
rect 14476 47058 14532 47068
rect 14364 47012 14420 47022
rect 14140 46900 14196 46910
rect 13916 46676 13972 46686
rect 13916 46582 13972 46620
rect 14140 46340 14196 46844
rect 14252 46786 14308 46798
rect 14252 46734 14254 46786
rect 14306 46734 14308 46786
rect 14252 46676 14308 46734
rect 14364 46786 14420 46956
rect 14364 46734 14366 46786
rect 14418 46734 14420 46786
rect 14364 46722 14420 46734
rect 14252 46610 14308 46620
rect 15260 46676 15316 46686
rect 15260 46582 15316 46620
rect 14700 46562 14756 46574
rect 14700 46510 14702 46562
rect 14754 46510 14756 46562
rect 14140 46274 14196 46284
rect 14588 46340 14644 46350
rect 14252 46228 14308 46238
rect 14028 45892 14084 45902
rect 13916 45780 13972 45790
rect 13916 45686 13972 45724
rect 14028 45778 14084 45836
rect 14028 45726 14030 45778
rect 14082 45726 14084 45778
rect 14028 45444 14084 45726
rect 14028 45378 14084 45388
rect 14252 45666 14308 46172
rect 14252 45614 14254 45666
rect 14306 45614 14308 45666
rect 13804 44548 13860 44558
rect 13804 44434 13860 44492
rect 13804 44382 13806 44434
rect 13858 44382 13860 44434
rect 13804 44370 13860 44382
rect 12460 43762 12852 43764
rect 12460 43710 12574 43762
rect 12626 43710 12852 43762
rect 12460 43708 12852 43710
rect 12572 43698 12628 43708
rect 12348 43598 12350 43650
rect 12402 43598 12404 43650
rect 12348 43586 12404 43598
rect 12012 43540 12068 43550
rect 11900 43538 12068 43540
rect 11900 43486 12014 43538
rect 12066 43486 12068 43538
rect 11900 43484 12068 43486
rect 11900 43204 11956 43484
rect 12012 43474 12068 43484
rect 11900 43138 11956 43148
rect 12124 42980 12180 42990
rect 11788 42924 12068 42980
rect 11564 42642 11732 42644
rect 11564 42590 11566 42642
rect 11618 42590 11732 42642
rect 11564 42588 11732 42590
rect 11564 42420 11620 42588
rect 11676 42420 11732 42588
rect 11788 42754 11844 42766
rect 11788 42702 11790 42754
rect 11842 42702 11844 42754
rect 11788 42644 11844 42702
rect 11788 42578 11844 42588
rect 11676 42364 11844 42420
rect 11564 42354 11620 42364
rect 11452 42140 11620 42196
rect 11228 41970 11284 42028
rect 11228 41918 11230 41970
rect 11282 41918 11284 41970
rect 11228 41906 11284 41918
rect 11452 41972 11508 41982
rect 11116 41358 11118 41410
rect 11170 41358 11172 41410
rect 11116 41346 11172 41358
rect 11116 41188 11172 41198
rect 11116 40516 11172 41132
rect 11228 40964 11284 40974
rect 11228 40962 11396 40964
rect 11228 40910 11230 40962
rect 11282 40910 11396 40962
rect 11228 40908 11396 40910
rect 11228 40898 11284 40908
rect 11228 40516 11284 40526
rect 11116 40460 11228 40516
rect 11228 40384 11284 40460
rect 11116 40292 11172 40302
rect 11116 40198 11172 40236
rect 11340 40292 11396 40908
rect 11452 40514 11508 41916
rect 11564 41298 11620 42140
rect 11788 41300 11844 42364
rect 12012 41970 12068 42924
rect 12012 41918 12014 41970
rect 12066 41918 12068 41970
rect 12012 41410 12068 41918
rect 12124 41972 12180 42924
rect 12348 42868 12404 42878
rect 12348 42644 12404 42812
rect 12348 42578 12404 42588
rect 12796 41972 12852 43708
rect 13468 43652 13524 43662
rect 13580 43652 13636 43708
rect 13468 43650 13636 43652
rect 13468 43598 13470 43650
rect 13522 43598 13636 43650
rect 13468 43596 13636 43598
rect 13804 44100 13860 44110
rect 13468 43586 13524 43596
rect 12908 43540 12964 43550
rect 12908 43446 12964 43484
rect 13356 43540 13412 43550
rect 13020 43428 13076 43438
rect 13020 43334 13076 43372
rect 13356 42644 13412 43484
rect 13020 42530 13076 42542
rect 13020 42478 13022 42530
rect 13074 42478 13076 42530
rect 12908 41972 12964 41982
rect 12796 41970 12964 41972
rect 12796 41918 12910 41970
rect 12962 41918 12964 41970
rect 12796 41916 12964 41918
rect 12124 41906 12180 41916
rect 12572 41860 12628 41870
rect 12572 41858 12740 41860
rect 12572 41806 12574 41858
rect 12626 41806 12740 41858
rect 12572 41804 12740 41806
rect 12572 41794 12628 41804
rect 12012 41358 12014 41410
rect 12066 41358 12068 41410
rect 12012 41346 12068 41358
rect 12460 41636 12516 41646
rect 11564 41246 11566 41298
rect 11618 41246 11620 41298
rect 11564 40852 11620 41246
rect 11732 41244 11844 41300
rect 12460 41298 12516 41580
rect 12460 41246 12462 41298
rect 12514 41246 12516 41298
rect 11732 41076 11788 41244
rect 12460 41076 12516 41246
rect 11732 41020 11844 41076
rect 11564 40786 11620 40796
rect 11676 40628 11732 40638
rect 11676 40534 11732 40572
rect 11452 40462 11454 40514
rect 11506 40462 11508 40514
rect 11452 40450 11508 40462
rect 11340 40226 11396 40236
rect 11564 40404 11620 40414
rect 10892 39900 11060 39956
rect 10668 39566 10670 39618
rect 10722 39566 10724 39618
rect 10668 39554 10724 39566
rect 10780 39730 10836 39742
rect 10780 39678 10782 39730
rect 10834 39678 10836 39730
rect 10332 39340 10612 39396
rect 10220 39218 10276 39228
rect 9996 38882 10052 38892
rect 10444 39060 10500 39070
rect 10332 38836 10388 38846
rect 10220 38834 10388 38836
rect 10220 38782 10334 38834
rect 10386 38782 10388 38834
rect 10220 38780 10388 38782
rect 9772 38722 9828 38734
rect 9772 38670 9774 38722
rect 9826 38670 9828 38722
rect 9772 38668 9828 38670
rect 10108 38724 10164 38734
rect 9772 38612 9940 38668
rect 9772 37940 9828 37950
rect 9772 37846 9828 37884
rect 9772 37266 9828 37278
rect 9772 37214 9774 37266
rect 9826 37214 9828 37266
rect 9548 36978 9604 36988
rect 9660 37156 9716 37166
rect 9436 36764 9604 36820
rect 9436 36596 9492 36606
rect 9100 36428 9268 36484
rect 9324 36484 9380 36494
rect 8988 36148 9044 36158
rect 8988 35922 9044 36092
rect 8988 35870 8990 35922
rect 9042 35870 9044 35922
rect 8988 35858 9044 35870
rect 9100 34244 9156 36428
rect 9324 36390 9380 36428
rect 9436 36482 9492 36540
rect 9436 36430 9438 36482
rect 9490 36430 9492 36482
rect 9436 36418 9492 36430
rect 9212 36260 9268 36270
rect 9212 36258 9380 36260
rect 9212 36206 9214 36258
rect 9266 36206 9380 36258
rect 9212 36204 9380 36206
rect 9212 36194 9268 36204
rect 9324 36148 9380 36204
rect 9324 35476 9380 36092
rect 9324 35410 9380 35420
rect 9548 35700 9604 36764
rect 9100 34178 9156 34188
rect 9212 35364 9268 35374
rect 9212 34356 9268 35308
rect 8988 34018 9044 34030
rect 8988 33966 8990 34018
rect 9042 33966 9044 34018
rect 8988 33796 9044 33966
rect 8988 33730 9044 33740
rect 8876 33394 8932 33404
rect 9212 33124 9268 34300
rect 9212 33030 9268 33068
rect 9548 32788 9604 35644
rect 9660 35026 9716 37100
rect 9772 35252 9828 37214
rect 9884 36036 9940 38612
rect 10108 38274 10164 38668
rect 10108 38222 10110 38274
rect 10162 38222 10164 38274
rect 10108 38210 10164 38222
rect 10220 38052 10276 38780
rect 10332 38770 10388 38780
rect 10332 38276 10388 38286
rect 10332 38162 10388 38220
rect 10332 38110 10334 38162
rect 10386 38110 10388 38162
rect 10332 38098 10388 38110
rect 9996 37380 10052 37390
rect 9996 37286 10052 37324
rect 10220 37268 10276 37996
rect 10444 38052 10500 39004
rect 10444 37986 10500 37996
rect 10556 37716 10612 39340
rect 10668 38948 10724 38958
rect 10780 38948 10836 39678
rect 10892 38948 10948 38958
rect 10780 38946 10948 38948
rect 10780 38894 10894 38946
rect 10946 38894 10948 38946
rect 10780 38892 10948 38894
rect 10668 38834 10724 38892
rect 10892 38882 10948 38892
rect 10668 38782 10670 38834
rect 10722 38782 10724 38834
rect 10668 38770 10724 38782
rect 10780 38722 10836 38734
rect 10780 38670 10782 38722
rect 10834 38670 10836 38722
rect 10668 37828 10724 37838
rect 10668 37734 10724 37772
rect 10220 37202 10276 37212
rect 10332 37660 10612 37716
rect 10220 37044 10276 37054
rect 10220 36950 10276 36988
rect 9996 36932 10052 36942
rect 9996 36706 10052 36876
rect 9996 36654 9998 36706
rect 10050 36654 10052 36706
rect 9996 36642 10052 36654
rect 10108 36484 10164 36494
rect 10332 36484 10388 37660
rect 10556 37492 10612 37502
rect 10556 37398 10612 37436
rect 10668 37380 10724 37390
rect 10556 37266 10612 37278
rect 10556 37214 10558 37266
rect 10610 37214 10612 37266
rect 10556 37044 10612 37214
rect 10556 36978 10612 36988
rect 10668 36932 10724 37324
rect 10668 36596 10724 36876
rect 10108 36390 10164 36428
rect 10220 36428 10388 36484
rect 10556 36540 10724 36596
rect 9884 35970 9940 35980
rect 10108 35812 10164 35822
rect 10108 35698 10164 35756
rect 10108 35646 10110 35698
rect 10162 35646 10164 35698
rect 10108 35476 10164 35646
rect 10108 35410 10164 35420
rect 9772 35186 9828 35196
rect 9660 34974 9662 35026
rect 9714 34974 9716 35026
rect 9660 34962 9716 34974
rect 9884 35028 9940 35038
rect 9884 33570 9940 34972
rect 9884 33518 9886 33570
rect 9938 33518 9940 33570
rect 9884 33506 9940 33518
rect 9996 34244 10052 34254
rect 9548 32722 9604 32732
rect 9660 33348 9716 33358
rect 9100 32564 9156 32574
rect 9100 32470 9156 32508
rect 9212 32004 9268 32014
rect 9212 31666 9268 31948
rect 9212 31614 9214 31666
rect 9266 31614 9268 31666
rect 9212 31602 9268 31614
rect 9324 31778 9380 31790
rect 9324 31726 9326 31778
rect 9378 31726 9380 31778
rect 8540 30942 8542 30994
rect 8594 30942 8596 30994
rect 8540 30930 8596 30942
rect 8652 30994 8820 30996
rect 8652 30942 8766 30994
rect 8818 30942 8820 30994
rect 8652 30940 8820 30942
rect 8428 30322 8484 30380
rect 8428 30270 8430 30322
rect 8482 30270 8484 30322
rect 8428 30258 8484 30270
rect 8316 29314 8372 29326
rect 8316 29262 8318 29314
rect 8370 29262 8372 29314
rect 8316 29092 8372 29262
rect 8316 29026 8372 29036
rect 8540 29204 8596 29214
rect 8316 28642 8372 28654
rect 8316 28590 8318 28642
rect 8370 28590 8372 28642
rect 8316 27860 8372 28590
rect 8428 27860 8484 27870
rect 8316 27804 8428 27860
rect 8428 27728 8484 27804
rect 7756 26852 7924 26908
rect 7980 26852 8036 26862
rect 7532 26126 7534 26178
rect 7586 26126 7588 26178
rect 7532 26114 7588 26126
rect 7868 26850 8036 26852
rect 7868 26798 7982 26850
rect 8034 26798 8036 26850
rect 7868 26796 8036 26798
rect 7868 25844 7924 26796
rect 7980 26786 8036 26796
rect 8092 26852 8260 26908
rect 8316 27524 8372 27534
rect 8092 26628 8148 26852
rect 7868 25618 7924 25788
rect 7868 25566 7870 25618
rect 7922 25566 7924 25618
rect 7868 25508 7924 25566
rect 7868 25442 7924 25452
rect 7980 26572 8148 26628
rect 7420 25282 7476 25294
rect 7420 25230 7422 25282
rect 7474 25230 7476 25282
rect 7420 24836 7476 25230
rect 7420 24770 7476 24780
rect 7084 24670 7086 24722
rect 7138 24670 7140 24722
rect 7084 24276 7140 24670
rect 6524 24098 6580 24108
rect 6748 24220 7140 24276
rect 6748 23940 6804 24220
rect 7308 24164 7364 24174
rect 6300 23884 6580 23940
rect 5964 23378 6132 23380
rect 5964 23326 5966 23378
rect 6018 23326 6132 23378
rect 5964 23324 6132 23326
rect 5964 22482 6020 23324
rect 5964 22430 5966 22482
rect 6018 22430 6020 22482
rect 5852 21700 5908 21710
rect 5180 21532 5572 21588
rect 5740 21698 5908 21700
rect 5740 21646 5854 21698
rect 5906 21646 5908 21698
rect 5740 21644 5908 21646
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4844 21196 5012 21252
rect 5068 21476 5124 21486
rect 4508 21026 4564 21038
rect 4508 20974 4510 21026
rect 4562 20974 4564 21026
rect 4508 20914 4564 20974
rect 4508 20862 4510 20914
rect 4562 20862 4564 20914
rect 4508 20850 4564 20862
rect 4508 20356 4564 20366
rect 4844 20356 4900 21196
rect 4956 21028 5012 21038
rect 4956 20914 5012 20972
rect 4956 20862 4958 20914
rect 5010 20862 5012 20914
rect 4956 20850 5012 20862
rect 4564 20300 4900 20356
rect 4956 20356 5012 20366
rect 4508 20130 4564 20300
rect 4508 20078 4510 20130
rect 4562 20078 4564 20130
rect 4508 20066 4564 20078
rect 4956 20130 5012 20300
rect 4956 20078 4958 20130
rect 5010 20078 5012 20130
rect 4956 20066 5012 20078
rect 4060 18958 4062 19010
rect 4114 18958 4116 19010
rect 3388 18452 3444 18462
rect 3388 18358 3444 18396
rect 4060 18340 4116 18958
rect 4060 18274 4116 18284
rect 4172 18676 4228 18686
rect 4284 18676 4340 19964
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 5068 19348 5124 21420
rect 5180 19684 5236 21532
rect 5516 21028 5572 21038
rect 5180 19618 5236 19628
rect 5292 20242 5348 20254
rect 5292 20190 5294 20242
rect 5346 20190 5348 20242
rect 4956 19236 5012 19246
rect 5068 19216 5124 19292
rect 4228 18620 4340 18676
rect 4508 19010 4564 19022
rect 4508 18958 4510 19010
rect 4562 18958 4564 19010
rect 4508 18676 4564 18958
rect 2268 17714 2324 17724
rect 4060 17780 4116 17790
rect 4172 17780 4228 18620
rect 4508 18610 4564 18620
rect 4620 18340 4676 18350
rect 4620 18246 4676 18284
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4060 17778 4228 17780
rect 4060 17726 4062 17778
rect 4114 17726 4228 17778
rect 4060 17724 4228 17726
rect 4508 17780 4564 17790
rect 4060 17714 4116 17724
rect 4508 17686 4564 17724
rect 4844 17780 4900 17790
rect 4620 17108 4676 17118
rect 4620 17014 4676 17052
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4844 14644 4900 17724
rect 4956 17778 5012 19180
rect 4956 17726 4958 17778
rect 5010 17726 5012 17778
rect 4956 17714 5012 17726
rect 5068 18450 5124 18462
rect 5068 18398 5070 18450
rect 5122 18398 5124 18450
rect 5068 17108 5124 18398
rect 5292 17220 5348 20190
rect 5516 20188 5572 20972
rect 5628 20916 5684 20926
rect 5628 20822 5684 20860
rect 5516 20132 5684 20188
rect 5628 17780 5684 20132
rect 5740 18450 5796 21644
rect 5852 21634 5908 21644
rect 5964 21588 6020 22430
rect 6412 22260 6468 22270
rect 6412 22166 6468 22204
rect 6412 21812 6468 21822
rect 6188 21700 6244 21710
rect 6188 21606 6244 21644
rect 5964 20916 6020 21532
rect 6076 20916 6132 20926
rect 5964 20914 6132 20916
rect 5964 20862 6078 20914
rect 6130 20862 6132 20914
rect 5964 20860 6132 20862
rect 5852 20244 5908 20254
rect 6076 20244 6132 20860
rect 6412 20916 6468 21756
rect 5852 20242 6020 20244
rect 5852 20190 5854 20242
rect 5906 20190 6020 20242
rect 5852 20188 6020 20190
rect 5852 20178 5908 20188
rect 5852 19348 5908 19358
rect 5852 19254 5908 19292
rect 5740 18398 5742 18450
rect 5794 18398 5796 18450
rect 5740 18386 5796 18398
rect 5740 17780 5796 17790
rect 5628 17778 5796 17780
rect 5628 17726 5742 17778
rect 5794 17726 5796 17778
rect 5628 17724 5796 17726
rect 5740 17714 5796 17724
rect 5292 17164 5796 17220
rect 5068 17106 5460 17108
rect 5068 17054 5070 17106
rect 5122 17054 5460 17106
rect 5068 17052 5460 17054
rect 5068 17042 5124 17052
rect 5292 16884 5348 16894
rect 4956 14644 5012 14654
rect 4284 14642 5012 14644
rect 4284 14590 4958 14642
rect 5010 14590 5012 14642
rect 4284 14588 5012 14590
rect 4284 13746 4340 14588
rect 4284 13694 4286 13746
rect 4338 13694 4340 13746
rect 4284 13682 4340 13694
rect 3948 13634 4004 13646
rect 3948 13582 3950 13634
rect 4002 13582 4004 13634
rect 3836 12964 3892 12974
rect 3948 12964 4004 13582
rect 4284 13522 4340 13534
rect 4284 13470 4286 13522
rect 4338 13470 4340 13522
rect 4284 13076 4340 13470
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4844 13188 4900 14588
rect 4956 14578 5012 14588
rect 4284 13010 4340 13020
rect 4732 13132 5012 13188
rect 3836 12962 4004 12964
rect 3836 12910 3838 12962
rect 3890 12910 4004 12962
rect 3836 12908 4004 12910
rect 3836 12898 3892 12908
rect 3500 12852 3556 12862
rect 3500 12758 3556 12796
rect 4284 12852 4340 12862
rect 3612 12738 3668 12750
rect 3612 12686 3614 12738
rect 3666 12686 3668 12738
rect 3612 12180 3668 12686
rect 3612 12114 3668 12124
rect 4172 12180 4228 12190
rect 4172 12086 4228 12124
rect 4284 12066 4340 12796
rect 4732 12850 4788 13132
rect 4732 12798 4734 12850
rect 4786 12798 4788 12850
rect 4732 12786 4788 12798
rect 4956 12852 5012 13132
rect 4956 12796 5124 12852
rect 4508 12738 4564 12750
rect 4508 12686 4510 12738
rect 4562 12686 4564 12738
rect 4508 12180 4564 12686
rect 4844 12740 4900 12750
rect 4844 12738 5012 12740
rect 4844 12686 4846 12738
rect 4898 12686 5012 12738
rect 4844 12684 5012 12686
rect 4844 12674 4900 12684
rect 4508 12114 4564 12124
rect 4284 12014 4286 12066
rect 4338 12014 4340 12066
rect 4284 12002 4340 12014
rect 4620 12068 4676 12078
rect 4620 12066 4900 12068
rect 4620 12014 4622 12066
rect 4674 12014 4900 12066
rect 4620 12012 4900 12014
rect 4620 12002 4676 12012
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4844 11396 4900 12012
rect 4844 11330 4900 11340
rect 4844 10612 4900 10622
rect 4284 10610 4900 10612
rect 4284 10558 4846 10610
rect 4898 10558 4900 10610
rect 4284 10556 4900 10558
rect 4284 9826 4340 10556
rect 4844 10546 4900 10556
rect 4956 10500 5012 12684
rect 5068 11506 5124 12796
rect 5068 11454 5070 11506
rect 5122 11454 5124 11506
rect 5068 11172 5124 11454
rect 5068 11106 5124 11116
rect 5068 10500 5124 10510
rect 4956 10498 5124 10500
rect 4956 10446 5070 10498
rect 5122 10446 5124 10498
rect 4956 10444 5124 10446
rect 4956 10388 5012 10444
rect 5068 10434 5124 10444
rect 4844 10332 5012 10388
rect 5292 10386 5348 16828
rect 5404 16882 5460 17052
rect 5404 16830 5406 16882
rect 5458 16830 5460 16882
rect 5404 15426 5460 16830
rect 5404 15374 5406 15426
rect 5458 15374 5460 15426
rect 5404 14644 5460 15374
rect 5628 14644 5684 14654
rect 5404 14588 5628 14644
rect 5404 13746 5460 14588
rect 5628 14512 5684 14588
rect 5404 13694 5406 13746
rect 5458 13694 5460 13746
rect 5404 12964 5460 13694
rect 5740 13746 5796 17164
rect 5964 16882 6020 20188
rect 6076 20178 6132 20188
rect 6188 20692 6244 20702
rect 6188 20130 6244 20636
rect 6188 20078 6190 20130
rect 6242 20078 6244 20130
rect 6188 20066 6244 20078
rect 6300 19348 6356 19358
rect 6412 19348 6468 20860
rect 6300 19346 6468 19348
rect 6300 19294 6302 19346
rect 6354 19294 6468 19346
rect 6300 19292 6468 19294
rect 6524 19348 6580 23884
rect 6636 23938 6804 23940
rect 6636 23886 6750 23938
rect 6802 23886 6804 23938
rect 6636 23884 6804 23886
rect 6636 23156 6692 23884
rect 6748 23874 6804 23884
rect 7084 23940 7140 23950
rect 6636 21924 6692 23100
rect 6972 23604 7028 23614
rect 6972 23042 7028 23548
rect 6972 22990 6974 23042
rect 7026 22990 7028 23042
rect 6972 22978 7028 22990
rect 6636 21858 6692 21868
rect 6748 22484 6804 22494
rect 6636 21588 6692 21598
rect 6636 21494 6692 21532
rect 6636 20690 6692 20702
rect 6636 20638 6638 20690
rect 6690 20638 6692 20690
rect 6636 20356 6692 20638
rect 6636 20290 6692 20300
rect 6300 19282 6356 19292
rect 6524 19282 6580 19292
rect 6636 19684 6692 19694
rect 6636 19012 6692 19628
rect 6748 19346 6804 22428
rect 6860 22146 6916 22158
rect 6860 22094 6862 22146
rect 6914 22094 6916 22146
rect 6860 21812 6916 22094
rect 6860 21746 6916 21756
rect 6860 20804 6916 20814
rect 6860 20132 6916 20748
rect 7084 20188 7140 23884
rect 7308 21810 7364 24108
rect 7644 24164 7700 24174
rect 7644 24050 7700 24108
rect 7644 23998 7646 24050
rect 7698 23998 7700 24050
rect 7644 23986 7700 23998
rect 7868 23604 7924 23614
rect 7868 23380 7924 23548
rect 7868 22370 7924 23324
rect 7980 22932 8036 26572
rect 8092 24724 8148 24734
rect 8092 23154 8148 24668
rect 8316 23268 8372 27468
rect 8428 27188 8484 27198
rect 8540 27188 8596 29148
rect 8428 27186 8596 27188
rect 8428 27134 8430 27186
rect 8482 27134 8596 27186
rect 8428 27132 8596 27134
rect 8652 27300 8708 30940
rect 8764 30930 8820 30940
rect 8988 30996 9044 31006
rect 8988 30902 9044 30940
rect 9324 30996 9380 31726
rect 9660 31668 9716 33292
rect 9996 33346 10052 34188
rect 10108 34132 10164 34170
rect 10108 34066 10164 34076
rect 10108 33908 10164 33918
rect 10220 33908 10276 36428
rect 10444 36372 10500 36382
rect 10444 36258 10500 36316
rect 10444 36206 10446 36258
rect 10498 36206 10500 36258
rect 10332 35474 10388 35486
rect 10332 35422 10334 35474
rect 10386 35422 10388 35474
rect 10332 35364 10388 35422
rect 10332 35298 10388 35308
rect 10164 33852 10276 33908
rect 10332 34802 10388 34814
rect 10332 34750 10334 34802
rect 10386 34750 10388 34802
rect 10108 33814 10164 33852
rect 9996 33294 9998 33346
rect 10050 33294 10052 33346
rect 9996 33282 10052 33294
rect 9884 33124 9940 33134
rect 9660 31602 9716 31612
rect 9772 33122 9940 33124
rect 9772 33070 9886 33122
rect 9938 33070 9940 33122
rect 9772 33068 9940 33070
rect 8876 30882 8932 30894
rect 8876 30830 8878 30882
rect 8930 30830 8932 30882
rect 8876 30436 8932 30830
rect 8876 30370 8932 30380
rect 8876 30212 8932 30222
rect 8876 29540 8932 30156
rect 9324 30212 9380 30940
rect 9660 31332 9716 31342
rect 9660 30994 9716 31276
rect 9660 30942 9662 30994
rect 9714 30942 9716 30994
rect 9660 30930 9716 30942
rect 9772 30548 9828 33068
rect 9884 33058 9940 33068
rect 10220 32562 10276 32574
rect 10220 32510 10222 32562
rect 10274 32510 10276 32562
rect 9996 32450 10052 32462
rect 9996 32398 9998 32450
rect 10050 32398 10052 32450
rect 9772 30482 9828 30492
rect 9884 32004 9940 32014
rect 9772 30322 9828 30334
rect 9772 30270 9774 30322
rect 9826 30270 9828 30322
rect 9548 30212 9604 30222
rect 9324 30210 9604 30212
rect 9324 30158 9550 30210
rect 9602 30158 9604 30210
rect 9324 30156 9604 30158
rect 9212 30100 9268 30110
rect 9212 30006 9268 30044
rect 8876 29538 9044 29540
rect 8876 29486 8878 29538
rect 8930 29486 9044 29538
rect 8876 29484 9044 29486
rect 8876 29474 8932 29484
rect 8988 27972 9044 29484
rect 9324 28980 9380 30156
rect 9548 30146 9604 30156
rect 9772 29426 9828 30270
rect 9884 29650 9940 31948
rect 9996 31108 10052 32398
rect 10108 32338 10164 32350
rect 10108 32286 10110 32338
rect 10162 32286 10164 32338
rect 10108 31892 10164 32286
rect 10220 32004 10276 32510
rect 10220 31938 10276 31948
rect 10108 31826 10164 31836
rect 10332 31220 10388 34750
rect 10444 31444 10500 36206
rect 10556 35698 10612 36540
rect 10780 36484 10836 38670
rect 10892 38052 10948 38062
rect 10892 37044 10948 37996
rect 10892 36978 10948 36988
rect 11004 36708 11060 39900
rect 11564 39842 11620 40348
rect 11788 40180 11844 41020
rect 12460 41010 12516 41020
rect 12012 40962 12068 40974
rect 12012 40910 12014 40962
rect 12066 40910 12068 40962
rect 12012 40516 12068 40910
rect 12012 40402 12068 40460
rect 12012 40350 12014 40402
rect 12066 40350 12068 40402
rect 12012 40338 12068 40350
rect 12124 40404 12180 40414
rect 12180 40348 12292 40404
rect 12124 40310 12180 40348
rect 11788 40124 12068 40180
rect 11564 39790 11566 39842
rect 11618 39790 11620 39842
rect 11564 39778 11620 39790
rect 11676 40068 11732 40078
rect 11452 39508 11508 39518
rect 11452 39414 11508 39452
rect 11676 39508 11732 40012
rect 11788 39620 11844 39630
rect 12012 39620 12068 40124
rect 11788 39618 11956 39620
rect 11788 39566 11790 39618
rect 11842 39566 11956 39618
rect 11788 39564 11956 39566
rect 11788 39554 11844 39564
rect 11564 39396 11620 39406
rect 11228 38274 11284 38286
rect 11228 38222 11230 38274
rect 11282 38222 11284 38274
rect 11116 37828 11172 37866
rect 11116 37762 11172 37772
rect 11116 37604 11172 37614
rect 11116 37378 11172 37548
rect 11116 37326 11118 37378
rect 11170 37326 11172 37378
rect 11116 37314 11172 37326
rect 11228 37380 11284 38222
rect 11564 38162 11620 39340
rect 11676 38836 11732 39452
rect 11900 39508 11956 39564
rect 12012 39618 12180 39620
rect 12012 39566 12014 39618
rect 12066 39566 12180 39618
rect 12012 39564 12180 39566
rect 12012 39554 12068 39564
rect 11788 38836 11844 38846
rect 11676 38834 11844 38836
rect 11676 38782 11790 38834
rect 11842 38782 11844 38834
rect 11676 38780 11844 38782
rect 11788 38770 11844 38780
rect 11564 38110 11566 38162
rect 11618 38110 11620 38162
rect 11564 38098 11620 38110
rect 11676 38164 11732 38174
rect 11228 37378 11396 37380
rect 11228 37326 11230 37378
rect 11282 37326 11396 37378
rect 11228 37324 11396 37326
rect 11228 37314 11284 37324
rect 11228 37156 11284 37166
rect 11228 37042 11284 37100
rect 11228 36990 11230 37042
rect 11282 36990 11284 37042
rect 11228 36978 11284 36990
rect 11004 36652 11172 36708
rect 10892 36596 10948 36634
rect 10892 36530 10948 36540
rect 10780 36418 10836 36428
rect 10668 36370 10724 36382
rect 10668 36318 10670 36370
rect 10722 36318 10724 36370
rect 10668 35924 10724 36318
rect 10892 36370 10948 36382
rect 10892 36318 10894 36370
rect 10946 36318 10948 36370
rect 10892 36260 10948 36318
rect 10892 36194 10948 36204
rect 10892 35924 10948 35934
rect 10668 35922 10948 35924
rect 10668 35870 10894 35922
rect 10946 35870 10948 35922
rect 10668 35868 10948 35870
rect 10892 35858 10948 35868
rect 10556 35646 10558 35698
rect 10610 35646 10612 35698
rect 10556 35634 10612 35646
rect 10780 35700 10836 35710
rect 10780 35606 10836 35644
rect 11004 35698 11060 35710
rect 11004 35646 11006 35698
rect 11058 35646 11060 35698
rect 11004 35476 11060 35646
rect 10668 35420 11060 35476
rect 10444 31378 10500 31388
rect 10556 34914 10612 34926
rect 10556 34862 10558 34914
rect 10610 34862 10612 34914
rect 10556 34018 10612 34862
rect 10556 33966 10558 34018
rect 10610 33966 10612 34018
rect 10556 31556 10612 33966
rect 10220 31164 10388 31220
rect 10444 31220 10500 31230
rect 10220 31108 10276 31164
rect 9996 31042 10052 31052
rect 10108 31052 10276 31108
rect 10108 30996 10164 31052
rect 10108 30902 10164 30940
rect 10332 30996 10388 31006
rect 10332 30902 10388 30940
rect 9884 29598 9886 29650
rect 9938 29598 9940 29650
rect 9884 29586 9940 29598
rect 10220 30882 10276 30894
rect 10220 30830 10222 30882
rect 10274 30830 10276 30882
rect 9772 29374 9774 29426
rect 9826 29374 9828 29426
rect 9380 28924 9604 28980
rect 9324 28914 9380 28924
rect 8988 27878 9044 27916
rect 9100 28642 9156 28654
rect 9100 28590 9102 28642
rect 9154 28590 9156 28642
rect 9100 28420 9156 28590
rect 8428 27122 8484 27132
rect 8652 26908 8708 27244
rect 8876 27860 8932 27870
rect 8540 26852 8708 26908
rect 8764 27188 8820 27198
rect 8540 26786 8596 26796
rect 8652 26290 8708 26302
rect 8652 26238 8654 26290
rect 8706 26238 8708 26290
rect 8316 23202 8372 23212
rect 8540 26180 8596 26190
rect 8092 23102 8094 23154
rect 8146 23102 8148 23154
rect 8092 23090 8148 23102
rect 8540 23044 8596 26124
rect 8652 24164 8708 26238
rect 8764 25618 8820 27132
rect 8764 25566 8766 25618
rect 8818 25566 8820 25618
rect 8764 25554 8820 25566
rect 8876 24836 8932 27804
rect 8988 26850 9044 26862
rect 8988 26798 8990 26850
rect 9042 26798 9044 26850
rect 8988 25730 9044 26798
rect 8988 25678 8990 25730
rect 9042 25678 9044 25730
rect 8988 25666 9044 25678
rect 9100 25732 9156 28364
rect 9548 28642 9604 28924
rect 9548 28590 9550 28642
rect 9602 28590 9604 28642
rect 9436 27186 9492 27198
rect 9436 27134 9438 27186
rect 9490 27134 9492 27186
rect 9436 26852 9492 27134
rect 9436 26786 9492 26796
rect 9548 26628 9604 28590
rect 9660 28532 9716 28542
rect 9660 28438 9716 28476
rect 9772 28418 9828 29374
rect 9884 29428 9940 29438
rect 9884 29202 9940 29372
rect 9884 29150 9886 29202
rect 9938 29150 9940 29202
rect 9884 29138 9940 29150
rect 9996 29204 10052 29214
rect 9772 28366 9774 28418
rect 9826 28366 9828 28418
rect 9772 27972 9828 28366
rect 9996 28084 10052 29148
rect 10220 28980 10276 30830
rect 10444 30212 10500 31164
rect 10108 28924 10276 28980
rect 10332 30156 10500 30212
rect 10556 30996 10612 31500
rect 10108 28196 10164 28924
rect 10332 28868 10388 30156
rect 10444 29988 10500 29998
rect 10444 29894 10500 29932
rect 10108 28130 10164 28140
rect 10220 28866 10388 28868
rect 10220 28814 10334 28866
rect 10386 28814 10388 28866
rect 10220 28812 10388 28814
rect 9772 27858 9828 27916
rect 9772 27806 9774 27858
rect 9826 27806 9828 27858
rect 9772 27794 9828 27806
rect 9884 28028 10052 28084
rect 9884 27412 9940 28028
rect 10108 27972 10164 27982
rect 9996 27860 10052 27898
rect 9996 27794 10052 27804
rect 10108 27634 10164 27916
rect 10108 27582 10110 27634
rect 10162 27582 10164 27634
rect 10108 27570 10164 27582
rect 9884 27356 10164 27412
rect 9436 26572 9604 26628
rect 9996 27076 10052 27086
rect 9100 25666 9156 25676
rect 9212 26180 9268 26190
rect 9212 25618 9268 26124
rect 9212 25566 9214 25618
rect 9266 25566 9268 25618
rect 9212 25554 9268 25566
rect 8876 24742 8932 24780
rect 9324 25396 9380 25406
rect 8652 24108 8820 24164
rect 8652 23940 8708 23950
rect 8652 23846 8708 23884
rect 8764 23938 8820 24108
rect 8764 23886 8766 23938
rect 8818 23886 8820 23938
rect 8764 23604 8820 23886
rect 8764 23538 8820 23548
rect 8988 23716 9044 23726
rect 8988 23380 9044 23660
rect 8988 23266 9044 23324
rect 8988 23214 8990 23266
rect 9042 23214 9044 23266
rect 8988 23202 9044 23214
rect 8652 23044 8708 23054
rect 8540 23042 8708 23044
rect 8540 22990 8654 23042
rect 8706 22990 8708 23042
rect 8540 22988 8708 22990
rect 7980 22876 8148 22932
rect 7868 22318 7870 22370
rect 7922 22318 7924 22370
rect 7868 22306 7924 22318
rect 7308 21758 7310 21810
rect 7362 21758 7364 21810
rect 7308 21028 7364 21758
rect 7420 22258 7476 22270
rect 7420 22206 7422 22258
rect 7474 22206 7476 22258
rect 7420 21700 7476 22206
rect 7420 21634 7476 21644
rect 7980 21698 8036 21710
rect 7980 21646 7982 21698
rect 8034 21646 8036 21698
rect 7868 21588 7924 21598
rect 7308 20962 7364 20972
rect 7532 21586 7924 21588
rect 7532 21534 7870 21586
rect 7922 21534 7924 21586
rect 7532 21532 7924 21534
rect 7532 20914 7588 21532
rect 7532 20862 7534 20914
rect 7586 20862 7588 20914
rect 7532 20850 7588 20862
rect 7308 20804 7364 20814
rect 7308 20710 7364 20748
rect 6860 20066 6916 20076
rect 6972 20132 7140 20188
rect 7196 20244 7252 20254
rect 7868 20242 7924 21532
rect 7980 21140 8036 21646
rect 8092 21700 8148 22876
rect 8092 21634 8148 21644
rect 8204 22482 8260 22494
rect 8204 22430 8206 22482
rect 8258 22430 8260 22482
rect 8204 21364 8260 22430
rect 8204 21298 8260 21308
rect 8540 21474 8596 21486
rect 8540 21422 8542 21474
rect 8594 21422 8596 21474
rect 8540 21364 8596 21422
rect 8540 21298 8596 21308
rect 7980 20804 8036 21084
rect 7980 20738 8036 20748
rect 8428 21252 8484 21262
rect 8428 20580 8484 21196
rect 8428 20486 8484 20524
rect 7868 20190 7870 20242
rect 7922 20190 7924 20242
rect 7196 20132 7364 20188
rect 7868 20178 7924 20190
rect 6860 19908 6916 19918
rect 6972 19908 7028 20132
rect 7084 20020 7140 20030
rect 7084 19926 7140 19964
rect 7196 20018 7252 20030
rect 7196 19966 7198 20018
rect 7250 19966 7252 20018
rect 6860 19906 7028 19908
rect 6860 19854 6862 19906
rect 6914 19854 7028 19906
rect 6860 19852 7028 19854
rect 6860 19458 6916 19852
rect 7196 19796 7252 19966
rect 6860 19406 6862 19458
rect 6914 19406 6916 19458
rect 6860 19394 6916 19406
rect 6972 19740 7252 19796
rect 6748 19294 6750 19346
rect 6802 19294 6804 19346
rect 6748 19282 6804 19294
rect 6636 18946 6692 18956
rect 5964 16830 5966 16882
rect 6018 16830 6020 16882
rect 5964 16818 6020 16830
rect 6076 18676 6132 18686
rect 6076 17442 6132 18620
rect 6748 18340 6804 18350
rect 6524 17780 6580 17790
rect 6524 17686 6580 17724
rect 6076 17390 6078 17442
rect 6130 17390 6132 17442
rect 5740 13694 5742 13746
rect 5794 13694 5796 13746
rect 5740 13682 5796 13694
rect 5852 15876 5908 15886
rect 6076 15876 6132 17390
rect 6412 16212 6468 16222
rect 6412 16118 6468 16156
rect 5852 15874 6132 15876
rect 5852 15822 5854 15874
rect 5906 15822 6132 15874
rect 5852 15820 6132 15822
rect 6748 15874 6804 18284
rect 6972 16212 7028 19740
rect 7308 19684 7364 20132
rect 7084 19628 7364 19684
rect 7644 20018 7700 20030
rect 7644 19966 7646 20018
rect 7698 19966 7700 20018
rect 7084 19346 7140 19628
rect 7084 19294 7086 19346
rect 7138 19294 7140 19346
rect 7084 19282 7140 19294
rect 7420 19458 7476 19470
rect 7420 19406 7422 19458
rect 7474 19406 7476 19458
rect 7084 18564 7140 18574
rect 7084 17778 7140 18508
rect 7084 17726 7086 17778
rect 7138 17726 7140 17778
rect 7084 17714 7140 17726
rect 6972 16146 7028 16156
rect 7420 17442 7476 19406
rect 7532 19460 7588 19470
rect 7532 19346 7588 19404
rect 7532 19294 7534 19346
rect 7586 19294 7588 19346
rect 7532 19236 7588 19294
rect 7532 19170 7588 19180
rect 7420 17390 7422 17442
rect 7474 17390 7476 17442
rect 6748 15822 6750 15874
rect 6802 15822 6804 15874
rect 5740 13076 5796 13086
rect 5628 12964 5684 12974
rect 5404 12962 5684 12964
rect 5404 12910 5630 12962
rect 5682 12910 5684 12962
rect 5404 12908 5684 12910
rect 5628 12898 5684 12908
rect 5404 12180 5460 12190
rect 5404 12086 5460 12124
rect 5740 11394 5796 13020
rect 5740 11342 5742 11394
rect 5794 11342 5796 11394
rect 5740 11330 5796 11342
rect 5292 10334 5294 10386
rect 5346 10334 5348 10386
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4284 9774 4286 9826
rect 4338 9774 4340 9826
rect 4284 9268 4340 9774
rect 4844 9826 4900 10332
rect 4844 9774 4846 9826
rect 4898 9774 4900 9826
rect 4844 9762 4900 9774
rect 4956 9716 5012 9726
rect 4956 9622 5012 9660
rect 4396 9268 4452 9278
rect 4284 9266 4452 9268
rect 4284 9214 4398 9266
rect 4450 9214 4452 9266
rect 4284 9212 4452 9214
rect 4396 9202 4452 9212
rect 4844 9268 4900 9278
rect 4844 9174 4900 9212
rect 4284 9044 4340 9054
rect 4284 8950 4340 8988
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 5292 8428 5348 10334
rect 5740 9716 5796 9726
rect 5740 9622 5796 9660
rect 5180 8372 5348 8428
rect 5180 7362 5236 8372
rect 5292 8306 5348 8316
rect 5516 9042 5572 9054
rect 5516 8990 5518 9042
rect 5570 8990 5572 9042
rect 5180 7310 5182 7362
rect 5234 7310 5236 7362
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 5180 6692 5236 7310
rect 4956 6636 5236 6692
rect 4732 6578 4788 6590
rect 4732 6526 4734 6578
rect 4786 6526 4788 6578
rect 4732 6244 4788 6526
rect 4844 6580 4900 6590
rect 4844 6486 4900 6524
rect 4956 6244 5012 6636
rect 4732 6188 5012 6244
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4956 5012 5012 6188
rect 5068 6466 5124 6478
rect 5068 6414 5070 6466
rect 5122 6414 5124 6466
rect 5068 5236 5124 6414
rect 5516 6468 5572 8990
rect 5852 8428 5908 15820
rect 6748 15204 6804 15822
rect 6748 15138 6804 15148
rect 7196 15876 7252 15886
rect 7420 15876 7476 17390
rect 7532 17780 7588 17790
rect 7532 16212 7588 17724
rect 7644 17108 7700 19966
rect 8204 19906 8260 19918
rect 8204 19854 8206 19906
rect 8258 19854 8260 19906
rect 7980 19348 8036 19358
rect 7980 19254 8036 19292
rect 8204 19124 8260 19854
rect 8204 19058 8260 19068
rect 8428 19012 8484 19022
rect 8428 18918 8484 18956
rect 8652 18676 8708 22988
rect 9100 22148 9156 22158
rect 8428 18620 8708 18676
rect 8764 22146 9156 22148
rect 8764 22094 9102 22146
rect 9154 22094 9156 22146
rect 8764 22092 9156 22094
rect 7980 18562 8036 18574
rect 7980 18510 7982 18562
rect 8034 18510 8036 18562
rect 7980 18452 8036 18510
rect 7980 18386 8036 18396
rect 7868 17780 7924 17790
rect 7868 17686 7924 17724
rect 8428 17780 8484 18620
rect 8428 17648 8484 17724
rect 8540 18452 8596 18462
rect 7644 17042 7700 17052
rect 8540 17106 8596 18396
rect 8764 18450 8820 22092
rect 9100 22082 9156 22092
rect 8988 21812 9044 21822
rect 8988 21476 9044 21756
rect 8988 21410 9044 21420
rect 9100 21700 9156 21710
rect 8764 18398 8766 18450
rect 8818 18398 8820 18450
rect 8764 18386 8820 18398
rect 8876 20804 8932 20814
rect 8876 17220 8932 20748
rect 8988 20692 9044 20702
rect 8988 20598 9044 20636
rect 9100 20188 9156 21644
rect 8988 20132 9156 20188
rect 8988 19906 9044 20132
rect 8988 19854 8990 19906
rect 9042 19854 9044 19906
rect 8988 19346 9044 19854
rect 8988 19294 8990 19346
rect 9042 19294 9044 19346
rect 8988 19282 9044 19294
rect 8988 17444 9044 17454
rect 9324 17444 9380 25340
rect 9436 21700 9492 26572
rect 9660 26404 9716 26414
rect 9548 25730 9604 25742
rect 9548 25678 9550 25730
rect 9602 25678 9604 25730
rect 9548 23380 9604 25678
rect 9660 25620 9716 26348
rect 9660 25488 9716 25564
rect 9772 26292 9828 26302
rect 9772 26178 9828 26236
rect 9772 26126 9774 26178
rect 9826 26126 9828 26178
rect 9772 24052 9828 26126
rect 9996 25396 10052 27020
rect 10108 25844 10164 27356
rect 10220 26068 10276 28812
rect 10332 28802 10388 28812
rect 10444 29652 10500 29662
rect 10444 28308 10500 29596
rect 10332 27636 10388 27646
rect 10332 27188 10388 27580
rect 10332 27056 10388 27132
rect 10332 26516 10388 26526
rect 10332 26422 10388 26460
rect 10220 26002 10276 26012
rect 10444 25956 10500 28252
rect 10556 26964 10612 30940
rect 10668 34692 10724 35420
rect 11004 35252 11060 35262
rect 11004 34916 11060 35196
rect 11004 34822 11060 34860
rect 10668 34020 10724 34636
rect 11116 34690 11172 36652
rect 11116 34638 11118 34690
rect 11170 34638 11172 34690
rect 11116 34626 11172 34638
rect 11340 34356 11396 37324
rect 11564 36820 11620 36830
rect 11452 36484 11508 36494
rect 11452 35924 11508 36428
rect 11564 36482 11620 36764
rect 11564 36430 11566 36482
rect 11618 36430 11620 36482
rect 11564 36418 11620 36430
rect 11452 35868 11620 35924
rect 11340 34290 11396 34300
rect 10780 34132 10836 34142
rect 10780 34038 10836 34076
rect 10668 30212 10724 33964
rect 10780 33684 10836 33694
rect 10780 33570 10836 33628
rect 10780 33518 10782 33570
rect 10834 33518 10836 33570
rect 10780 33506 10836 33518
rect 11452 32676 11508 32686
rect 11228 32562 11284 32574
rect 11228 32510 11230 32562
rect 11282 32510 11284 32562
rect 11228 32452 11284 32510
rect 10780 31780 10836 31790
rect 10780 30994 10836 31724
rect 10780 30942 10782 30994
rect 10834 30942 10836 30994
rect 10780 30930 10836 30942
rect 11116 31778 11172 31790
rect 11116 31726 11118 31778
rect 11170 31726 11172 31778
rect 11004 30882 11060 30894
rect 11004 30830 11006 30882
rect 11058 30830 11060 30882
rect 11004 30660 11060 30830
rect 11004 30594 11060 30604
rect 11116 30548 11172 31726
rect 11228 31220 11284 32396
rect 11452 31668 11508 32620
rect 11228 31154 11284 31164
rect 11340 31666 11508 31668
rect 11340 31614 11454 31666
rect 11506 31614 11508 31666
rect 11340 31612 11508 31614
rect 11228 30994 11284 31006
rect 11228 30942 11230 30994
rect 11282 30942 11284 30994
rect 11228 30884 11284 30942
rect 11228 30818 11284 30828
rect 11116 30482 11172 30492
rect 11340 30436 11396 31612
rect 11452 31602 11508 31612
rect 11228 30380 11396 30436
rect 11452 30994 11508 31006
rect 11452 30942 11454 30994
rect 11506 30942 11508 30994
rect 11116 30324 11172 30334
rect 10668 30146 10724 30156
rect 11004 30212 11060 30222
rect 11004 30118 11060 30156
rect 11116 30210 11172 30268
rect 11116 30158 11118 30210
rect 11170 30158 11172 30210
rect 11116 29652 11172 30158
rect 11228 29988 11284 30380
rect 11228 29922 11284 29932
rect 11340 30212 11396 30222
rect 11116 29586 11172 29596
rect 11340 29650 11396 30156
rect 11340 29598 11342 29650
rect 11394 29598 11396 29650
rect 11340 29586 11396 29598
rect 11452 29986 11508 30942
rect 11452 29934 11454 29986
rect 11506 29934 11508 29986
rect 11452 29652 11508 29934
rect 10780 29540 10836 29550
rect 10780 29446 10836 29484
rect 11340 29428 11396 29438
rect 11116 29426 11396 29428
rect 11116 29374 11342 29426
rect 11394 29374 11396 29426
rect 11116 29372 11396 29374
rect 11004 29316 11060 29326
rect 11004 29222 11060 29260
rect 10892 28756 10948 28766
rect 11116 28756 11172 29372
rect 11340 29362 11396 29372
rect 11228 29204 11284 29214
rect 11228 29110 11284 29148
rect 10892 28754 11172 28756
rect 10892 28702 10894 28754
rect 10946 28702 11172 28754
rect 10892 28700 11172 28702
rect 10892 28690 10948 28700
rect 10668 28642 10724 28654
rect 10668 28590 10670 28642
rect 10722 28590 10724 28642
rect 10668 28532 10724 28590
rect 10668 28466 10724 28476
rect 10780 28420 10836 28430
rect 10780 28326 10836 28364
rect 11004 28418 11060 28430
rect 11004 28366 11006 28418
rect 11058 28366 11060 28418
rect 11004 27972 11060 28366
rect 11060 27916 11172 27972
rect 11004 27906 11060 27916
rect 10556 26898 10612 26908
rect 10892 26964 10948 27002
rect 10892 26898 10948 26908
rect 11004 26850 11060 26862
rect 11004 26798 11006 26850
rect 11058 26798 11060 26850
rect 11004 26516 11060 26798
rect 10444 25890 10500 25900
rect 10556 26460 11060 26516
rect 10108 25788 10276 25844
rect 9996 25330 10052 25340
rect 10108 25506 10164 25518
rect 10108 25454 10110 25506
rect 10162 25454 10164 25506
rect 9884 24948 9940 24958
rect 10108 24948 10164 25454
rect 10220 25172 10276 25788
rect 10556 25506 10612 26460
rect 10556 25454 10558 25506
rect 10610 25454 10612 25506
rect 10556 25442 10612 25454
rect 10668 26290 10724 26302
rect 10668 26238 10670 26290
rect 10722 26238 10724 26290
rect 10668 26068 10724 26238
rect 11004 26292 11060 26302
rect 11004 26198 11060 26236
rect 10444 25284 10500 25294
rect 10444 25190 10500 25228
rect 10220 25106 10276 25116
rect 9884 24946 10164 24948
rect 9884 24894 9886 24946
rect 9938 24894 10164 24946
rect 9884 24892 10164 24894
rect 9884 24882 9940 24892
rect 10444 24836 10500 24846
rect 10444 24742 10500 24780
rect 9996 24724 10052 24734
rect 9772 23986 9828 23996
rect 9884 24164 9940 24174
rect 9660 23380 9716 23390
rect 9548 23378 9716 23380
rect 9548 23326 9662 23378
rect 9714 23326 9716 23378
rect 9548 23324 9716 23326
rect 9548 23156 9604 23166
rect 9548 22482 9604 23100
rect 9548 22430 9550 22482
rect 9602 22430 9604 22482
rect 9548 22418 9604 22430
rect 9660 21812 9716 23324
rect 9884 22372 9940 24108
rect 9660 21746 9716 21756
rect 9772 22316 9940 22372
rect 9436 21634 9492 21644
rect 9772 21588 9828 22316
rect 9660 21532 9828 21588
rect 9884 22148 9940 22158
rect 9436 20804 9492 20814
rect 9436 20710 9492 20748
rect 9548 19012 9604 19022
rect 8988 17442 9380 17444
rect 8988 17390 8990 17442
rect 9042 17390 9380 17442
rect 8988 17388 9380 17390
rect 9436 19010 9604 19012
rect 9436 18958 9550 19010
rect 9602 18958 9604 19010
rect 9436 18956 9604 18958
rect 8988 17378 9044 17388
rect 8876 17164 9156 17220
rect 8540 17054 8542 17106
rect 8594 17054 8596 17106
rect 7756 16884 7812 16894
rect 7644 16212 7700 16222
rect 7532 16210 7700 16212
rect 7532 16158 7646 16210
rect 7698 16158 7700 16210
rect 7532 16156 7700 16158
rect 7644 16146 7700 16156
rect 7196 15874 7476 15876
rect 7196 15822 7198 15874
rect 7250 15822 7476 15874
rect 7196 15820 7476 15822
rect 7196 14754 7252 15820
rect 7196 14702 7198 14754
rect 7250 14702 7252 14754
rect 7196 14690 7252 14702
rect 7308 15316 7364 15326
rect 6412 14644 6468 14654
rect 6412 14550 6468 14588
rect 6860 14644 6916 14654
rect 6860 14550 6916 14588
rect 7308 14642 7364 15260
rect 7308 14590 7310 14642
rect 7362 14590 7364 14642
rect 7308 14578 7364 14590
rect 7756 14644 7812 16828
rect 8540 16884 8596 17054
rect 9100 17106 9156 17164
rect 9100 17054 9102 17106
rect 9154 17054 9156 17106
rect 9100 17042 9156 17054
rect 8540 16818 8596 16828
rect 8092 16098 8148 16110
rect 8092 16046 8094 16098
rect 8146 16046 8148 16098
rect 8092 14644 8148 16046
rect 8764 16100 8820 16110
rect 9436 16100 9492 18956
rect 9548 18946 9604 18956
rect 9660 18452 9716 21532
rect 9772 20916 9828 20926
rect 9772 20822 9828 20860
rect 9884 20188 9940 22092
rect 9996 21810 10052 24668
rect 10220 24498 10276 24510
rect 10220 24446 10222 24498
rect 10274 24446 10276 24498
rect 10220 24388 10276 24446
rect 10220 24322 10276 24332
rect 10556 24164 10612 24174
rect 10556 23828 10612 24108
rect 10556 23734 10612 23772
rect 9996 21758 9998 21810
rect 10050 21758 10052 21810
rect 9996 21746 10052 21758
rect 10108 23044 10164 23054
rect 10668 23044 10724 26012
rect 10892 25956 10948 25966
rect 10780 25394 10836 25406
rect 10780 25342 10782 25394
rect 10834 25342 10836 25394
rect 10780 25172 10836 25342
rect 10780 23716 10836 25116
rect 10780 23650 10836 23660
rect 10892 23604 10948 25900
rect 11116 25060 11172 27916
rect 11228 27074 11284 27086
rect 11228 27022 11230 27074
rect 11282 27022 11284 27074
rect 11228 26852 11284 27022
rect 11228 26786 11284 26796
rect 11452 27074 11508 29596
rect 11452 27022 11454 27074
rect 11506 27022 11508 27074
rect 11452 26404 11508 27022
rect 11564 26740 11620 35868
rect 11676 34580 11732 38108
rect 11900 37828 11956 39452
rect 12012 39284 12068 39294
rect 12012 38834 12068 39228
rect 12124 39172 12180 39564
rect 12236 39396 12292 40348
rect 12572 40290 12628 40302
rect 12572 40238 12574 40290
rect 12626 40238 12628 40290
rect 12460 39508 12516 39518
rect 12460 39414 12516 39452
rect 12236 39330 12292 39340
rect 12572 39284 12628 40238
rect 12684 39956 12740 41804
rect 12684 39890 12740 39900
rect 12796 41410 12852 41422
rect 12796 41358 12798 41410
rect 12850 41358 12852 41410
rect 12796 39732 12852 41358
rect 12908 41300 12964 41916
rect 13020 41972 13076 42478
rect 13244 42196 13300 42206
rect 13244 41972 13300 42140
rect 13356 42194 13412 42588
rect 13580 43428 13636 43438
rect 13356 42142 13358 42194
rect 13410 42142 13412 42194
rect 13356 42130 13412 42142
rect 13468 42196 13524 42206
rect 13468 42102 13524 42140
rect 13580 42194 13636 43372
rect 13580 42142 13582 42194
rect 13634 42142 13636 42194
rect 13580 42130 13636 42142
rect 13692 42642 13748 42654
rect 13692 42590 13694 42642
rect 13746 42590 13748 42642
rect 13692 42084 13748 42590
rect 13692 42018 13748 42028
rect 13244 41916 13524 41972
rect 13020 41906 13076 41916
rect 12908 41234 12964 41244
rect 13020 41524 13076 41534
rect 12908 41076 12964 41086
rect 13020 41076 13076 41468
rect 12908 41074 13076 41076
rect 12908 41022 12910 41074
rect 12962 41022 13076 41074
rect 12908 41020 13076 41022
rect 13356 41300 13412 41310
rect 12908 41010 12964 41020
rect 13020 40852 13076 40862
rect 13020 40516 13076 40796
rect 13020 40422 13076 40460
rect 12908 39732 12964 39742
rect 12796 39676 12908 39732
rect 12572 39218 12628 39228
rect 12124 39116 12292 39172
rect 12012 38782 12014 38834
rect 12066 38782 12068 38834
rect 12012 38770 12068 38782
rect 12124 38052 12180 38062
rect 11900 37156 11956 37772
rect 12012 37826 12068 37838
rect 12012 37774 12014 37826
rect 12066 37774 12068 37826
rect 12012 37380 12068 37774
rect 12124 37604 12180 37996
rect 12124 37490 12180 37548
rect 12124 37438 12126 37490
rect 12178 37438 12180 37490
rect 12124 37426 12180 37438
rect 12012 37314 12068 37324
rect 12124 37268 12180 37278
rect 11900 37100 12068 37156
rect 11676 34514 11732 34524
rect 11788 35922 11844 35934
rect 11788 35870 11790 35922
rect 11842 35870 11844 35922
rect 11788 35700 11844 35870
rect 11788 34244 11844 35644
rect 11900 35698 11956 35710
rect 11900 35646 11902 35698
rect 11954 35646 11956 35698
rect 11900 35252 11956 35646
rect 11900 35186 11956 35196
rect 12012 35140 12068 37100
rect 12124 37044 12180 37212
rect 12124 36594 12180 36988
rect 12124 36542 12126 36594
rect 12178 36542 12180 36594
rect 12124 36530 12180 36542
rect 12012 35074 12068 35084
rect 12124 35028 12180 35038
rect 12124 34934 12180 34972
rect 11900 34914 11956 34926
rect 11900 34862 11902 34914
rect 11954 34862 11956 34914
rect 11900 34580 11956 34862
rect 12236 34692 12292 39116
rect 12460 39060 12516 39070
rect 12460 38966 12516 39004
rect 12348 38836 12404 38846
rect 12348 38742 12404 38780
rect 12684 38834 12740 38846
rect 12684 38782 12686 38834
rect 12738 38782 12740 38834
rect 12572 38722 12628 38734
rect 12572 38670 12574 38722
rect 12626 38670 12628 38722
rect 12572 38164 12628 38670
rect 12684 38724 12740 38782
rect 12684 38658 12740 38668
rect 12908 38276 12964 39676
rect 13244 39284 13300 39294
rect 13244 39060 13300 39228
rect 12908 38210 12964 38220
rect 13020 39058 13300 39060
rect 13020 39006 13246 39058
rect 13298 39006 13300 39058
rect 13020 39004 13300 39006
rect 12572 38098 12628 38108
rect 12572 37826 12628 37838
rect 12572 37774 12574 37826
rect 12626 37774 12628 37826
rect 12572 37716 12628 37774
rect 12572 37156 12628 37660
rect 12908 37826 12964 37838
rect 12908 37774 12910 37826
rect 12962 37774 12964 37826
rect 12796 37604 12852 37614
rect 12684 37268 12740 37278
rect 12684 37174 12740 37212
rect 12796 37266 12852 37548
rect 12796 37214 12798 37266
rect 12850 37214 12852 37266
rect 12796 37202 12852 37214
rect 12572 37090 12628 37100
rect 12796 36708 12852 36718
rect 12796 36260 12852 36652
rect 12908 36484 12964 37774
rect 12908 36418 12964 36428
rect 12908 36260 12964 36270
rect 12796 36258 12964 36260
rect 12796 36206 12910 36258
rect 12962 36206 12964 36258
rect 12796 36204 12964 36206
rect 12684 36148 12740 36158
rect 12348 35700 12404 35738
rect 12348 35634 12404 35644
rect 12348 34692 12404 34702
rect 12236 34690 12404 34692
rect 12236 34638 12350 34690
rect 12402 34638 12404 34690
rect 12236 34636 12404 34638
rect 11900 34514 11956 34524
rect 11900 34356 11956 34366
rect 11900 34262 11956 34300
rect 12236 34356 12292 34366
rect 12236 34262 12292 34300
rect 11788 34178 11844 34188
rect 12348 33684 12404 34636
rect 12348 33618 12404 33628
rect 12460 34690 12516 34702
rect 12460 34638 12462 34690
rect 12514 34638 12516 34690
rect 12460 33348 12516 34638
rect 12572 34692 12628 34702
rect 12572 34598 12628 34636
rect 12684 33796 12740 36092
rect 12908 36148 12964 36204
rect 12908 36082 12964 36092
rect 13020 35922 13076 39004
rect 13244 38994 13300 39004
rect 13356 38668 13412 41244
rect 13020 35870 13022 35922
rect 13074 35870 13076 35922
rect 13020 35858 13076 35870
rect 13132 38612 13412 38668
rect 13468 40404 13524 41916
rect 13692 41076 13748 41086
rect 13692 40626 13748 41020
rect 13692 40574 13694 40626
rect 13746 40574 13748 40626
rect 13580 40404 13636 40414
rect 13468 40402 13636 40404
rect 13468 40350 13582 40402
rect 13634 40350 13636 40402
rect 13468 40348 13636 40350
rect 13468 38668 13524 40348
rect 13580 40338 13636 40348
rect 13692 40404 13748 40574
rect 13692 40338 13748 40348
rect 13692 39620 13748 39630
rect 13580 39396 13636 39406
rect 13580 39302 13636 39340
rect 13692 39058 13748 39564
rect 13692 39006 13694 39058
rect 13746 39006 13748 39058
rect 13468 38612 13636 38668
rect 13132 37378 13188 38612
rect 13580 37604 13636 38612
rect 13580 37538 13636 37548
rect 13132 37326 13134 37378
rect 13186 37326 13188 37378
rect 13132 35028 13188 37326
rect 13692 37380 13748 39006
rect 13804 37604 13860 44044
rect 14252 43540 14308 45614
rect 14476 45780 14532 45790
rect 14476 45106 14532 45724
rect 14476 45054 14478 45106
rect 14530 45054 14532 45106
rect 14364 44660 14420 44670
rect 14364 44322 14420 44604
rect 14364 44270 14366 44322
rect 14418 44270 14420 44322
rect 14364 44100 14420 44270
rect 14364 44034 14420 44044
rect 14252 43474 14308 43484
rect 14364 43538 14420 43550
rect 14364 43486 14366 43538
rect 14418 43486 14420 43538
rect 13916 43428 13972 43438
rect 13916 43334 13972 43372
rect 13916 42868 13972 42878
rect 13916 42754 13972 42812
rect 14252 42868 14308 42878
rect 14252 42774 14308 42812
rect 13916 42702 13918 42754
rect 13970 42702 13972 42754
rect 13916 42690 13972 42702
rect 14364 42756 14420 43486
rect 14364 42662 14420 42700
rect 14140 42644 14196 42654
rect 14140 42550 14196 42588
rect 14140 42196 14196 42206
rect 14140 41970 14196 42140
rect 14140 41918 14142 41970
rect 14194 41918 14196 41970
rect 14140 41906 14196 41918
rect 14364 41860 14420 41870
rect 14364 41766 14420 41804
rect 14476 41524 14532 45054
rect 14588 44324 14644 46284
rect 14700 45890 14756 46510
rect 15260 46004 15316 46014
rect 14700 45838 14702 45890
rect 14754 45838 14756 45890
rect 14700 45826 14756 45838
rect 14924 46002 15316 46004
rect 14924 45950 15262 46002
rect 15314 45950 15316 46002
rect 14924 45948 15316 45950
rect 14812 45218 14868 45230
rect 14812 45166 14814 45218
rect 14866 45166 14868 45218
rect 14812 45108 14868 45166
rect 14812 45042 14868 45052
rect 14924 44434 14980 45948
rect 15260 45938 15316 45948
rect 14924 44382 14926 44434
rect 14978 44382 14980 44434
rect 14924 44370 14980 44382
rect 15372 45890 15428 51996
rect 15708 51602 15764 52110
rect 15932 52164 15988 52174
rect 15708 51550 15710 51602
rect 15762 51550 15764 51602
rect 15708 51538 15764 51550
rect 15820 51604 15876 51614
rect 15596 51380 15652 51390
rect 15484 51378 15652 51380
rect 15484 51326 15598 51378
rect 15650 51326 15652 51378
rect 15484 51324 15652 51326
rect 15484 50370 15540 51324
rect 15596 51314 15652 51324
rect 15820 50820 15876 51548
rect 15932 51378 15988 52108
rect 15932 51326 15934 51378
rect 15986 51326 15988 51378
rect 15932 51314 15988 51326
rect 16044 52162 16100 52332
rect 16044 52110 16046 52162
rect 16098 52110 16100 52162
rect 16044 51380 16100 52110
rect 16044 51314 16100 51324
rect 15820 50754 15876 50764
rect 15484 50318 15486 50370
rect 15538 50318 15540 50370
rect 15484 50306 15540 50318
rect 15596 50484 15652 50494
rect 15596 50260 15652 50428
rect 15596 50194 15652 50204
rect 15820 50482 15876 50494
rect 15820 50430 15822 50482
rect 15874 50430 15876 50482
rect 15708 50036 15764 50046
rect 15708 49942 15764 49980
rect 15820 49698 15876 50430
rect 16156 50260 16212 53004
rect 16492 52834 16548 52846
rect 16492 52782 16494 52834
rect 16546 52782 16548 52834
rect 16492 52724 16548 52782
rect 16492 52658 16548 52668
rect 16268 51154 16324 51166
rect 16268 51102 16270 51154
rect 16322 51102 16324 51154
rect 16268 50820 16324 51102
rect 16492 51044 16548 51054
rect 16380 50820 16436 50830
rect 16268 50818 16436 50820
rect 16268 50766 16382 50818
rect 16434 50766 16436 50818
rect 16268 50764 16436 50766
rect 16156 50194 16212 50204
rect 16380 50036 16436 50764
rect 16492 50482 16548 50988
rect 16716 50820 16772 53004
rect 16940 52834 16996 52846
rect 16940 52782 16942 52834
rect 16994 52782 16996 52834
rect 16940 52276 16996 52782
rect 16940 52210 16996 52220
rect 16716 50754 16772 50764
rect 16940 51266 16996 51278
rect 16940 51214 16942 51266
rect 16994 51214 16996 51266
rect 16492 50430 16494 50482
rect 16546 50430 16548 50482
rect 16492 50418 16548 50430
rect 16380 49970 16436 49980
rect 16940 49924 16996 51214
rect 17052 50596 17108 53004
rect 17164 53284 17220 53294
rect 17164 52274 17220 53228
rect 17164 52222 17166 52274
rect 17218 52222 17220 52274
rect 17164 52210 17220 52222
rect 17276 52948 17332 53452
rect 17276 52164 17332 52892
rect 17276 52098 17332 52108
rect 17052 50530 17108 50540
rect 17164 52052 17220 52062
rect 17164 51604 17220 51996
rect 16940 49858 16996 49868
rect 15820 49646 15822 49698
rect 15874 49646 15876 49698
rect 15820 49634 15876 49646
rect 16044 49700 16100 49710
rect 15484 49586 15540 49598
rect 15484 49534 15486 49586
rect 15538 49534 15540 49586
rect 15484 49364 15540 49534
rect 15484 49298 15540 49308
rect 15596 49028 15652 49038
rect 15596 48580 15652 48972
rect 16044 48804 16100 49644
rect 16492 49698 16548 49710
rect 16492 49646 16494 49698
rect 16546 49646 16548 49698
rect 16492 49252 16548 49646
rect 16940 49700 16996 49710
rect 16940 49606 16996 49644
rect 16492 49186 16548 49196
rect 16044 48710 16100 48748
rect 16380 49140 16436 49150
rect 15484 48468 15540 48478
rect 15484 48354 15540 48412
rect 15484 48302 15486 48354
rect 15538 48302 15540 48354
rect 15484 48290 15540 48302
rect 15372 45838 15374 45890
rect 15426 45838 15428 45890
rect 14812 44324 14868 44334
rect 14588 44322 14868 44324
rect 14588 44270 14814 44322
rect 14866 44270 14868 44322
rect 14588 44268 14868 44270
rect 14812 44258 14868 44268
rect 14924 44212 14980 44222
rect 14924 44118 14980 44156
rect 14588 44098 14644 44110
rect 14588 44046 14590 44098
rect 14642 44046 14644 44098
rect 14588 43540 14644 44046
rect 15372 43876 15428 45838
rect 15148 43820 15428 43876
rect 15484 48020 15540 48030
rect 14700 43764 14756 43774
rect 14700 43670 14756 43708
rect 14700 43540 14756 43550
rect 14588 43538 14756 43540
rect 14588 43486 14702 43538
rect 14754 43486 14756 43538
rect 14588 43484 14756 43486
rect 14028 41468 14532 41524
rect 14588 41972 14644 41982
rect 14028 40852 14084 41468
rect 14140 41188 14196 41198
rect 14140 41094 14196 41132
rect 14252 41076 14308 41086
rect 14252 40982 14308 41020
rect 14364 41074 14420 41086
rect 14364 41022 14366 41074
rect 14418 41022 14420 41074
rect 14028 40796 14196 40852
rect 13916 40628 13972 40638
rect 13916 40534 13972 40572
rect 14028 39394 14084 39406
rect 14028 39342 14030 39394
rect 14082 39342 14084 39394
rect 14028 39172 14084 39342
rect 14028 39106 14084 39116
rect 14140 39060 14196 40796
rect 14364 40628 14420 41022
rect 14364 40562 14420 40572
rect 14476 40740 14532 40750
rect 14476 40626 14532 40684
rect 14476 40574 14478 40626
rect 14530 40574 14532 40626
rect 14476 40562 14532 40574
rect 14364 40402 14420 40414
rect 14364 40350 14366 40402
rect 14418 40350 14420 40402
rect 14364 39844 14420 40350
rect 14588 39844 14644 41916
rect 14700 40628 14756 43484
rect 15036 43538 15092 43550
rect 15036 43486 15038 43538
rect 15090 43486 15092 43538
rect 15036 43428 15092 43486
rect 15148 43428 15204 43820
rect 15484 43764 15540 47964
rect 15596 47572 15652 48524
rect 15708 48692 15764 48702
rect 15708 48466 15764 48636
rect 15708 48414 15710 48466
rect 15762 48414 15764 48466
rect 15708 48402 15764 48414
rect 16156 48580 16212 48590
rect 16156 48356 16212 48524
rect 16044 48354 16212 48356
rect 16044 48302 16158 48354
rect 16210 48302 16212 48354
rect 16044 48300 16212 48302
rect 15932 48244 15988 48254
rect 15932 48150 15988 48188
rect 15596 47506 15652 47516
rect 15708 47460 15764 47470
rect 15708 47366 15764 47404
rect 15932 47460 15988 47470
rect 16044 47460 16100 48300
rect 16156 48290 16212 48300
rect 15932 47458 16100 47460
rect 15932 47406 15934 47458
rect 15986 47406 16100 47458
rect 15932 47404 16100 47406
rect 16268 48130 16324 48142
rect 16268 48078 16270 48130
rect 16322 48078 16324 48130
rect 16268 47458 16324 48078
rect 16268 47406 16270 47458
rect 16322 47406 16324 47458
rect 15820 47234 15876 47246
rect 15820 47182 15822 47234
rect 15874 47182 15876 47234
rect 15708 47124 15764 47134
rect 15596 45332 15652 45342
rect 15596 45238 15652 45276
rect 15708 45108 15764 47068
rect 15820 46788 15876 47182
rect 15932 47124 15988 47404
rect 16268 47394 16324 47406
rect 15932 47058 15988 47068
rect 15820 46722 15876 46732
rect 15820 46564 15876 46574
rect 16380 46564 16436 49084
rect 16940 49140 16996 49150
rect 16940 49046 16996 49084
rect 15820 46562 16436 46564
rect 15820 46510 15822 46562
rect 15874 46510 16382 46562
rect 16434 46510 16436 46562
rect 15820 46508 16436 46510
rect 15820 46498 15876 46508
rect 16044 45780 16100 45790
rect 16044 45686 16100 45724
rect 15260 43708 15540 43764
rect 15596 45052 15764 45108
rect 15260 43540 15316 43708
rect 15260 43484 15428 43540
rect 15036 43372 15316 43428
rect 15148 43092 15204 43102
rect 15148 42866 15204 43036
rect 15148 42814 15150 42866
rect 15202 42814 15204 42866
rect 15148 42802 15204 42814
rect 14924 42196 14980 42206
rect 14924 42102 14980 42140
rect 14812 41970 14868 41982
rect 14812 41918 14814 41970
rect 14866 41918 14868 41970
rect 14812 41410 14868 41918
rect 15036 41970 15092 41982
rect 15036 41918 15038 41970
rect 15090 41918 15092 41970
rect 15036 41748 15092 41918
rect 15036 41682 15092 41692
rect 14812 41358 14814 41410
rect 14866 41358 14868 41410
rect 14812 41346 14868 41358
rect 15260 41636 15316 43372
rect 15260 41412 15316 41580
rect 15260 41346 15316 41356
rect 15372 41300 15428 43484
rect 15484 43426 15540 43438
rect 15484 43374 15486 43426
rect 15538 43374 15540 43426
rect 15484 43316 15540 43374
rect 15484 43250 15540 43260
rect 15596 42532 15652 45052
rect 16156 44994 16212 45006
rect 16156 44942 16158 44994
rect 16210 44942 16212 44994
rect 16156 44772 16212 44942
rect 16156 44706 16212 44716
rect 16156 44548 16212 44558
rect 16380 44548 16436 46508
rect 16492 48804 16548 48814
rect 16492 45892 16548 48748
rect 16940 48468 16996 48478
rect 16940 48374 16996 48412
rect 17164 47572 17220 51548
rect 17500 50596 17556 56140
rect 17612 55972 17668 55982
rect 17612 55878 17668 55916
rect 18172 55970 18228 55982
rect 18172 55918 18174 55970
rect 18226 55918 18228 55970
rect 18172 55524 18228 55918
rect 18508 55636 18564 56252
rect 18620 56242 18676 56252
rect 18508 55570 18564 55580
rect 17836 55074 17892 55086
rect 17836 55022 17838 55074
rect 17890 55022 17892 55074
rect 17836 54964 17892 55022
rect 18172 55076 18228 55468
rect 18956 55410 19012 56702
rect 19180 56754 19236 56924
rect 19180 56702 19182 56754
rect 19234 56702 19236 56754
rect 19180 55970 19236 56702
rect 19180 55918 19182 55970
rect 19234 55918 19236 55970
rect 19180 55906 19236 55918
rect 19292 56194 19348 56206
rect 19292 56142 19294 56194
rect 19346 56142 19348 56194
rect 18956 55358 18958 55410
rect 19010 55358 19012 55410
rect 18956 55346 19012 55358
rect 18732 55300 18788 55310
rect 18732 55206 18788 55244
rect 19180 55300 19236 55310
rect 19068 55188 19124 55198
rect 19068 55094 19124 55132
rect 18172 55020 18564 55076
rect 17836 54898 17892 54908
rect 17612 54404 17668 54414
rect 17612 54402 17780 54404
rect 17612 54350 17614 54402
rect 17666 54350 17780 54402
rect 17612 54348 17780 54350
rect 17612 54338 17668 54348
rect 17724 54292 17780 54348
rect 17612 53506 17668 53518
rect 17612 53454 17614 53506
rect 17666 53454 17668 53506
rect 17612 51268 17668 53454
rect 17724 51492 17780 54236
rect 18060 54402 18116 54414
rect 18060 54350 18062 54402
rect 18114 54350 18116 54402
rect 18060 53506 18116 54350
rect 18508 54180 18564 55020
rect 19068 54628 19124 54638
rect 19180 54628 19236 55244
rect 19068 54626 19236 54628
rect 19068 54574 19070 54626
rect 19122 54574 19236 54626
rect 19068 54572 19236 54574
rect 19292 54628 19348 56142
rect 19068 54562 19124 54572
rect 19292 54562 19348 54572
rect 18620 54404 18676 54414
rect 19404 54404 19460 57036
rect 19516 55860 19572 55870
rect 19516 55766 19572 55804
rect 19628 54740 19684 57260
rect 20524 57204 20580 58158
rect 20636 57540 20692 59388
rect 20972 58212 21028 58222
rect 20972 58118 21028 58156
rect 20972 57540 21028 57550
rect 20636 57538 21028 57540
rect 20636 57486 20974 57538
rect 21026 57486 21028 57538
rect 20636 57484 21028 57486
rect 20188 57092 20244 57102
rect 20188 56978 20244 57036
rect 20188 56926 20190 56978
rect 20242 56926 20244 56978
rect 20188 56914 20244 56926
rect 19852 56644 19908 56682
rect 19852 56578 19908 56588
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 20188 55970 20244 55982
rect 20188 55918 20190 55970
rect 20242 55918 20244 55970
rect 20076 55860 20132 55870
rect 20076 55766 20132 55804
rect 20188 55748 20244 55918
rect 20244 55692 20356 55748
rect 20188 55682 20244 55692
rect 19740 55298 19796 55310
rect 19740 55246 19742 55298
rect 19794 55246 19796 55298
rect 19740 55188 19796 55246
rect 19964 55300 20020 55310
rect 19964 55206 20020 55244
rect 19740 55122 19796 55132
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 20188 54740 20244 54750
rect 19684 54684 19796 54740
rect 18620 54402 18788 54404
rect 18620 54350 18622 54402
rect 18674 54350 18788 54402
rect 18620 54348 18788 54350
rect 18620 54338 18676 54348
rect 18508 54124 18676 54180
rect 18508 53844 18564 53854
rect 18508 53750 18564 53788
rect 18060 53454 18062 53506
rect 18114 53454 18116 53506
rect 18060 52948 18116 53454
rect 18284 53060 18340 53070
rect 18060 52882 18116 52892
rect 18172 53058 18340 53060
rect 18172 53006 18286 53058
rect 18338 53006 18340 53058
rect 18172 53004 18340 53006
rect 18060 52722 18116 52734
rect 18060 52670 18062 52722
rect 18114 52670 18116 52722
rect 17836 52164 17892 52174
rect 17836 51602 17892 52108
rect 17836 51550 17838 51602
rect 17890 51550 17892 51602
rect 17836 51538 17892 51550
rect 17724 51426 17780 51436
rect 17612 50820 17668 51212
rect 17612 50754 17668 50764
rect 18060 51380 18116 52670
rect 18172 52052 18228 53004
rect 18284 52994 18340 53004
rect 18172 51986 18228 51996
rect 18284 52836 18340 52846
rect 18284 52388 18340 52780
rect 18284 52162 18340 52332
rect 18396 52722 18452 52734
rect 18396 52670 18398 52722
rect 18450 52670 18452 52722
rect 18396 52274 18452 52670
rect 18396 52222 18398 52274
rect 18450 52222 18452 52274
rect 18396 52210 18452 52222
rect 18284 52110 18286 52162
rect 18338 52110 18340 52162
rect 18284 51940 18340 52110
rect 18284 51874 18340 51884
rect 18620 51604 18676 54124
rect 18732 53732 18788 54348
rect 18732 53666 18788 53676
rect 19068 54348 19460 54404
rect 19516 54628 19572 54638
rect 19628 54608 19684 54684
rect 19516 54514 19572 54572
rect 19516 54462 19518 54514
rect 19570 54462 19572 54514
rect 19068 53954 19124 54348
rect 19068 53902 19070 53954
rect 19122 53902 19124 53954
rect 19068 53620 19124 53902
rect 19404 54180 19460 54190
rect 19404 53730 19460 54124
rect 19516 53956 19572 54462
rect 19516 53890 19572 53900
rect 19404 53678 19406 53730
rect 19458 53678 19460 53730
rect 19404 53666 19460 53678
rect 19628 53844 19684 53854
rect 19628 53730 19684 53788
rect 19628 53678 19630 53730
rect 19682 53678 19684 53730
rect 19628 53666 19684 53678
rect 19740 53730 19796 54684
rect 19964 54628 20020 54638
rect 19964 54514 20020 54572
rect 19964 54462 19966 54514
rect 20018 54462 20020 54514
rect 19964 54450 20020 54462
rect 19740 53678 19742 53730
rect 19794 53678 19796 53730
rect 19740 53666 19796 53678
rect 19068 53284 19124 53564
rect 19516 53506 19572 53518
rect 19516 53454 19518 53506
rect 19570 53454 19572 53506
rect 19516 53396 19572 53454
rect 19516 53330 19572 53340
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 19068 53218 19124 53228
rect 19852 53060 19908 53070
rect 19852 52966 19908 53004
rect 18956 52836 19012 52846
rect 18956 52742 19012 52780
rect 19516 52834 19572 52846
rect 19516 52782 19518 52834
rect 19570 52782 19572 52834
rect 18508 51548 18676 51604
rect 18732 52722 18788 52734
rect 18732 52670 18734 52722
rect 18786 52670 18788 52722
rect 18284 51380 18340 51390
rect 18060 51378 18340 51380
rect 18060 51326 18286 51378
rect 18338 51326 18340 51378
rect 18060 51324 18340 51326
rect 17500 50540 17780 50596
rect 17612 50372 17668 50382
rect 17724 50372 17780 50540
rect 17612 50370 17780 50372
rect 17612 50318 17614 50370
rect 17666 50318 17780 50370
rect 17612 50316 17780 50318
rect 17276 49924 17332 49934
rect 17276 47684 17332 49868
rect 17612 49812 17668 50316
rect 17836 50260 17892 50270
rect 17724 50148 17780 50158
rect 17724 49922 17780 50092
rect 17836 50034 17892 50204
rect 17836 49982 17838 50034
rect 17890 49982 17892 50034
rect 17836 49970 17892 49982
rect 18060 50034 18116 51324
rect 18284 51314 18340 51324
rect 18172 50820 18228 50830
rect 18172 50706 18228 50764
rect 18172 50654 18174 50706
rect 18226 50654 18228 50706
rect 18172 50428 18228 50654
rect 18396 50596 18452 50606
rect 18172 50372 18340 50428
rect 18060 49982 18062 50034
rect 18114 49982 18116 50034
rect 18060 49970 18116 49982
rect 18172 50260 18228 50270
rect 17724 49870 17726 49922
rect 17778 49870 17780 49922
rect 17724 49858 17780 49870
rect 18172 49812 18228 50204
rect 17612 49746 17668 49756
rect 18060 49756 18228 49812
rect 17388 49700 17444 49710
rect 17388 49138 17444 49644
rect 18060 49364 18116 49756
rect 17388 49086 17390 49138
rect 17442 49086 17444 49138
rect 17388 49074 17444 49086
rect 17500 49252 17556 49262
rect 17276 47628 17444 47684
rect 16828 47516 17220 47572
rect 16604 46676 16660 46686
rect 16604 46582 16660 46620
rect 16492 45826 16548 45836
rect 16604 45444 16660 45454
rect 16492 44996 16548 45006
rect 16492 44902 16548 44940
rect 16212 44492 16436 44548
rect 15820 44324 15876 44334
rect 16044 44324 16100 44334
rect 15820 44230 15876 44268
rect 15932 44322 16100 44324
rect 15932 44270 16046 44322
rect 16098 44270 16100 44322
rect 15932 44268 16100 44270
rect 15708 44100 15764 44110
rect 15708 42754 15764 44044
rect 15708 42702 15710 42754
rect 15762 42702 15764 42754
rect 15708 42690 15764 42702
rect 15820 43988 15876 43998
rect 15596 42476 15764 42532
rect 15596 42308 15652 42318
rect 15596 41972 15652 42252
rect 15596 41840 15652 41916
rect 15484 41300 15540 41310
rect 15372 41298 15652 41300
rect 15372 41246 15486 41298
rect 15538 41246 15652 41298
rect 15372 41244 15652 41246
rect 14700 40562 14756 40572
rect 15036 41076 15092 41086
rect 15036 40628 15092 41020
rect 15372 41076 15428 41244
rect 15484 41234 15540 41244
rect 15372 41010 15428 41020
rect 15036 40626 15204 40628
rect 15036 40574 15038 40626
rect 15090 40574 15204 40626
rect 15036 40572 15204 40574
rect 15036 40562 15092 40572
rect 14700 40404 14756 40414
rect 14700 40402 14980 40404
rect 14700 40350 14702 40402
rect 14754 40350 14980 40402
rect 14700 40348 14980 40350
rect 14700 40338 14756 40348
rect 14812 39956 14868 39966
rect 14588 39788 14756 39844
rect 14364 39778 14420 39788
rect 14588 39620 14644 39630
rect 14140 38994 14196 39004
rect 14364 39618 14644 39620
rect 14364 39566 14590 39618
rect 14642 39566 14644 39618
rect 14364 39564 14644 39566
rect 14028 38948 14084 38958
rect 13804 37538 13860 37548
rect 13916 38050 13972 38062
rect 13916 37998 13918 38050
rect 13970 37998 13972 38050
rect 13692 37324 13860 37380
rect 13356 37268 13412 37278
rect 13132 34962 13188 34972
rect 13244 37266 13412 37268
rect 13244 37214 13358 37266
rect 13410 37214 13412 37266
rect 13244 37212 13412 37214
rect 13020 34692 13076 34702
rect 13244 34692 13300 37212
rect 13356 37202 13412 37212
rect 13580 37268 13636 37278
rect 13076 34636 13300 34692
rect 13356 36820 13412 36830
rect 13356 35700 13412 36764
rect 13580 36708 13636 37212
rect 13692 37156 13748 37166
rect 13692 37062 13748 37100
rect 13580 36642 13636 36652
rect 13804 36708 13860 37324
rect 13916 37044 13972 37998
rect 13916 36978 13972 36988
rect 13804 36642 13860 36652
rect 13916 36482 13972 36494
rect 13916 36430 13918 36482
rect 13970 36430 13972 36482
rect 13804 36372 13860 36382
rect 13580 36316 13804 36372
rect 13468 35924 13524 35934
rect 13468 35830 13524 35868
rect 12796 34244 12852 34254
rect 12796 34150 12852 34188
rect 13020 34130 13076 34636
rect 13020 34078 13022 34130
rect 13074 34078 13076 34130
rect 13020 34066 13076 34078
rect 13020 33908 13076 33918
rect 13020 33796 13076 33852
rect 12684 33740 13076 33796
rect 12908 33572 12964 33582
rect 12908 33460 12964 33516
rect 12460 33282 12516 33292
rect 12684 33458 12964 33460
rect 12684 33406 12910 33458
rect 12962 33406 12964 33458
rect 12684 33404 12964 33406
rect 11788 33236 11844 33246
rect 11788 33234 11956 33236
rect 11788 33182 11790 33234
rect 11842 33182 11956 33234
rect 11788 33180 11956 33182
rect 11788 33170 11844 33180
rect 11676 32562 11732 32574
rect 11676 32510 11678 32562
rect 11730 32510 11732 32562
rect 11676 32452 11732 32510
rect 11676 32386 11732 32396
rect 11676 31780 11732 31790
rect 11676 30324 11732 31724
rect 11900 30996 11956 33180
rect 12460 33122 12516 33134
rect 12460 33070 12462 33122
rect 12514 33070 12516 33122
rect 12124 32900 12180 32910
rect 12124 32674 12180 32844
rect 12124 32622 12126 32674
rect 12178 32622 12180 32674
rect 12124 32610 12180 32622
rect 12348 32452 12404 32462
rect 12348 32358 12404 32396
rect 12460 32004 12516 33070
rect 12572 33012 12628 33022
rect 12572 32562 12628 32956
rect 12572 32510 12574 32562
rect 12626 32510 12628 32562
rect 12572 32116 12628 32510
rect 12572 32050 12628 32060
rect 12684 32564 12740 33404
rect 12908 33394 12964 33404
rect 12348 31948 12516 32004
rect 12012 31892 12068 31902
rect 12012 31556 12068 31836
rect 12012 31462 12068 31500
rect 12236 31444 12292 31454
rect 11900 30930 11956 30940
rect 12124 31332 12180 31342
rect 12124 31218 12180 31276
rect 12124 31166 12126 31218
rect 12178 31166 12180 31218
rect 11676 30258 11732 30268
rect 11788 30548 11844 30558
rect 11676 30098 11732 30110
rect 11676 30046 11678 30098
rect 11730 30046 11732 30098
rect 11676 29764 11732 30046
rect 11676 29698 11732 29708
rect 11676 29540 11732 29550
rect 11676 28532 11732 29484
rect 11788 29204 11844 30492
rect 11900 30324 11956 30334
rect 11900 30210 11956 30268
rect 11900 30158 11902 30210
rect 11954 30158 11956 30210
rect 11900 30146 11956 30158
rect 12012 30322 12068 30334
rect 12012 30270 12014 30322
rect 12066 30270 12068 30322
rect 11788 29148 11956 29204
rect 11788 28756 11844 28766
rect 11788 28662 11844 28700
rect 11676 28476 11844 28532
rect 11788 26908 11844 28476
rect 11900 27858 11956 29148
rect 11900 27806 11902 27858
rect 11954 27806 11956 27858
rect 11900 27794 11956 27806
rect 12012 27636 12068 30270
rect 12124 29650 12180 31166
rect 12236 29764 12292 31388
rect 12348 30100 12404 31948
rect 12460 31554 12516 31566
rect 12460 31502 12462 31554
rect 12514 31502 12516 31554
rect 12460 31332 12516 31502
rect 12460 31266 12516 31276
rect 12572 31556 12628 31566
rect 12572 30322 12628 31500
rect 12684 31218 12740 32508
rect 12908 31892 12964 31902
rect 13020 31892 13076 33740
rect 12908 31890 13076 31892
rect 12908 31838 12910 31890
rect 12962 31838 13076 31890
rect 12908 31836 13076 31838
rect 13244 33796 13300 33806
rect 12908 31780 12964 31836
rect 12908 31714 12964 31724
rect 12684 31166 12686 31218
rect 12738 31166 12740 31218
rect 12684 31154 12740 31166
rect 13132 31668 13188 31678
rect 13132 31218 13188 31612
rect 13132 31166 13134 31218
rect 13186 31166 13188 31218
rect 13132 31154 13188 31166
rect 12572 30270 12574 30322
rect 12626 30270 12628 30322
rect 12572 30258 12628 30270
rect 13132 30324 13188 30334
rect 12348 30034 12404 30044
rect 12908 30100 12964 30110
rect 12908 29988 12964 30044
rect 12908 29986 13076 29988
rect 12908 29934 12910 29986
rect 12962 29934 13076 29986
rect 12908 29932 13076 29934
rect 12908 29922 12964 29932
rect 12236 29698 12292 29708
rect 12796 29876 12852 29886
rect 12124 29598 12126 29650
rect 12178 29598 12180 29650
rect 12124 29586 12180 29598
rect 12684 29652 12740 29662
rect 12684 29558 12740 29596
rect 12796 28756 12852 29820
rect 12572 28644 12628 28654
rect 12348 28532 12404 28542
rect 12348 28438 12404 28476
rect 12572 28418 12628 28588
rect 12572 28366 12574 28418
rect 12626 28366 12628 28418
rect 12572 28354 12628 28366
rect 12684 28644 12740 28654
rect 12796 28644 12852 28700
rect 12684 28642 12852 28644
rect 12684 28590 12686 28642
rect 12738 28590 12852 28642
rect 12684 28588 12852 28590
rect 12908 29540 12964 29550
rect 12908 28642 12964 29484
rect 13020 28756 13076 29932
rect 13132 29204 13188 30268
rect 13244 29540 13300 33740
rect 13356 31780 13412 35644
rect 13468 35252 13524 35262
rect 13468 33796 13524 35196
rect 13468 33730 13524 33740
rect 13580 32900 13636 36316
rect 13804 36278 13860 36316
rect 13692 35812 13748 35822
rect 13692 34356 13748 35756
rect 13692 34290 13748 34300
rect 13804 35698 13860 35710
rect 13804 35646 13806 35698
rect 13858 35646 13860 35698
rect 13804 35588 13860 35646
rect 13692 34130 13748 34142
rect 13692 34078 13694 34130
rect 13746 34078 13748 34130
rect 13692 33796 13748 34078
rect 13692 33730 13748 33740
rect 13804 33236 13860 35532
rect 13916 35364 13972 36430
rect 13916 35298 13972 35308
rect 13804 33170 13860 33180
rect 13916 34914 13972 34926
rect 13916 34862 13918 34914
rect 13970 34862 13972 34914
rect 13468 32844 13636 32900
rect 13916 32900 13972 34862
rect 14028 34020 14084 38892
rect 14252 38834 14308 38846
rect 14252 38782 14254 38834
rect 14306 38782 14308 38834
rect 14252 38276 14308 38782
rect 14364 38668 14420 39564
rect 14588 39554 14644 39564
rect 14700 39396 14756 39788
rect 14476 39340 14756 39396
rect 14476 38948 14532 39340
rect 14476 38816 14532 38892
rect 14588 39058 14644 39070
rect 14588 39006 14590 39058
rect 14642 39006 14644 39058
rect 14364 38612 14532 38668
rect 14252 38210 14308 38220
rect 14364 37938 14420 37950
rect 14364 37886 14366 37938
rect 14418 37886 14420 37938
rect 14364 37828 14420 37886
rect 14140 37772 14420 37828
rect 14140 34242 14196 37772
rect 14364 37604 14420 37614
rect 14252 36708 14308 36718
rect 14252 35922 14308 36652
rect 14364 36260 14420 37548
rect 14476 36596 14532 38612
rect 14588 37154 14644 39006
rect 14812 38946 14868 39900
rect 14924 39618 14980 40348
rect 14924 39566 14926 39618
rect 14978 39566 14980 39618
rect 14924 39554 14980 39566
rect 15036 39730 15092 39742
rect 15036 39678 15038 39730
rect 15090 39678 15092 39730
rect 15036 39172 15092 39678
rect 15148 39620 15204 40572
rect 15260 40516 15316 40526
rect 15260 40422 15316 40460
rect 15372 40402 15428 40414
rect 15372 40350 15374 40402
rect 15426 40350 15428 40402
rect 15372 40180 15428 40350
rect 15372 39844 15428 40124
rect 15372 39778 15428 39788
rect 15372 39620 15428 39630
rect 15148 39618 15428 39620
rect 15148 39566 15374 39618
rect 15426 39566 15428 39618
rect 15148 39564 15428 39566
rect 15372 39554 15428 39564
rect 15148 39396 15204 39406
rect 15148 39302 15204 39340
rect 15036 39106 15092 39116
rect 14812 38894 14814 38946
rect 14866 38894 14868 38946
rect 14812 38836 14868 38894
rect 14812 38770 14868 38780
rect 14924 39060 14980 39070
rect 14924 38668 14980 39004
rect 15484 39060 15540 39070
rect 15484 38966 15540 39004
rect 15372 38948 15428 38958
rect 15372 38854 15428 38892
rect 15596 38948 15652 41244
rect 15708 40964 15764 42476
rect 15820 41188 15876 43932
rect 15932 42866 15988 44268
rect 16044 44258 16100 44268
rect 16156 43316 16212 44492
rect 16380 44100 16436 44110
rect 16380 44006 16436 44044
rect 16156 43250 16212 43260
rect 16268 43652 16324 43662
rect 15932 42814 15934 42866
rect 15986 42814 15988 42866
rect 15932 42802 15988 42814
rect 16156 43092 16212 43102
rect 16044 42644 16100 42654
rect 16044 42550 16100 42588
rect 16156 42642 16212 43036
rect 16156 42590 16158 42642
rect 16210 42590 16212 42642
rect 16156 42578 16212 42590
rect 15932 42532 15988 42542
rect 15932 42438 15988 42476
rect 16044 41858 16100 41870
rect 16044 41806 16046 41858
rect 16098 41806 16100 41858
rect 16044 41636 16100 41806
rect 16044 41570 16100 41580
rect 15820 41132 16212 41188
rect 15932 40964 15988 40974
rect 15708 40962 15988 40964
rect 15708 40910 15934 40962
rect 15986 40910 15988 40962
rect 15708 40908 15988 40910
rect 15708 39396 15764 39406
rect 15708 39058 15764 39340
rect 15708 39006 15710 39058
rect 15762 39006 15764 39058
rect 15708 38994 15764 39006
rect 14588 37102 14590 37154
rect 14642 37102 14644 37154
rect 14588 37090 14644 37102
rect 14700 38612 14980 38668
rect 14476 36530 14532 36540
rect 14588 36708 14644 36718
rect 14588 36482 14644 36652
rect 14588 36430 14590 36482
rect 14642 36430 14644 36482
rect 14588 36418 14644 36430
rect 14476 36372 14532 36382
rect 14476 36278 14532 36316
rect 14364 36194 14420 36204
rect 14252 35870 14254 35922
rect 14306 35870 14308 35922
rect 14252 35700 14308 35870
rect 14252 35634 14308 35644
rect 14588 35700 14644 35710
rect 14140 34190 14142 34242
rect 14194 34190 14196 34242
rect 14140 34178 14196 34190
rect 14252 35140 14308 35150
rect 14252 35026 14308 35084
rect 14252 34974 14254 35026
rect 14306 34974 14308 35026
rect 14252 34916 14308 34974
rect 14028 33954 14084 33964
rect 14252 33684 14308 34860
rect 14476 34804 14532 34814
rect 14364 34748 14476 34804
rect 14364 34130 14420 34748
rect 14476 34710 14532 34748
rect 14364 34078 14366 34130
rect 14418 34078 14420 34130
rect 14364 34066 14420 34078
rect 14588 33908 14644 35644
rect 13468 32676 13524 32844
rect 13804 32788 13860 32798
rect 13804 32694 13860 32732
rect 13468 32544 13524 32620
rect 13580 32674 13636 32686
rect 13580 32622 13582 32674
rect 13634 32622 13636 32674
rect 13580 32564 13636 32622
rect 13916 32564 13972 32844
rect 13580 32498 13636 32508
rect 13804 32508 13972 32564
rect 14028 33628 14308 33684
rect 14364 33852 14644 33908
rect 13692 31892 13748 31902
rect 13580 31780 13636 31790
rect 13356 31778 13636 31780
rect 13356 31726 13582 31778
rect 13634 31726 13636 31778
rect 13356 31724 13636 31726
rect 13244 29408 13300 29484
rect 13132 29148 13412 29204
rect 13020 28690 13076 28700
rect 13132 28868 13188 28878
rect 12908 28590 12910 28642
rect 12962 28590 12964 28642
rect 12012 27580 12404 27636
rect 12124 27188 12180 27198
rect 12124 27094 12180 27132
rect 12012 27076 12068 27086
rect 12012 26982 12068 27020
rect 11564 26674 11620 26684
rect 11676 26852 11732 26862
rect 11788 26852 11956 26908
rect 11900 26796 12068 26852
rect 11228 26348 11452 26404
rect 11228 26290 11284 26348
rect 11452 26338 11508 26348
rect 11676 26402 11732 26796
rect 11676 26350 11678 26402
rect 11730 26350 11732 26402
rect 11676 26338 11732 26350
rect 11228 26238 11230 26290
rect 11282 26238 11284 26290
rect 11228 26226 11284 26238
rect 11452 26180 11508 26190
rect 11452 26086 11508 26124
rect 11564 26178 11620 26190
rect 11564 26126 11566 26178
rect 11618 26126 11620 26178
rect 11564 25508 11620 26126
rect 11676 25620 11732 25630
rect 11676 25526 11732 25564
rect 11452 25452 11620 25508
rect 11788 25508 11844 25518
rect 11340 25394 11396 25406
rect 11340 25342 11342 25394
rect 11394 25342 11396 25394
rect 11340 25284 11396 25342
rect 11340 25218 11396 25228
rect 11116 25004 11396 25060
rect 11004 24834 11060 24846
rect 11004 24782 11006 24834
rect 11058 24782 11060 24834
rect 11004 23828 11060 24782
rect 11004 23762 11060 23772
rect 11228 23940 11284 23950
rect 10892 23548 11060 23604
rect 10892 23268 10948 23278
rect 10892 23174 10948 23212
rect 10108 23042 10724 23044
rect 10108 22990 10110 23042
rect 10162 22990 10724 23042
rect 10108 22988 10724 22990
rect 10780 23156 10836 23166
rect 8764 16098 9492 16100
rect 8764 16046 8766 16098
rect 8818 16046 9492 16098
rect 8764 16044 9492 16046
rect 9548 17666 9604 17678
rect 9548 17614 9550 17666
rect 9602 17614 9604 17666
rect 8764 16034 8820 16044
rect 8316 15316 8372 15326
rect 8316 15222 8372 15260
rect 8652 15204 8708 15214
rect 7756 14642 8036 14644
rect 7756 14590 7758 14642
rect 7810 14590 8036 14642
rect 7756 14588 8036 14590
rect 7756 14578 7812 14588
rect 7980 13972 8036 14588
rect 8092 14578 8148 14588
rect 8204 14754 8260 14766
rect 8204 14702 8206 14754
rect 8258 14702 8260 14754
rect 8204 14306 8260 14702
rect 8204 14254 8206 14306
rect 8258 14254 8260 14306
rect 8092 13972 8148 13982
rect 7980 13970 8148 13972
rect 7980 13918 8094 13970
rect 8146 13918 8148 13970
rect 7980 13916 8148 13918
rect 6188 12964 6244 12974
rect 6076 12962 6244 12964
rect 6076 12910 6190 12962
rect 6242 12910 6244 12962
rect 6076 12908 6244 12910
rect 6076 11282 6132 12908
rect 6188 12898 6244 12908
rect 8092 12964 8148 13916
rect 6188 12404 6244 12414
rect 6188 12310 6244 12348
rect 8092 12404 8148 12908
rect 6972 12180 7028 12190
rect 6636 11396 6692 11406
rect 6636 11302 6692 11340
rect 6076 11230 6078 11282
rect 6130 11230 6132 11282
rect 6076 11218 6132 11230
rect 6972 11282 7028 12124
rect 8092 11506 8148 12348
rect 8092 11454 8094 11506
rect 8146 11454 8148 11506
rect 8092 11442 8148 11454
rect 6972 11230 6974 11282
rect 7026 11230 7028 11282
rect 6972 11218 7028 11230
rect 6076 9604 6132 9614
rect 5964 9602 6132 9604
rect 5964 9550 6078 9602
rect 6130 9550 6132 9602
rect 5964 9548 6132 9550
rect 5964 9042 6020 9548
rect 6076 9538 6132 9548
rect 5964 8990 5966 9042
rect 6018 8990 6020 9042
rect 5964 8978 6020 8990
rect 7644 9156 7700 9166
rect 5740 8372 5908 8428
rect 6748 8372 6804 8382
rect 5516 5908 5572 6412
rect 5628 6580 5684 6590
rect 5628 6468 5684 6524
rect 5740 6468 5796 8372
rect 6748 8278 6804 8316
rect 7196 8036 7252 8046
rect 6188 7586 6244 7598
rect 6188 7534 6190 7586
rect 6242 7534 6244 7586
rect 5628 6466 5796 6468
rect 5628 6414 5630 6466
rect 5682 6414 5796 6466
rect 5628 6412 5796 6414
rect 5628 6402 5684 6412
rect 5628 5908 5684 5918
rect 5516 5906 5684 5908
rect 5516 5854 5630 5906
rect 5682 5854 5684 5906
rect 5516 5852 5684 5854
rect 5068 5170 5124 5180
rect 4956 4956 5124 5012
rect 4284 4116 4340 4126
rect 4284 800 4340 4060
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 5068 3556 5124 4956
rect 5628 4338 5684 5852
rect 5628 4286 5630 4338
rect 5682 4286 5684 4338
rect 5628 4274 5684 4286
rect 5740 3780 5796 6412
rect 5852 7474 5908 7486
rect 5852 7422 5854 7474
rect 5906 7422 5908 7474
rect 5852 5346 5908 7422
rect 6076 5908 6132 5918
rect 6188 5908 6244 7534
rect 6748 6690 6804 6702
rect 6748 6638 6750 6690
rect 6802 6638 6804 6690
rect 6524 6468 6580 6478
rect 6076 5906 6244 5908
rect 6076 5854 6078 5906
rect 6130 5854 6244 5906
rect 6076 5852 6244 5854
rect 6300 6466 6580 6468
rect 6300 6414 6526 6466
rect 6578 6414 6580 6466
rect 6300 6412 6580 6414
rect 6076 5842 6132 5852
rect 5852 5294 5854 5346
rect 5906 5294 5908 5346
rect 5852 5282 5908 5294
rect 5964 5236 6020 5246
rect 5964 5142 6020 5180
rect 6076 4340 6132 4350
rect 6300 4340 6356 6412
rect 6524 6402 6580 6412
rect 6636 6132 6692 6142
rect 6636 5122 6692 6076
rect 6636 5070 6638 5122
rect 6690 5070 6692 5122
rect 6636 5058 6692 5070
rect 6748 4900 6804 6638
rect 7196 6580 7252 7980
rect 7644 6692 7700 9100
rect 8204 8428 8260 14254
rect 8428 12180 8484 12190
rect 8428 12086 8484 12124
rect 8540 11282 8596 11294
rect 8540 11230 8542 11282
rect 8594 11230 8596 11282
rect 8540 11172 8596 11230
rect 8540 11106 8596 11116
rect 8428 9940 8484 9950
rect 8652 9940 8708 15148
rect 8764 14756 8820 14766
rect 8764 14642 8820 14700
rect 8764 14590 8766 14642
rect 8818 14590 8820 14642
rect 8764 13972 8820 14590
rect 9548 14644 9604 17614
rect 9660 17108 9716 18396
rect 9772 20132 9940 20188
rect 10108 20188 10164 22988
rect 10220 22484 10276 22494
rect 10220 22390 10276 22428
rect 10668 22484 10724 22494
rect 10780 22484 10836 23100
rect 10668 22482 10836 22484
rect 10668 22430 10670 22482
rect 10722 22430 10836 22482
rect 10668 22428 10836 22430
rect 10668 22418 10724 22428
rect 10556 21700 10612 21710
rect 10444 21698 10612 21700
rect 10444 21646 10558 21698
rect 10610 21646 10612 21698
rect 10444 21644 10612 21646
rect 10332 21586 10388 21598
rect 10332 21534 10334 21586
rect 10386 21534 10388 21586
rect 10332 20916 10388 21534
rect 10332 20850 10388 20860
rect 10332 20580 10388 20590
rect 10108 20132 10276 20188
rect 9772 17668 9828 20132
rect 9996 19906 10052 19918
rect 9996 19854 9998 19906
rect 10050 19854 10052 19906
rect 9884 19236 9940 19246
rect 9996 19236 10052 19854
rect 9884 19234 10052 19236
rect 9884 19182 9886 19234
rect 9938 19182 10052 19234
rect 9884 19180 10052 19182
rect 10108 19348 10164 19358
rect 9884 19170 9940 19180
rect 10108 18450 10164 19292
rect 10220 19124 10276 20132
rect 10220 18676 10276 19068
rect 10220 18610 10276 18620
rect 10108 18398 10110 18450
rect 10162 18398 10164 18450
rect 10108 18386 10164 18398
rect 9884 17668 9940 17678
rect 9772 17666 9940 17668
rect 9772 17614 9886 17666
rect 9938 17614 9940 17666
rect 9772 17612 9940 17614
rect 9884 17602 9940 17612
rect 9772 17108 9828 17118
rect 9660 17106 9828 17108
rect 9660 17054 9774 17106
rect 9826 17054 9828 17106
rect 9660 17052 9828 17054
rect 9772 17042 9828 17052
rect 10220 17108 10276 17118
rect 10220 17014 10276 17052
rect 10332 16658 10388 20524
rect 10444 20020 10500 21644
rect 10556 21634 10612 21644
rect 10668 21588 10724 21598
rect 10668 20188 10724 21532
rect 10892 20804 10948 20814
rect 10892 20690 10948 20748
rect 10892 20638 10894 20690
rect 10946 20638 10948 20690
rect 10892 20626 10948 20638
rect 11004 20188 11060 23548
rect 11228 23380 11284 23884
rect 11116 23324 11228 23380
rect 11116 22820 11172 23324
rect 11228 23314 11284 23324
rect 11228 23156 11284 23166
rect 11228 23062 11284 23100
rect 11116 22764 11284 22820
rect 11116 22260 11172 22270
rect 11116 22166 11172 22204
rect 10668 20132 10836 20188
rect 10668 20020 10724 20030
rect 10444 19964 10668 20020
rect 10668 19926 10724 19964
rect 10780 19906 10836 20132
rect 10780 19854 10782 19906
rect 10834 19854 10836 19906
rect 10780 19842 10836 19854
rect 10892 20132 11060 20188
rect 11116 20244 11172 20254
rect 10556 19348 10612 19358
rect 10892 19348 10948 20132
rect 10556 19346 10948 19348
rect 10556 19294 10558 19346
rect 10610 19294 10948 19346
rect 10556 19292 10948 19294
rect 11004 19348 11060 19358
rect 10556 19282 10612 19292
rect 11004 19254 11060 19292
rect 10556 18676 10612 18686
rect 10556 18582 10612 18620
rect 11116 18226 11172 20188
rect 11116 18174 11118 18226
rect 11170 18174 11172 18226
rect 11116 18162 11172 18174
rect 11228 17668 11284 22764
rect 11340 19348 11396 25004
rect 11452 24724 11508 25452
rect 11788 25414 11844 25452
rect 11564 25284 11620 25294
rect 11564 25190 11620 25228
rect 11900 25282 11956 25294
rect 11900 25230 11902 25282
rect 11954 25230 11956 25282
rect 11900 24946 11956 25230
rect 11900 24894 11902 24946
rect 11954 24894 11956 24946
rect 11900 24882 11956 24894
rect 11564 24724 11620 24734
rect 11452 24722 11620 24724
rect 11452 24670 11566 24722
rect 11618 24670 11620 24722
rect 11452 24668 11620 24670
rect 11564 24658 11620 24668
rect 11900 24722 11956 24734
rect 11900 24670 11902 24722
rect 11954 24670 11956 24722
rect 11452 24388 11508 24398
rect 11452 23938 11508 24332
rect 11788 24164 11844 24174
rect 11900 24164 11956 24670
rect 11788 24162 11956 24164
rect 11788 24110 11790 24162
rect 11842 24110 11956 24162
rect 11788 24108 11956 24110
rect 11788 24098 11844 24108
rect 11452 23886 11454 23938
rect 11506 23886 11508 23938
rect 11452 23874 11508 23886
rect 11676 23828 11732 23838
rect 11676 23734 11732 23772
rect 11900 23716 11956 23726
rect 11788 23380 11844 23390
rect 11788 23286 11844 23324
rect 11900 23156 11956 23660
rect 11788 23100 11956 23156
rect 11564 22930 11620 22942
rect 11564 22878 11566 22930
rect 11618 22878 11620 22930
rect 11564 22482 11620 22878
rect 11564 22430 11566 22482
rect 11618 22430 11620 22482
rect 11564 22418 11620 22430
rect 11452 22260 11508 22270
rect 11452 21810 11508 22204
rect 11452 21758 11454 21810
rect 11506 21758 11508 21810
rect 11452 21746 11508 21758
rect 11676 21476 11732 21486
rect 11564 20690 11620 20702
rect 11564 20638 11566 20690
rect 11618 20638 11620 20690
rect 11564 20020 11620 20638
rect 11676 20578 11732 21420
rect 11788 21474 11844 23100
rect 11788 21422 11790 21474
rect 11842 21422 11844 21474
rect 11788 21362 11844 21422
rect 11788 21310 11790 21362
rect 11842 21310 11844 21362
rect 11788 21298 11844 21310
rect 11900 22930 11956 22942
rect 11900 22878 11902 22930
rect 11954 22878 11956 22930
rect 11788 20804 11844 20814
rect 11788 20710 11844 20748
rect 11676 20526 11678 20578
rect 11730 20526 11732 20578
rect 11676 20514 11732 20526
rect 11452 19348 11508 19358
rect 11340 19346 11508 19348
rect 11340 19294 11454 19346
rect 11506 19294 11508 19346
rect 11340 19292 11508 19294
rect 11452 19282 11508 19292
rect 11564 19124 11620 19964
rect 11564 19058 11620 19068
rect 11676 20130 11732 20142
rect 11676 20078 11678 20130
rect 11730 20078 11732 20130
rect 11340 19012 11396 19022
rect 11340 18674 11396 18956
rect 11340 18622 11342 18674
rect 11394 18622 11396 18674
rect 11340 18610 11396 18622
rect 11676 18564 11732 20078
rect 11900 19348 11956 22878
rect 12012 22260 12068 26796
rect 12236 26850 12292 26862
rect 12236 26798 12238 26850
rect 12290 26798 12292 26850
rect 12124 26404 12180 26414
rect 12124 23378 12180 26348
rect 12236 25844 12292 26798
rect 12236 25778 12292 25788
rect 12348 25508 12404 27580
rect 12460 27300 12516 27310
rect 12460 26962 12516 27244
rect 12460 26910 12462 26962
rect 12514 26910 12516 26962
rect 12460 26852 12516 26910
rect 12460 26786 12516 26796
rect 12572 26290 12628 26302
rect 12572 26238 12574 26290
rect 12626 26238 12628 26290
rect 12348 25442 12404 25452
rect 12460 26180 12516 26190
rect 12236 24948 12292 24958
rect 12236 24836 12292 24892
rect 12236 24834 12404 24836
rect 12236 24782 12238 24834
rect 12290 24782 12404 24834
rect 12236 24780 12404 24782
rect 12236 24770 12292 24780
rect 12124 23326 12126 23378
rect 12178 23326 12180 23378
rect 12124 22930 12180 23326
rect 12124 22878 12126 22930
rect 12178 22878 12180 22930
rect 12124 22866 12180 22878
rect 12348 22372 12404 24780
rect 12460 24050 12516 26124
rect 12572 25844 12628 26238
rect 12572 25778 12628 25788
rect 12572 25508 12628 25518
rect 12572 25414 12628 25452
rect 12460 23998 12462 24050
rect 12514 23998 12516 24050
rect 12460 23828 12516 23998
rect 12460 23762 12516 23772
rect 12348 22316 12516 22372
rect 12012 22194 12068 22204
rect 12124 22146 12180 22158
rect 12124 22094 12126 22146
rect 12178 22094 12180 22146
rect 12012 21362 12068 21374
rect 12012 21310 12014 21362
rect 12066 21310 12068 21362
rect 12012 20188 12068 21310
rect 12124 21364 12180 22094
rect 12236 22148 12292 22158
rect 12236 22054 12292 22092
rect 12348 22146 12404 22158
rect 12348 22094 12350 22146
rect 12402 22094 12404 22146
rect 12348 22036 12404 22094
rect 12124 21298 12180 21308
rect 12236 21588 12292 21598
rect 12124 21140 12180 21150
rect 12124 20356 12180 21084
rect 12236 20804 12292 21532
rect 12348 21140 12404 21980
rect 12348 21074 12404 21084
rect 12236 20738 12292 20748
rect 12348 20916 12404 20926
rect 12236 20580 12292 20590
rect 12348 20580 12404 20860
rect 12236 20578 12404 20580
rect 12236 20526 12238 20578
rect 12290 20526 12404 20578
rect 12236 20524 12404 20526
rect 12236 20514 12292 20524
rect 12124 20300 12404 20356
rect 12012 20132 12180 20188
rect 12012 20020 12068 20030
rect 12012 19926 12068 19964
rect 12124 19572 12180 20132
rect 11900 19282 11956 19292
rect 12012 19516 12180 19572
rect 11564 18508 11732 18564
rect 11788 19124 11844 19134
rect 10332 16606 10334 16658
rect 10386 16606 10388 16658
rect 10332 16594 10388 16606
rect 10556 17612 11284 17668
rect 11340 18226 11396 18238
rect 11340 18174 11342 18226
rect 11394 18174 11396 18226
rect 10220 15988 10276 15998
rect 9660 15204 9716 15214
rect 9660 15110 9716 15148
rect 9996 15204 10052 15214
rect 9548 14530 9604 14588
rect 9548 14478 9550 14530
rect 9602 14478 9604 14530
rect 8876 13972 8932 13982
rect 8764 13970 8932 13972
rect 8764 13918 8878 13970
rect 8930 13918 8932 13970
rect 8764 13916 8932 13918
rect 9548 13972 9604 14478
rect 9996 14530 10052 15148
rect 9996 14478 9998 14530
rect 10050 14478 10052 14530
rect 9996 14466 10052 14478
rect 9660 13972 9716 13982
rect 10108 13972 10164 13982
rect 9548 13970 10164 13972
rect 9548 13918 9662 13970
rect 9714 13918 10110 13970
rect 10162 13918 10164 13970
rect 9548 13916 10164 13918
rect 8876 13906 8932 13916
rect 8764 12964 8820 12974
rect 8764 12740 8820 12908
rect 9324 12740 9380 12750
rect 8764 12646 8820 12684
rect 8988 12738 9380 12740
rect 8988 12686 9326 12738
rect 9378 12686 9380 12738
rect 8988 12684 9380 12686
rect 8988 11394 9044 12684
rect 9324 12674 9380 12684
rect 9660 12404 9716 13916
rect 10108 13748 10164 13916
rect 10108 13682 10164 13692
rect 10108 13412 10164 13422
rect 9884 12852 9940 12862
rect 9884 12758 9940 12796
rect 8988 11342 8990 11394
rect 9042 11342 9044 11394
rect 8988 11330 9044 11342
rect 9100 12402 9716 12404
rect 9100 12350 9662 12402
rect 9714 12350 9716 12402
rect 9100 12348 9716 12350
rect 9100 12178 9156 12348
rect 9660 12338 9716 12348
rect 10108 12740 10164 13356
rect 10220 13188 10276 15932
rect 10556 15538 10612 17612
rect 10668 17108 10724 17118
rect 11340 17108 11396 18174
rect 10668 17106 11396 17108
rect 10668 17054 10670 17106
rect 10722 17054 11396 17106
rect 10668 17052 11396 17054
rect 10668 17042 10724 17052
rect 11228 16884 11284 16894
rect 11228 16790 11284 16828
rect 10556 15486 10558 15538
rect 10610 15486 10612 15538
rect 10556 15474 10612 15486
rect 10892 16658 10948 16670
rect 10892 16606 10894 16658
rect 10946 16606 10948 16658
rect 10892 15540 10948 16606
rect 11116 15874 11172 15886
rect 11116 15822 11118 15874
rect 11170 15822 11172 15874
rect 11004 15540 11060 15550
rect 10892 15538 11060 15540
rect 10892 15486 11006 15538
rect 11058 15486 11060 15538
rect 10892 15484 11060 15486
rect 11004 15474 11060 15484
rect 10556 13748 10612 13758
rect 10556 13654 10612 13692
rect 10892 13748 10948 13758
rect 10220 13186 10724 13188
rect 10220 13134 10222 13186
rect 10274 13134 10724 13186
rect 10220 13132 10724 13134
rect 10220 13122 10276 13132
rect 10444 12964 10500 12974
rect 10444 12870 10500 12908
rect 10108 12402 10164 12684
rect 10108 12350 10110 12402
rect 10162 12350 10164 12402
rect 10108 12338 10164 12350
rect 10668 12402 10724 13132
rect 10892 13074 10948 13692
rect 11116 13412 11172 15822
rect 11564 15204 11620 18508
rect 11676 18338 11732 18350
rect 11676 18286 11678 18338
rect 11730 18286 11732 18338
rect 11676 18226 11732 18286
rect 11676 18174 11678 18226
rect 11730 18174 11732 18226
rect 11676 18162 11732 18174
rect 11788 16322 11844 19068
rect 12012 17108 12068 19516
rect 12124 19348 12180 19358
rect 12348 19348 12404 20300
rect 12460 20188 12516 22316
rect 12684 22148 12740 28588
rect 12908 28578 12964 28590
rect 12796 26852 12852 26862
rect 12796 26066 12852 26796
rect 13020 26852 13076 26862
rect 12908 26180 12964 26190
rect 12908 26086 12964 26124
rect 12796 26014 12798 26066
rect 12850 26014 12852 26066
rect 12796 26002 12852 26014
rect 13020 25618 13076 26796
rect 13020 25566 13022 25618
rect 13074 25566 13076 25618
rect 13020 25554 13076 25566
rect 13132 25508 13188 28812
rect 13244 28196 13300 28206
rect 13244 28082 13300 28140
rect 13244 28030 13246 28082
rect 13298 28030 13300 28082
rect 13244 28018 13300 28030
rect 13356 27636 13412 29148
rect 13356 27570 13412 27580
rect 13132 25442 13188 25452
rect 13244 26404 13300 26414
rect 13244 24834 13300 26348
rect 13468 26292 13524 31724
rect 13580 31714 13636 31724
rect 13692 31220 13748 31836
rect 13580 31218 13748 31220
rect 13580 31166 13694 31218
rect 13746 31166 13748 31218
rect 13580 31164 13748 31166
rect 13580 29988 13636 31164
rect 13692 31154 13748 31164
rect 13804 30994 13860 32508
rect 13916 31780 13972 31790
rect 14028 31780 14084 33628
rect 14252 33458 14308 33470
rect 14252 33406 14254 33458
rect 14306 33406 14308 33458
rect 14252 33236 14308 33406
rect 14364 33346 14420 33852
rect 14364 33294 14366 33346
rect 14418 33294 14420 33346
rect 14364 33282 14420 33294
rect 14252 33170 14308 33180
rect 14700 32900 14756 38612
rect 14812 38500 14868 38510
rect 14812 38050 14868 38444
rect 14812 37998 14814 38050
rect 14866 37998 14868 38050
rect 14812 37986 14868 37998
rect 14924 38388 14980 38398
rect 14924 37378 14980 38332
rect 15148 38276 15204 38286
rect 15036 38164 15092 38202
rect 15036 38098 15092 38108
rect 15036 37940 15092 37950
rect 15036 37846 15092 37884
rect 14924 37326 14926 37378
rect 14978 37326 14980 37378
rect 14924 37314 14980 37326
rect 14812 37266 14868 37278
rect 14812 37214 14814 37266
rect 14866 37214 14868 37266
rect 14812 36258 14868 37214
rect 14812 36206 14814 36258
rect 14866 36206 14868 36258
rect 14812 36194 14868 36206
rect 14924 36260 14980 36270
rect 14924 35698 14980 36204
rect 15036 35924 15092 35934
rect 15036 35830 15092 35868
rect 14924 35646 14926 35698
rect 14978 35646 14980 35698
rect 14924 35634 14980 35646
rect 15148 35810 15204 38220
rect 15372 37604 15428 37614
rect 15260 37268 15316 37278
rect 15260 37044 15316 37212
rect 15260 36978 15316 36988
rect 15148 35758 15150 35810
rect 15202 35758 15204 35810
rect 15148 35138 15204 35758
rect 15148 35086 15150 35138
rect 15202 35086 15204 35138
rect 15148 35074 15204 35086
rect 15260 36484 15316 36494
rect 15260 34916 15316 36428
rect 15036 34860 15316 34916
rect 13916 31778 14084 31780
rect 13916 31726 13918 31778
rect 13970 31726 14084 31778
rect 13916 31724 14084 31726
rect 14140 32844 14756 32900
rect 14812 34132 14868 34142
rect 14812 33458 14868 34076
rect 14812 33406 14814 33458
rect 14866 33406 14868 33458
rect 13916 31714 13972 31724
rect 13804 30942 13806 30994
rect 13858 30942 13860 30994
rect 13804 30930 13860 30942
rect 14140 31666 14196 32844
rect 14812 32788 14868 33406
rect 15036 33346 15092 34860
rect 15148 34692 15204 34702
rect 15148 34598 15204 34636
rect 15372 34244 15428 37548
rect 15596 37268 15652 38892
rect 15596 37202 15652 37212
rect 15820 37266 15876 40908
rect 15932 40898 15988 40908
rect 16044 40404 16100 40414
rect 15932 40290 15988 40302
rect 15932 40238 15934 40290
rect 15986 40238 15988 40290
rect 15932 38276 15988 40238
rect 16044 39058 16100 40348
rect 16156 39730 16212 41132
rect 16268 40516 16324 43596
rect 16604 43652 16660 45388
rect 16828 44100 16884 47516
rect 17276 47460 17332 47470
rect 16940 47458 17332 47460
rect 16940 47406 17278 47458
rect 17330 47406 17332 47458
rect 16940 47404 17332 47406
rect 16940 46898 16996 47404
rect 17276 47394 17332 47404
rect 16940 46846 16942 46898
rect 16994 46846 16996 46898
rect 16940 46834 16996 46846
rect 17388 46116 17444 47628
rect 17388 46050 17444 46060
rect 17388 45892 17444 45902
rect 17388 45798 17444 45836
rect 16940 45668 16996 45678
rect 16940 45330 16996 45612
rect 16940 45278 16942 45330
rect 16994 45278 16996 45330
rect 16940 45266 16996 45278
rect 17276 44100 17332 44110
rect 16828 44098 16996 44100
rect 16828 44046 16830 44098
rect 16882 44046 16996 44098
rect 16828 44044 16996 44046
rect 16828 44034 16884 44044
rect 16828 43876 16884 43886
rect 16828 43762 16884 43820
rect 16828 43710 16830 43762
rect 16882 43710 16884 43762
rect 16828 43698 16884 43710
rect 16604 43650 16772 43652
rect 16604 43598 16606 43650
rect 16658 43598 16772 43650
rect 16604 43596 16772 43598
rect 16604 43586 16660 43596
rect 16380 43540 16436 43550
rect 16380 43446 16436 43484
rect 16492 43426 16548 43438
rect 16492 43374 16494 43426
rect 16546 43374 16548 43426
rect 16380 43316 16436 43326
rect 16380 42532 16436 43260
rect 16492 42644 16548 43374
rect 16492 42578 16548 42588
rect 16380 42466 16436 42476
rect 16604 42532 16660 42542
rect 16492 41972 16548 41982
rect 16604 41972 16660 42476
rect 16492 41970 16660 41972
rect 16492 41918 16494 41970
rect 16546 41918 16660 41970
rect 16492 41916 16660 41918
rect 16492 41906 16548 41916
rect 16380 40964 16436 41002
rect 16380 40898 16436 40908
rect 16604 40852 16660 40862
rect 16268 40450 16324 40460
rect 16380 40740 16436 40750
rect 16380 40514 16436 40684
rect 16380 40462 16382 40514
rect 16434 40462 16436 40514
rect 16380 40450 16436 40462
rect 16492 40516 16548 40526
rect 16492 40422 16548 40460
rect 16604 40402 16660 40796
rect 16604 40350 16606 40402
rect 16658 40350 16660 40402
rect 16604 40338 16660 40350
rect 16716 39844 16772 43596
rect 16940 41858 16996 44044
rect 17276 44006 17332 44044
rect 17500 44100 17556 49196
rect 18060 49026 18116 49308
rect 18060 48974 18062 49026
rect 18114 48974 18116 49026
rect 18060 48962 18116 48974
rect 18172 49476 18228 49486
rect 18172 48916 18228 49420
rect 18172 48822 18228 48860
rect 17948 48356 18004 48366
rect 17948 48242 18004 48300
rect 18284 48356 18340 50372
rect 18396 49476 18452 50540
rect 18508 50036 18564 51548
rect 18620 51378 18676 51390
rect 18620 51326 18622 51378
rect 18674 51326 18676 51378
rect 18620 50260 18676 51326
rect 18732 50372 18788 52670
rect 19292 52612 19348 52622
rect 18844 51828 18900 51838
rect 18844 51602 18900 51772
rect 18844 51550 18846 51602
rect 18898 51550 18900 51602
rect 18844 51538 18900 51550
rect 19292 51492 19348 52556
rect 19404 52500 19460 52510
rect 19404 52274 19460 52444
rect 19404 52222 19406 52274
rect 19458 52222 19460 52274
rect 19404 52210 19460 52222
rect 19404 51492 19460 51502
rect 19292 51490 19460 51492
rect 19292 51438 19406 51490
rect 19458 51438 19460 51490
rect 19292 51436 19460 51438
rect 19404 51426 19460 51436
rect 18956 51268 19012 51278
rect 18956 51174 19012 51212
rect 18732 50278 18788 50316
rect 19180 50706 19236 50718
rect 19180 50654 19182 50706
rect 19234 50654 19236 50706
rect 18620 50194 18676 50204
rect 19068 50148 19124 50158
rect 19180 50148 19236 50654
rect 19516 50428 19572 52782
rect 19964 52722 20020 52734
rect 19964 52670 19966 52722
rect 20018 52670 20020 52722
rect 19964 52274 20020 52670
rect 19964 52222 19966 52274
rect 20018 52222 20020 52274
rect 19964 52210 20020 52222
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 20188 51604 20244 54684
rect 20300 54628 20356 55692
rect 20300 54562 20356 54572
rect 20524 54404 20580 57148
rect 20748 56642 20804 56654
rect 20748 56590 20750 56642
rect 20802 56590 20804 56642
rect 20636 55412 20692 55422
rect 20636 55318 20692 55356
rect 20748 54740 20804 56590
rect 20748 54674 20804 54684
rect 20300 54348 20580 54404
rect 20636 54404 20692 54414
rect 20636 54402 20804 54404
rect 20636 54350 20638 54402
rect 20690 54350 20804 54402
rect 20636 54348 20804 54350
rect 20300 53060 20356 54348
rect 20636 54338 20692 54348
rect 20524 53956 20580 53966
rect 20412 53844 20468 53854
rect 20412 53750 20468 53788
rect 20524 53842 20580 53900
rect 20524 53790 20526 53842
rect 20578 53790 20580 53842
rect 20524 53778 20580 53790
rect 20636 53506 20692 53518
rect 20636 53454 20638 53506
rect 20690 53454 20692 53506
rect 20636 53284 20692 53454
rect 20524 53228 20692 53284
rect 20524 53170 20580 53228
rect 20524 53118 20526 53170
rect 20578 53118 20580 53170
rect 20524 53106 20580 53118
rect 20412 53060 20468 53070
rect 20300 53058 20468 53060
rect 20300 53006 20414 53058
rect 20466 53006 20468 53058
rect 20300 53004 20468 53006
rect 20412 52994 20468 53004
rect 20636 53058 20692 53070
rect 20636 53006 20638 53058
rect 20690 53006 20692 53058
rect 20636 52948 20692 53006
rect 20636 52500 20692 52892
rect 20636 52434 20692 52444
rect 20524 52388 20580 52398
rect 20524 52274 20580 52332
rect 20524 52222 20526 52274
rect 20578 52222 20580 52274
rect 20524 52210 20580 52222
rect 20636 52164 20692 52174
rect 20076 51548 20244 51604
rect 20300 51940 20356 51950
rect 20076 51378 20132 51548
rect 20076 51326 20078 51378
rect 20130 51326 20132 51378
rect 19740 51268 19796 51278
rect 19796 51212 20020 51268
rect 19740 51174 19796 51212
rect 19964 50706 20020 51212
rect 20076 50932 20132 51326
rect 20076 50866 20132 50876
rect 19964 50654 19966 50706
rect 20018 50654 20020 50706
rect 19964 50642 20020 50654
rect 20300 50594 20356 51884
rect 20300 50542 20302 50594
rect 20354 50542 20356 50594
rect 20300 50428 20356 50542
rect 19516 50372 19684 50428
rect 20300 50372 20468 50428
rect 19124 50092 19236 50148
rect 19292 50148 19348 50158
rect 19068 50082 19124 50092
rect 19292 50036 19348 50092
rect 18508 49980 18788 50036
rect 18508 49812 18564 49822
rect 18508 49718 18564 49756
rect 18396 49410 18452 49420
rect 18396 49140 18452 49150
rect 18396 49046 18452 49084
rect 18396 48802 18452 48814
rect 18396 48750 18398 48802
rect 18450 48750 18452 48802
rect 18396 48580 18452 48750
rect 18396 48514 18452 48524
rect 18508 48804 18564 48814
rect 18732 48804 18788 49980
rect 18508 48802 18788 48804
rect 18508 48750 18510 48802
rect 18562 48750 18788 48802
rect 18508 48748 18788 48750
rect 19180 50034 19348 50036
rect 19180 49982 19294 50034
rect 19346 49982 19348 50034
rect 19180 49980 19348 49982
rect 18284 48290 18340 48300
rect 17948 48190 17950 48242
rect 18002 48190 18004 48242
rect 17836 48132 17892 48142
rect 17836 48038 17892 48076
rect 17612 47572 17668 47582
rect 17612 47478 17668 47516
rect 17948 47348 18004 48190
rect 18508 48244 18564 48748
rect 18508 48178 18564 48188
rect 19180 48468 19236 49980
rect 19292 49970 19348 49980
rect 19404 50036 19460 50046
rect 18172 48020 18228 48030
rect 18396 48020 18452 48030
rect 17724 47236 17780 47246
rect 17724 44324 17780 47180
rect 17836 46674 17892 46686
rect 17836 46622 17838 46674
rect 17890 46622 17892 46674
rect 17836 46564 17892 46622
rect 17836 46498 17892 46508
rect 17948 46340 18004 47292
rect 18060 47570 18116 47582
rect 18060 47518 18062 47570
rect 18114 47518 18116 47570
rect 18060 47012 18116 47518
rect 18172 47458 18228 47964
rect 18172 47406 18174 47458
rect 18226 47406 18228 47458
rect 18172 47394 18228 47406
rect 18284 48018 18452 48020
rect 18284 47966 18398 48018
rect 18450 47966 18452 48018
rect 18284 47964 18452 47966
rect 18060 46946 18116 46956
rect 17948 46274 18004 46284
rect 17836 46116 17892 46126
rect 17836 45332 17892 46060
rect 18172 45892 18228 45902
rect 18284 45892 18340 47964
rect 18396 47954 18452 47964
rect 18956 47572 19012 47582
rect 18508 47346 18564 47358
rect 18508 47294 18510 47346
rect 18562 47294 18564 47346
rect 18508 46786 18564 47294
rect 18508 46734 18510 46786
rect 18562 46734 18564 46786
rect 18508 46722 18564 46734
rect 18620 46452 18676 46462
rect 18172 45890 18340 45892
rect 18172 45838 18174 45890
rect 18226 45838 18340 45890
rect 18172 45836 18340 45838
rect 18508 46228 18564 46238
rect 18508 45890 18564 46172
rect 18508 45838 18510 45890
rect 18562 45838 18564 45890
rect 18172 45826 18228 45836
rect 18508 45826 18564 45838
rect 18284 45332 18340 45342
rect 17836 45276 18228 45332
rect 17836 45218 17892 45276
rect 17836 45166 17838 45218
rect 17890 45166 17892 45218
rect 17836 45154 17892 45166
rect 18060 45106 18116 45118
rect 18060 45054 18062 45106
rect 18114 45054 18116 45106
rect 17948 44436 18004 44446
rect 17724 44322 17892 44324
rect 17724 44270 17726 44322
rect 17778 44270 17892 44322
rect 17724 44268 17892 44270
rect 17724 44258 17780 44268
rect 17500 44034 17556 44044
rect 17052 43876 17108 43886
rect 17052 42756 17108 43820
rect 17724 43540 17780 43550
rect 17612 43538 17780 43540
rect 17612 43486 17726 43538
rect 17778 43486 17780 43538
rect 17612 43484 17780 43486
rect 17276 43316 17332 43326
rect 17052 42754 17220 42756
rect 17052 42702 17054 42754
rect 17106 42702 17220 42754
rect 17052 42700 17220 42702
rect 17052 42690 17108 42700
rect 16940 41806 16942 41858
rect 16994 41806 16996 41858
rect 16940 41636 16996 41806
rect 16940 41570 16996 41580
rect 16940 41076 16996 41086
rect 16940 40982 16996 41020
rect 16940 40740 16996 40750
rect 16940 40514 16996 40684
rect 16940 40462 16942 40514
rect 16994 40462 16996 40514
rect 16940 40450 16996 40462
rect 16604 39788 16772 39844
rect 16828 39844 16884 39854
rect 16156 39678 16158 39730
rect 16210 39678 16212 39730
rect 16156 39396 16212 39678
rect 16156 39330 16212 39340
rect 16268 39732 16324 39742
rect 16044 39006 16046 39058
rect 16098 39006 16100 39058
rect 16044 38500 16100 39006
rect 16268 39060 16324 39676
rect 16044 38434 16100 38444
rect 16156 38836 16212 38846
rect 15932 38210 15988 38220
rect 15820 37214 15822 37266
rect 15874 37214 15876 37266
rect 15820 37202 15876 37214
rect 15932 38050 15988 38062
rect 15932 37998 15934 38050
rect 15986 37998 15988 38050
rect 15484 36932 15540 36942
rect 15484 36482 15540 36876
rect 15484 36430 15486 36482
rect 15538 36430 15540 36482
rect 15484 36418 15540 36430
rect 15484 35140 15540 35150
rect 15484 35026 15540 35084
rect 15484 34974 15486 35026
rect 15538 34974 15540 35026
rect 15484 34962 15540 34974
rect 15708 35138 15764 35150
rect 15708 35086 15710 35138
rect 15762 35086 15764 35138
rect 15596 34244 15652 34254
rect 15372 34242 15652 34244
rect 15372 34190 15598 34242
rect 15650 34190 15652 34242
rect 15372 34188 15652 34190
rect 15596 34178 15652 34188
rect 15036 33294 15038 33346
rect 15090 33294 15092 33346
rect 14588 32732 14868 32788
rect 14924 33012 14980 33022
rect 14364 32676 14420 32686
rect 14364 32582 14420 32620
rect 14588 32674 14644 32732
rect 14588 32622 14590 32674
rect 14642 32622 14644 32674
rect 14588 32610 14644 32622
rect 14140 31614 14142 31666
rect 14194 31614 14196 31666
rect 13916 30882 13972 30894
rect 13916 30830 13918 30882
rect 13970 30830 13972 30882
rect 13692 30772 13748 30782
rect 13692 30210 13748 30716
rect 13692 30158 13694 30210
rect 13746 30158 13748 30210
rect 13692 30146 13748 30158
rect 13580 29922 13636 29932
rect 13468 26226 13524 26236
rect 13580 29428 13636 29438
rect 13244 24782 13246 24834
rect 13298 24782 13300 24834
rect 13244 24770 13300 24782
rect 13020 24052 13076 24062
rect 13020 23958 13076 23996
rect 13468 23492 13524 23502
rect 13468 23378 13524 23436
rect 13468 23326 13470 23378
rect 13522 23326 13524 23378
rect 13468 23314 13524 23326
rect 13580 23380 13636 29372
rect 13804 29428 13860 29438
rect 13804 29334 13860 29372
rect 13692 29316 13748 29326
rect 13692 28754 13748 29260
rect 13692 28702 13694 28754
rect 13746 28702 13748 28754
rect 13692 28532 13748 28702
rect 13692 28466 13748 28476
rect 13804 28420 13860 28430
rect 13692 28196 13748 28206
rect 13692 25620 13748 28140
rect 13804 28082 13860 28364
rect 13804 28030 13806 28082
rect 13858 28030 13860 28082
rect 13804 28018 13860 28030
rect 13916 27074 13972 30830
rect 14140 30324 14196 31614
rect 14252 32562 14308 32574
rect 14252 32510 14254 32562
rect 14306 32510 14308 32562
rect 14252 31556 14308 32510
rect 14700 32564 14756 32574
rect 14924 32564 14980 32956
rect 14700 32562 14980 32564
rect 14700 32510 14702 32562
rect 14754 32510 14980 32562
rect 14700 32508 14980 32510
rect 14700 32228 14756 32508
rect 14700 32162 14756 32172
rect 14924 32116 14980 32126
rect 14700 31780 14756 31790
rect 14588 31668 14644 31678
rect 14588 31574 14644 31612
rect 14252 31554 14532 31556
rect 14252 31502 14254 31554
rect 14306 31502 14532 31554
rect 14252 31500 14532 31502
rect 14252 31490 14308 31500
rect 14140 30258 14196 30268
rect 14364 30212 14420 30222
rect 14252 30210 14420 30212
rect 14252 30158 14366 30210
rect 14418 30158 14420 30210
rect 14252 30156 14420 30158
rect 14140 30098 14196 30110
rect 14140 30046 14142 30098
rect 14194 30046 14196 30098
rect 14028 29988 14084 29998
rect 14028 29538 14084 29932
rect 14140 29652 14196 30046
rect 14140 29586 14196 29596
rect 14252 29764 14308 30156
rect 14364 30146 14420 30156
rect 14028 29486 14030 29538
rect 14082 29486 14084 29538
rect 14028 29474 14084 29486
rect 14252 28980 14308 29708
rect 14364 29428 14420 29466
rect 14364 29362 14420 29372
rect 14364 29204 14420 29214
rect 14364 29110 14420 29148
rect 14252 28924 14420 28980
rect 14140 28644 14196 28654
rect 14140 28550 14196 28588
rect 14252 28308 14308 28318
rect 14252 28082 14308 28252
rect 14252 28030 14254 28082
rect 14306 28030 14308 28082
rect 14252 28018 14308 28030
rect 13916 27022 13918 27074
rect 13970 27022 13972 27074
rect 13916 26180 13972 27022
rect 14364 26852 14420 28924
rect 14476 28530 14532 31500
rect 14588 29650 14644 29662
rect 14588 29598 14590 29650
rect 14642 29598 14644 29650
rect 14588 28756 14644 29598
rect 14588 28690 14644 28700
rect 14476 28478 14478 28530
rect 14530 28478 14532 28530
rect 14476 28466 14532 28478
rect 14700 28420 14756 31724
rect 14812 30884 14868 30894
rect 14812 29204 14868 30828
rect 14924 29540 14980 32060
rect 15036 29876 15092 33294
rect 15148 34020 15204 34030
rect 15148 32004 15204 33964
rect 15260 33348 15316 33358
rect 15260 32004 15316 33292
rect 15372 32452 15428 32462
rect 15372 32450 15540 32452
rect 15372 32398 15374 32450
rect 15426 32398 15540 32450
rect 15372 32396 15540 32398
rect 15372 32386 15428 32396
rect 15484 32004 15540 32396
rect 15260 31948 15428 32004
rect 15148 31938 15204 31948
rect 15148 31778 15204 31790
rect 15148 31726 15150 31778
rect 15202 31726 15204 31778
rect 15148 31556 15204 31726
rect 15260 31780 15316 31790
rect 15260 31666 15316 31724
rect 15260 31614 15262 31666
rect 15314 31614 15316 31666
rect 15260 31602 15316 31614
rect 15148 31490 15204 31500
rect 15148 30996 15204 31006
rect 15148 30324 15204 30940
rect 15372 30994 15428 31948
rect 15708 31948 15764 35086
rect 15932 34916 15988 37998
rect 16156 37826 16212 38780
rect 16268 38274 16324 39004
rect 16268 38222 16270 38274
rect 16322 38222 16324 38274
rect 16268 38210 16324 38222
rect 16380 39284 16436 39294
rect 16380 38948 16436 39228
rect 16604 38948 16660 39788
rect 16716 39620 16772 39630
rect 16716 39526 16772 39564
rect 16828 39618 16884 39788
rect 17164 39732 17220 42700
rect 17276 42642 17332 43260
rect 17612 42980 17668 43484
rect 17724 43474 17780 43484
rect 17836 43092 17892 44268
rect 17948 43762 18004 44380
rect 17948 43710 17950 43762
rect 18002 43710 18004 43762
rect 17948 43540 18004 43710
rect 18060 43876 18116 45054
rect 18060 43650 18116 43820
rect 18060 43598 18062 43650
rect 18114 43598 18116 43650
rect 18060 43586 18116 43598
rect 18172 44322 18228 45276
rect 18284 45238 18340 45276
rect 18620 44884 18676 46396
rect 18620 44818 18676 44828
rect 18844 44994 18900 45006
rect 18844 44942 18846 44994
rect 18898 44942 18900 44994
rect 18172 44270 18174 44322
rect 18226 44270 18228 44322
rect 17948 43474 18004 43484
rect 17612 42914 17668 42924
rect 17724 43036 17892 43092
rect 17724 42756 17780 43036
rect 17500 42754 17780 42756
rect 17500 42702 17726 42754
rect 17778 42702 17780 42754
rect 17500 42700 17780 42702
rect 17276 42590 17278 42642
rect 17330 42590 17332 42642
rect 17276 42578 17332 42590
rect 17388 42644 17444 42654
rect 17388 42550 17444 42588
rect 17276 41860 17332 41870
rect 17276 40292 17332 41804
rect 17388 41410 17444 41422
rect 17388 41358 17390 41410
rect 17442 41358 17444 41410
rect 17388 41298 17444 41358
rect 17388 41246 17390 41298
rect 17442 41246 17444 41298
rect 17388 41234 17444 41246
rect 17388 40740 17444 40750
rect 17500 40740 17556 42700
rect 17724 42690 17780 42700
rect 17836 42866 17892 42878
rect 17836 42814 17838 42866
rect 17890 42814 17892 42866
rect 17836 42084 17892 42814
rect 17948 42532 18004 42542
rect 17948 42308 18004 42476
rect 18172 42420 18228 44270
rect 18284 44324 18340 44334
rect 18284 44230 18340 44268
rect 18396 44100 18452 44110
rect 18172 42308 18228 42364
rect 17948 42252 18228 42308
rect 18284 44098 18452 44100
rect 18284 44046 18398 44098
rect 18450 44046 18452 44098
rect 18284 44044 18452 44046
rect 17948 42194 18004 42252
rect 17948 42142 17950 42194
rect 18002 42142 18004 42194
rect 17948 42130 18004 42142
rect 17836 42018 17892 42028
rect 17612 41860 17668 41870
rect 17836 41860 17892 41870
rect 17668 41804 17780 41860
rect 17612 41794 17668 41804
rect 17724 41746 17780 41804
rect 17836 41766 17892 41804
rect 17724 41694 17726 41746
rect 17778 41694 17780 41746
rect 17724 41682 17780 41694
rect 17612 41410 17668 41422
rect 17612 41358 17614 41410
rect 17666 41358 17668 41410
rect 17612 41076 17668 41358
rect 17724 41412 17780 41422
rect 17724 41300 17780 41356
rect 17724 41298 18004 41300
rect 17724 41246 17726 41298
rect 17778 41246 18004 41298
rect 17724 41244 18004 41246
rect 17724 41234 17780 41244
rect 17612 41020 17780 41076
rect 17724 40852 17780 41020
rect 17444 40684 17556 40740
rect 17612 40796 17780 40852
rect 17836 40964 17892 40974
rect 17388 40674 17444 40684
rect 17276 40236 17444 40292
rect 17164 39666 17220 39676
rect 16828 39566 16830 39618
rect 16882 39566 16884 39618
rect 16716 39060 16772 39070
rect 16716 38966 16772 39004
rect 16828 39058 16884 39566
rect 17164 39508 17220 39518
rect 17164 39414 17220 39452
rect 17388 39506 17444 40236
rect 17500 40178 17556 40190
rect 17500 40126 17502 40178
rect 17554 40126 17556 40178
rect 17500 39620 17556 40126
rect 17612 39844 17668 40796
rect 17836 40740 17892 40908
rect 17724 40684 17892 40740
rect 17724 40626 17780 40684
rect 17724 40574 17726 40626
rect 17778 40574 17780 40626
rect 17724 40562 17780 40574
rect 17612 39778 17668 39788
rect 17948 40180 18004 41244
rect 18060 41188 18116 41198
rect 18060 40402 18116 41132
rect 18172 40962 18228 40974
rect 18172 40910 18174 40962
rect 18226 40910 18228 40962
rect 18172 40628 18228 40910
rect 18172 40562 18228 40572
rect 18060 40350 18062 40402
rect 18114 40350 18116 40402
rect 18060 40338 18116 40350
rect 18284 40404 18340 44044
rect 18396 44034 18452 44044
rect 18844 43652 18900 44942
rect 18956 44100 19012 47516
rect 19180 44996 19236 48412
rect 19292 48468 19348 48478
rect 19404 48468 19460 49980
rect 19628 49028 19684 50372
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 19852 49924 19908 49934
rect 19852 49830 19908 49868
rect 19292 48466 19460 48468
rect 19292 48414 19294 48466
rect 19346 48414 19460 48466
rect 19292 48412 19460 48414
rect 19516 49026 19684 49028
rect 19516 48974 19630 49026
rect 19682 48974 19684 49026
rect 19516 48972 19684 48974
rect 19292 48402 19348 48412
rect 19292 47348 19348 47358
rect 19292 47254 19348 47292
rect 19292 44996 19348 45006
rect 19180 44994 19348 44996
rect 19180 44942 19294 44994
rect 19346 44942 19348 44994
rect 19180 44940 19348 44942
rect 19292 44772 19348 44940
rect 19292 44706 19348 44716
rect 19292 44436 19348 44446
rect 19516 44436 19572 48972
rect 19628 48962 19684 48972
rect 20076 49028 20132 49038
rect 20076 48934 20132 48972
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 20188 48242 20244 48254
rect 20188 48190 20190 48242
rect 20242 48190 20244 48242
rect 19628 48132 19684 48142
rect 19628 47236 19684 48076
rect 19852 47572 19908 47582
rect 19852 47458 19908 47516
rect 20076 47572 20132 47582
rect 20188 47572 20244 48190
rect 20412 47796 20468 50372
rect 20524 49810 20580 49822
rect 20524 49758 20526 49810
rect 20578 49758 20580 49810
rect 20524 49140 20580 49758
rect 20524 49074 20580 49084
rect 20412 47730 20468 47740
rect 20636 48244 20692 52108
rect 20748 49812 20804 54348
rect 20860 52948 20916 57484
rect 20972 57474 21028 57484
rect 20972 56644 21028 56654
rect 20972 56306 21028 56588
rect 20972 56254 20974 56306
rect 21026 56254 21028 56306
rect 20972 55076 21028 56254
rect 20972 55010 21028 55020
rect 20860 52882 20916 52892
rect 21084 54402 21140 54414
rect 21084 54350 21086 54402
rect 21138 54350 21140 54402
rect 20860 52164 20916 52174
rect 20860 52070 20916 52108
rect 21084 52052 21140 54350
rect 21196 54180 21252 59500
rect 21308 55748 21364 59724
rect 21420 59714 21476 59724
rect 21868 59778 21924 59790
rect 21868 59726 21870 59778
rect 21922 59726 21924 59778
rect 21756 59218 21812 59230
rect 21756 59166 21758 59218
rect 21810 59166 21812 59218
rect 21756 58772 21812 59166
rect 21868 58884 21924 59726
rect 21868 58818 21924 58828
rect 21756 58706 21812 58716
rect 21868 58212 21924 58222
rect 21420 57540 21476 57550
rect 21420 57538 21588 57540
rect 21420 57486 21422 57538
rect 21474 57486 21588 57538
rect 21420 57484 21588 57486
rect 21420 57474 21476 57484
rect 21420 56084 21476 56094
rect 21420 55990 21476 56028
rect 21308 55682 21364 55692
rect 21532 55468 21588 57484
rect 21532 55412 21812 55468
rect 21196 54114 21252 54124
rect 21644 55076 21700 55086
rect 21308 53340 21588 53396
rect 21084 51986 21140 51996
rect 21196 53060 21252 53070
rect 21196 51602 21252 53004
rect 21196 51550 21198 51602
rect 21250 51550 21252 51602
rect 21196 51154 21252 51550
rect 21196 51102 21198 51154
rect 21250 51102 21252 51154
rect 21196 51090 21252 51102
rect 20860 50482 20916 50494
rect 20860 50430 20862 50482
rect 20914 50430 20916 50482
rect 20860 50148 20916 50430
rect 20860 50082 20916 50092
rect 20972 50372 21028 50382
rect 20748 49680 20804 49756
rect 20860 49140 20916 49150
rect 20860 49046 20916 49084
rect 20860 48356 20916 48366
rect 20860 48262 20916 48300
rect 20748 48244 20804 48254
rect 20636 48242 20804 48244
rect 20636 48190 20750 48242
rect 20802 48190 20804 48242
rect 20636 48188 20804 48190
rect 20188 47516 20580 47572
rect 20076 47478 20132 47516
rect 19852 47406 19854 47458
rect 19906 47406 19908 47458
rect 19852 47394 19908 47406
rect 20188 47348 20244 47358
rect 20188 47346 20468 47348
rect 20188 47294 20190 47346
rect 20242 47294 20468 47346
rect 20188 47292 20468 47294
rect 20188 47282 20244 47292
rect 20076 47236 20132 47246
rect 19628 47234 20132 47236
rect 19628 47182 20078 47234
rect 20130 47182 20132 47234
rect 19628 47180 20132 47182
rect 19628 46004 19684 47180
rect 20076 47170 20132 47180
rect 20188 47124 20244 47134
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 19628 45332 19684 45948
rect 19852 46674 19908 46686
rect 19852 46622 19854 46674
rect 19906 46622 19908 46674
rect 19852 45666 19908 46622
rect 19852 45614 19854 45666
rect 19906 45614 19908 45666
rect 19852 45602 19908 45614
rect 20188 45778 20244 47068
rect 20412 47012 20468 47292
rect 20188 45726 20190 45778
rect 20242 45726 20244 45778
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 19628 45276 19796 45332
rect 19740 44436 19796 45276
rect 20188 45108 20244 45726
rect 20300 46956 20412 47012
rect 20300 45892 20356 46956
rect 20412 46880 20468 46956
rect 20412 46564 20468 46574
rect 20412 46470 20468 46508
rect 20300 45444 20356 45836
rect 20524 45890 20580 47516
rect 20636 47458 20692 48188
rect 20748 48178 20804 48188
rect 20636 47406 20638 47458
rect 20690 47406 20692 47458
rect 20636 47124 20692 47406
rect 20636 47058 20692 47068
rect 20860 47572 20916 47582
rect 20524 45838 20526 45890
rect 20578 45838 20580 45890
rect 20412 45444 20468 45454
rect 20300 45388 20412 45444
rect 20188 45014 20244 45052
rect 19516 44380 19684 44436
rect 19068 44324 19124 44334
rect 19068 44230 19124 44268
rect 19180 44212 19236 44222
rect 19180 44118 19236 44156
rect 18956 44044 19124 44100
rect 18844 43586 18900 43596
rect 18732 43538 18788 43550
rect 18732 43486 18734 43538
rect 18786 43486 18788 43538
rect 18732 43428 18788 43486
rect 18956 43540 19012 43550
rect 18956 43446 19012 43484
rect 18732 43362 18788 43372
rect 18844 43426 18900 43438
rect 18844 43374 18846 43426
rect 18898 43374 18900 43426
rect 18396 42868 18452 42878
rect 18396 42774 18452 42812
rect 18732 42866 18788 42878
rect 18732 42814 18734 42866
rect 18786 42814 18788 42866
rect 18732 42756 18788 42814
rect 18732 42690 18788 42700
rect 18844 42644 18900 43374
rect 19068 42980 19124 44044
rect 19180 43426 19236 43438
rect 19180 43374 19182 43426
rect 19234 43374 19236 43426
rect 19180 43316 19236 43374
rect 19292 43428 19348 44380
rect 19516 44210 19572 44222
rect 19516 44158 19518 44210
rect 19570 44158 19572 44210
rect 19404 44098 19460 44110
rect 19404 44046 19406 44098
rect 19458 44046 19460 44098
rect 19404 43652 19460 44046
rect 19404 43586 19460 43596
rect 19516 44100 19572 44158
rect 19404 43428 19460 43438
rect 19292 43426 19460 43428
rect 19292 43374 19406 43426
rect 19458 43374 19460 43426
rect 19292 43372 19460 43374
rect 19404 43362 19460 43372
rect 19180 43250 19236 43260
rect 19068 42914 19124 42924
rect 19516 42868 19572 44044
rect 19628 43540 19684 44380
rect 19740 44370 19796 44380
rect 20300 44436 20356 44446
rect 20300 44210 20356 44380
rect 20300 44158 20302 44210
rect 20354 44158 20356 44210
rect 20300 44146 20356 44158
rect 20412 44210 20468 45388
rect 20524 45332 20580 45838
rect 20860 45668 20916 47516
rect 20524 45266 20580 45276
rect 20636 45612 20916 45668
rect 20412 44158 20414 44210
rect 20466 44158 20468 44210
rect 20412 44146 20468 44158
rect 20524 44210 20580 44222
rect 20524 44158 20526 44210
rect 20578 44158 20580 44210
rect 20076 44100 20132 44110
rect 20076 44098 20244 44100
rect 20076 44046 20078 44098
rect 20130 44046 20244 44098
rect 20076 44044 20244 44046
rect 20076 44034 20132 44044
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 20188 43764 20244 44044
rect 19628 43474 19684 43484
rect 19740 43708 20244 43764
rect 20412 43764 20468 43774
rect 19628 43316 19684 43326
rect 19740 43316 19796 43708
rect 19628 43314 19796 43316
rect 19628 43262 19630 43314
rect 19682 43262 19796 43314
rect 19628 43260 19796 43262
rect 20300 43540 20356 43550
rect 19628 42980 19684 43260
rect 19628 42914 19684 42924
rect 19516 42802 19572 42812
rect 19964 42644 20020 42654
rect 18844 42588 19460 42644
rect 18620 42532 18676 42542
rect 18620 42438 18676 42476
rect 18284 40338 18340 40348
rect 18396 42420 18452 42430
rect 18172 40290 18228 40302
rect 18172 40238 18174 40290
rect 18226 40238 18228 40290
rect 18172 40180 18228 40238
rect 18396 40180 18452 42364
rect 19180 42420 19236 42430
rect 18844 41858 18900 41870
rect 18844 41806 18846 41858
rect 18898 41806 18900 41858
rect 18620 41300 18676 41310
rect 18620 41206 18676 41244
rect 18732 41076 18788 41086
rect 18732 40852 18788 41020
rect 18732 40626 18788 40796
rect 18732 40574 18734 40626
rect 18786 40574 18788 40626
rect 18732 40562 18788 40574
rect 18508 40404 18564 40414
rect 18508 40310 18564 40348
rect 18844 40404 18900 41806
rect 19180 41300 19236 42364
rect 19404 42196 19460 42588
rect 19964 42550 20020 42588
rect 19516 42530 19572 42542
rect 19516 42478 19518 42530
rect 19570 42478 19572 42530
rect 19516 42420 19572 42478
rect 19516 42354 19572 42364
rect 19628 42532 19684 42542
rect 20300 42532 20356 43484
rect 20412 43538 20468 43708
rect 20412 43486 20414 43538
rect 20466 43486 20468 43538
rect 20412 43474 20468 43486
rect 20524 43316 20580 44158
rect 20524 43250 20580 43260
rect 20412 42532 20468 42542
rect 20300 42530 20468 42532
rect 20300 42478 20414 42530
rect 20466 42478 20468 42530
rect 20300 42476 20468 42478
rect 19516 42196 19572 42206
rect 19404 42194 19572 42196
rect 19404 42142 19518 42194
rect 19570 42142 19572 42194
rect 19404 42140 19572 42142
rect 19516 42130 19572 42140
rect 19628 42194 19684 42476
rect 20412 42420 20468 42476
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20412 42354 20468 42364
rect 19836 42298 20100 42308
rect 20636 42196 20692 45612
rect 20860 45444 20916 45454
rect 20860 45106 20916 45388
rect 20972 45218 21028 50316
rect 21308 50036 21364 53340
rect 21308 49970 21364 49980
rect 21420 53172 21476 53182
rect 21084 48468 21140 48478
rect 21084 48374 21140 48412
rect 21420 48468 21476 53116
rect 21532 53170 21588 53340
rect 21532 53118 21534 53170
rect 21586 53118 21588 53170
rect 21532 53106 21588 53118
rect 21644 53060 21700 55020
rect 21644 52994 21700 53004
rect 21756 55074 21812 55412
rect 21756 55022 21758 55074
rect 21810 55022 21812 55074
rect 21756 52612 21812 55022
rect 21868 55300 21924 58156
rect 21980 57652 22036 60174
rect 22540 60228 22596 60238
rect 22876 60228 22932 60238
rect 22540 60226 22932 60228
rect 22540 60174 22542 60226
rect 22594 60174 22878 60226
rect 22930 60174 22932 60226
rect 22540 60172 22932 60174
rect 22540 60162 22596 60172
rect 22876 60162 22932 60172
rect 23324 60002 23380 60014
rect 23324 59950 23326 60002
rect 23378 59950 23380 60002
rect 22764 59890 22820 59902
rect 22764 59838 22766 59890
rect 22818 59838 22820 59890
rect 22316 59780 22372 59790
rect 22316 59778 22596 59780
rect 22316 59726 22318 59778
rect 22370 59726 22596 59778
rect 22316 59724 22596 59726
rect 22316 59714 22372 59724
rect 22092 59106 22148 59118
rect 22092 59054 22094 59106
rect 22146 59054 22148 59106
rect 22092 58660 22148 59054
rect 22428 58994 22484 59006
rect 22428 58942 22430 58994
rect 22482 58942 22484 58994
rect 22092 58546 22148 58604
rect 22092 58494 22094 58546
rect 22146 58494 22148 58546
rect 22092 58482 22148 58494
rect 22316 58772 22372 58782
rect 22316 58434 22372 58716
rect 22316 58382 22318 58434
rect 22370 58382 22372 58434
rect 22316 58370 22372 58382
rect 21980 57650 22148 57652
rect 21980 57598 21982 57650
rect 22034 57598 22148 57650
rect 21980 57596 22148 57598
rect 21980 57586 22036 57596
rect 22092 57204 22148 57596
rect 22204 57428 22260 57438
rect 22204 57426 22372 57428
rect 22204 57374 22206 57426
rect 22258 57374 22372 57426
rect 22204 57372 22372 57374
rect 22204 57362 22260 57372
rect 22092 57148 22260 57204
rect 22092 56980 22148 56990
rect 22092 56754 22148 56924
rect 22204 56866 22260 57148
rect 22204 56814 22206 56866
rect 22258 56814 22260 56866
rect 22204 56802 22260 56814
rect 22092 56702 22094 56754
rect 22146 56702 22148 56754
rect 21980 56196 22036 56206
rect 21980 56082 22036 56140
rect 21980 56030 21982 56082
rect 22034 56030 22036 56082
rect 21980 55972 22036 56030
rect 22092 56084 22148 56702
rect 22316 56756 22372 57372
rect 22316 56662 22372 56700
rect 22428 56532 22484 58942
rect 22540 57764 22596 59724
rect 22764 58660 22820 59838
rect 22988 59890 23044 59902
rect 22988 59838 22990 59890
rect 23042 59838 23044 59890
rect 22988 59220 23044 59838
rect 23324 59668 23380 59950
rect 23324 59602 23380 59612
rect 23548 60002 23604 60014
rect 23548 59950 23550 60002
rect 23602 59950 23604 60002
rect 23548 59556 23604 59950
rect 24220 59778 24276 59790
rect 24220 59726 24222 59778
rect 24274 59726 24276 59778
rect 23548 59490 23604 59500
rect 24108 59668 24164 59678
rect 22988 59154 23044 59164
rect 23884 59220 23940 59230
rect 23884 59126 23940 59164
rect 24108 59218 24164 59612
rect 24108 59166 24110 59218
rect 24162 59166 24164 59218
rect 24108 59154 24164 59166
rect 23548 58994 23604 59006
rect 23548 58942 23550 58994
rect 23602 58942 23604 58994
rect 23548 58772 23604 58942
rect 23548 58706 23604 58716
rect 22764 58594 22820 58604
rect 23772 58434 23828 58446
rect 23772 58382 23774 58434
rect 23826 58382 23828 58434
rect 22876 58324 22932 58334
rect 23436 58324 23492 58334
rect 22876 58322 23492 58324
rect 22876 58270 22878 58322
rect 22930 58270 23438 58322
rect 23490 58270 23492 58322
rect 22876 58268 23492 58270
rect 22876 58258 22932 58268
rect 22540 57698 22596 57708
rect 23100 57762 23156 58268
rect 23436 58258 23492 58268
rect 23100 57710 23102 57762
rect 23154 57710 23156 57762
rect 23100 57698 23156 57710
rect 23548 58210 23604 58222
rect 23548 58158 23550 58210
rect 23602 58158 23604 58210
rect 23436 57650 23492 57662
rect 23436 57598 23438 57650
rect 23490 57598 23492 57650
rect 23212 57538 23268 57550
rect 23212 57486 23214 57538
rect 23266 57486 23268 57538
rect 22540 57428 22596 57438
rect 22540 57426 22708 57428
rect 22540 57374 22542 57426
rect 22594 57374 22708 57426
rect 22540 57372 22708 57374
rect 22540 57362 22596 57372
rect 22092 56018 22148 56028
rect 22316 56476 22484 56532
rect 22316 56082 22372 56476
rect 22540 56420 22596 56430
rect 22540 56306 22596 56364
rect 22540 56254 22542 56306
rect 22594 56254 22596 56306
rect 22540 56242 22596 56254
rect 22316 56030 22318 56082
rect 22370 56030 22372 56082
rect 22316 56018 22372 56030
rect 22428 56084 22484 56094
rect 21980 55906 22036 55916
rect 21868 54738 21924 55244
rect 22204 55074 22260 55086
rect 22204 55022 22206 55074
rect 22258 55022 22260 55074
rect 22204 54964 22260 55022
rect 22204 54898 22260 54908
rect 21868 54686 21870 54738
rect 21922 54686 21924 54738
rect 21868 54674 21924 54686
rect 22092 54404 22148 54414
rect 21980 53508 22036 53518
rect 21756 52546 21812 52556
rect 21868 53506 22036 53508
rect 21868 53454 21982 53506
rect 22034 53454 22036 53506
rect 21868 53452 22036 53454
rect 21532 52162 21588 52174
rect 21532 52110 21534 52162
rect 21586 52110 21588 52162
rect 21532 51716 21588 52110
rect 21868 52164 21924 53452
rect 21980 53442 22036 53452
rect 21980 53060 22036 53070
rect 21980 52966 22036 53004
rect 22092 52276 22148 54348
rect 22316 54402 22372 54414
rect 22316 54350 22318 54402
rect 22370 54350 22372 54402
rect 22316 53844 22372 54350
rect 22316 53778 22372 53788
rect 22428 53732 22484 56028
rect 22652 56082 22708 57372
rect 22764 57092 22820 57102
rect 22764 56998 22820 57036
rect 23212 56308 23268 57486
rect 23436 57540 23492 57598
rect 23436 57474 23492 57484
rect 23548 57090 23604 58158
rect 23548 57038 23550 57090
rect 23602 57038 23604 57090
rect 23548 57026 23604 57038
rect 23660 57650 23716 57662
rect 23660 57598 23662 57650
rect 23714 57598 23716 57650
rect 23660 57092 23716 57598
rect 23772 57540 23828 58382
rect 23772 57474 23828 57484
rect 24108 57540 24164 57550
rect 24220 57540 24276 59726
rect 24556 59778 24612 59790
rect 24556 59726 24558 59778
rect 24610 59726 24612 59778
rect 24556 59556 24612 59726
rect 24332 59500 24556 59556
rect 24332 59218 24388 59500
rect 24556 59490 24612 59500
rect 24668 59780 24724 59790
rect 24332 59166 24334 59218
rect 24386 59166 24388 59218
rect 24332 59154 24388 59166
rect 24556 58548 24612 58558
rect 24556 58454 24612 58492
rect 24444 58324 24500 58334
rect 24444 58230 24500 58268
rect 24164 57484 24276 57540
rect 24556 57538 24612 57550
rect 24556 57486 24558 57538
rect 24610 57486 24612 57538
rect 24108 57446 24164 57484
rect 24556 57204 24612 57486
rect 24108 57148 24612 57204
rect 23660 57026 23716 57036
rect 23996 57092 24052 57102
rect 23996 56998 24052 57036
rect 24108 56980 24164 57148
rect 24668 57092 24724 59724
rect 25228 59778 25284 59790
rect 25228 59726 25230 59778
rect 25282 59726 25284 59778
rect 25228 59668 25284 59726
rect 25228 59602 25284 59612
rect 24892 59556 24948 59566
rect 24892 59442 24948 59500
rect 24892 59390 24894 59442
rect 24946 59390 24948 59442
rect 24892 59378 24948 59390
rect 24780 58436 24836 58446
rect 24780 58342 24836 58380
rect 24108 56914 24164 56924
rect 24220 57036 24724 57092
rect 24780 57540 24836 57550
rect 23324 56866 23380 56878
rect 23324 56814 23326 56866
rect 23378 56814 23380 56866
rect 23324 56420 23380 56814
rect 23772 56868 23828 56878
rect 23772 56774 23828 56812
rect 23324 56354 23380 56364
rect 24108 56754 24164 56766
rect 24108 56702 24110 56754
rect 24162 56702 24164 56754
rect 24108 56420 24164 56702
rect 24108 56354 24164 56364
rect 23212 56242 23268 56252
rect 23660 56308 23716 56318
rect 23660 56214 23716 56252
rect 22652 56030 22654 56082
rect 22706 56030 22708 56082
rect 22652 55524 22708 56030
rect 23884 56082 23940 56094
rect 23884 56030 23886 56082
rect 23938 56030 23940 56082
rect 23772 55970 23828 55982
rect 23772 55918 23774 55970
rect 23826 55918 23828 55970
rect 23324 55636 23380 55646
rect 22988 55524 23044 55534
rect 22652 55522 23044 55524
rect 22652 55470 22990 55522
rect 23042 55470 23044 55522
rect 22652 55468 23044 55470
rect 22988 55458 23044 55468
rect 23324 55410 23380 55580
rect 23772 55524 23828 55918
rect 23884 55636 23940 56030
rect 23884 55570 23940 55580
rect 23996 55860 24052 55870
rect 23772 55458 23828 55468
rect 23324 55358 23326 55410
rect 23378 55358 23380 55410
rect 23324 55346 23380 55358
rect 22428 53638 22484 53676
rect 22540 55300 22596 55310
rect 22428 53172 22484 53182
rect 22540 53172 22596 55244
rect 23212 55074 23268 55086
rect 23772 55076 23828 55086
rect 23212 55022 23214 55074
rect 23266 55022 23268 55074
rect 22428 53170 22540 53172
rect 22428 53118 22430 53170
rect 22482 53118 22540 53170
rect 22428 53116 22540 53118
rect 22428 53106 22484 53116
rect 22540 53106 22596 53116
rect 22652 54964 22708 54974
rect 22652 53508 22708 54908
rect 22764 54740 22820 54750
rect 22764 54646 22820 54684
rect 23212 53732 23268 55022
rect 23548 55074 23828 55076
rect 23548 55022 23774 55074
rect 23826 55022 23828 55074
rect 23548 55020 23828 55022
rect 23324 54402 23380 54414
rect 23324 54350 23326 54402
rect 23378 54350 23380 54402
rect 23324 53956 23380 54350
rect 23324 53890 23380 53900
rect 23548 53844 23604 55020
rect 23772 55010 23828 55020
rect 23996 54738 24052 55804
rect 24220 55300 24276 57036
rect 24556 56866 24612 56878
rect 24556 56814 24558 56866
rect 24610 56814 24612 56866
rect 24332 56084 24388 56094
rect 24556 56084 24612 56814
rect 24332 56082 24612 56084
rect 24332 56030 24334 56082
rect 24386 56030 24612 56082
rect 24332 56028 24612 56030
rect 24332 56018 24388 56028
rect 23996 54686 23998 54738
rect 24050 54686 24052 54738
rect 23996 54674 24052 54686
rect 24108 55244 24276 55300
rect 23212 53666 23268 53676
rect 23436 53788 23604 53844
rect 22988 53620 23044 53630
rect 22988 53526 23044 53564
rect 23436 53620 23492 53788
rect 23660 53732 23716 53742
rect 22204 52946 22260 52958
rect 22204 52894 22206 52946
rect 22258 52894 22260 52946
rect 22204 52612 22260 52894
rect 22540 52948 22596 52958
rect 22540 52854 22596 52892
rect 22428 52836 22484 52846
rect 22428 52742 22484 52780
rect 22204 52546 22260 52556
rect 22652 52276 22708 53452
rect 22764 53506 22820 53518
rect 22764 53454 22766 53506
rect 22818 53454 22820 53506
rect 22764 53284 22820 53454
rect 22876 53508 22932 53518
rect 22876 53414 22932 53452
rect 22764 53218 22820 53228
rect 22876 53172 22932 53182
rect 22764 52276 22820 52286
rect 22092 52274 22484 52276
rect 22092 52222 22094 52274
rect 22146 52222 22484 52274
rect 22092 52220 22484 52222
rect 22652 52274 22820 52276
rect 22652 52222 22766 52274
rect 22818 52222 22820 52274
rect 22652 52220 22820 52222
rect 22092 52210 22148 52220
rect 21756 52052 21812 52062
rect 21532 51650 21588 51660
rect 21644 51940 21700 51950
rect 21532 51492 21588 51502
rect 21532 48692 21588 51436
rect 21644 51266 21700 51884
rect 21644 51214 21646 51266
rect 21698 51214 21700 51266
rect 21644 49924 21700 51214
rect 21644 49858 21700 49868
rect 21644 48916 21700 48926
rect 21644 48822 21700 48860
rect 21756 48914 21812 51996
rect 21868 51604 21924 52108
rect 22428 51940 22484 52220
rect 22764 52210 22820 52220
rect 22540 52164 22596 52174
rect 22540 52070 22596 52108
rect 22428 51884 22708 51940
rect 22092 51604 22148 51614
rect 21868 51602 22148 51604
rect 21868 51550 22094 51602
rect 22146 51550 22148 51602
rect 21868 51548 22148 51550
rect 21868 50818 21924 50830
rect 21868 50766 21870 50818
rect 21922 50766 21924 50818
rect 21868 50706 21924 50766
rect 21868 50654 21870 50706
rect 21922 50654 21924 50706
rect 21868 50642 21924 50654
rect 22092 50428 22148 51548
rect 22204 51156 22260 51166
rect 22204 51154 22484 51156
rect 22204 51102 22206 51154
rect 22258 51102 22484 51154
rect 22204 51100 22484 51102
rect 22204 51090 22260 51100
rect 22316 50708 22372 50718
rect 22092 50372 22260 50428
rect 22204 50260 22260 50372
rect 22204 50194 22260 50204
rect 22092 49924 22148 49934
rect 21980 49028 22036 49038
rect 21980 48934 22036 48972
rect 21756 48862 21758 48914
rect 21810 48862 21812 48914
rect 21756 48850 21812 48862
rect 21532 48636 21812 48692
rect 21420 48402 21476 48412
rect 21308 48356 21364 48366
rect 21308 47068 21364 48300
rect 21532 48354 21588 48366
rect 21532 48302 21534 48354
rect 21586 48302 21588 48354
rect 21532 47124 21588 48302
rect 21756 48242 21812 48636
rect 21756 48190 21758 48242
rect 21810 48190 21812 48242
rect 21308 47012 21476 47068
rect 21532 47058 21588 47068
rect 21644 47234 21700 47246
rect 21644 47182 21646 47234
rect 21698 47182 21700 47234
rect 21196 46786 21252 46798
rect 21196 46734 21198 46786
rect 21250 46734 21252 46786
rect 21196 45556 21252 46734
rect 21308 46674 21364 46686
rect 21308 46622 21310 46674
rect 21362 46622 21364 46674
rect 21308 45780 21364 46622
rect 21308 45714 21364 45724
rect 21420 45668 21476 47012
rect 21644 46452 21700 47182
rect 21644 46386 21700 46396
rect 21532 45668 21588 45678
rect 21420 45612 21532 45668
rect 21532 45574 21588 45612
rect 21196 45500 21364 45556
rect 20972 45166 20974 45218
rect 21026 45166 21028 45218
rect 20972 45154 21028 45166
rect 20860 45054 20862 45106
rect 20914 45054 20916 45106
rect 20860 45042 20916 45054
rect 21308 44772 21364 45500
rect 21644 45220 21700 45230
rect 20860 44434 20916 44446
rect 20860 44382 20862 44434
rect 20914 44382 20916 44434
rect 19628 42142 19630 42194
rect 19682 42142 19684 42194
rect 19628 42130 19684 42142
rect 20188 42140 20692 42196
rect 20748 44324 20804 44334
rect 19292 41970 19348 41982
rect 19292 41918 19294 41970
rect 19346 41918 19348 41970
rect 19292 41748 19348 41918
rect 19740 41970 19796 41982
rect 19740 41918 19742 41970
rect 19794 41918 19796 41970
rect 19740 41860 19796 41918
rect 19740 41794 19796 41804
rect 19852 41970 19908 41982
rect 19852 41918 19854 41970
rect 19906 41918 19908 41970
rect 19292 41682 19348 41692
rect 19180 41234 19236 41244
rect 19292 41524 19348 41534
rect 19068 41188 19124 41198
rect 19068 40628 19124 41132
rect 19292 41186 19348 41468
rect 19292 41134 19294 41186
rect 19346 41134 19348 41186
rect 19292 41122 19348 41134
rect 19404 41412 19460 41422
rect 19404 41186 19460 41356
rect 19628 41300 19684 41310
rect 19852 41300 19908 41918
rect 19628 41298 19908 41300
rect 19628 41246 19630 41298
rect 19682 41246 19908 41298
rect 19628 41244 19908 41246
rect 20188 41298 20244 42140
rect 20748 41972 20804 44268
rect 20860 43650 20916 44382
rect 20860 43598 20862 43650
rect 20914 43598 20916 43650
rect 20860 43586 20916 43598
rect 21196 43652 21252 43662
rect 21084 43428 21140 43438
rect 21084 43334 21140 43372
rect 21196 43426 21252 43596
rect 21308 43540 21364 44716
rect 21308 43474 21364 43484
rect 21532 44994 21588 45006
rect 21532 44942 21534 44994
rect 21586 44942 21588 44994
rect 21196 43374 21198 43426
rect 21250 43374 21252 43426
rect 21196 43362 21252 43374
rect 21420 43316 21476 43326
rect 20860 42530 20916 42542
rect 20860 42478 20862 42530
rect 20914 42478 20916 42530
rect 20860 42308 20916 42478
rect 20860 42242 20916 42252
rect 20860 41972 20916 41982
rect 21084 41972 21140 41982
rect 20748 41970 20916 41972
rect 20748 41918 20862 41970
rect 20914 41918 20916 41970
rect 20748 41916 20916 41918
rect 20860 41906 20916 41916
rect 20972 41916 21084 41972
rect 20524 41748 20580 41758
rect 20524 41654 20580 41692
rect 20188 41246 20190 41298
rect 20242 41246 20244 41298
rect 19628 41234 19684 41244
rect 19404 41134 19406 41186
rect 19458 41134 19460 41186
rect 19404 41122 19460 41134
rect 19740 41076 19796 41086
rect 19628 41074 19796 41076
rect 19628 41022 19742 41074
rect 19794 41022 19796 41074
rect 19628 41020 19796 41022
rect 19628 40852 19684 41020
rect 19740 41010 19796 41020
rect 19628 40786 19684 40796
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19180 40628 19236 40638
rect 19628 40628 19684 40638
rect 19068 40626 19348 40628
rect 19068 40574 19182 40626
rect 19234 40574 19348 40626
rect 19068 40572 19348 40574
rect 19180 40562 19236 40572
rect 18620 40292 18676 40302
rect 18620 40198 18676 40236
rect 18172 40124 18452 40180
rect 17612 39620 17668 39630
rect 17500 39618 17892 39620
rect 17500 39566 17614 39618
rect 17666 39566 17892 39618
rect 17500 39564 17892 39566
rect 17612 39554 17668 39564
rect 17388 39454 17390 39506
rect 17442 39454 17444 39506
rect 16828 39006 16830 39058
rect 16882 39006 16884 39058
rect 16828 38994 16884 39006
rect 16940 39284 16996 39294
rect 16380 38892 16660 38948
rect 16156 37774 16158 37826
rect 16210 37774 16212 37826
rect 16044 35812 16100 35822
rect 16044 35718 16100 35756
rect 16044 35028 16100 35038
rect 16044 34934 16100 34972
rect 15932 34850 15988 34860
rect 15820 34132 15876 34142
rect 15820 34038 15876 34076
rect 16044 34130 16100 34142
rect 16044 34078 16046 34130
rect 16098 34078 16100 34130
rect 15932 34018 15988 34030
rect 15932 33966 15934 34018
rect 15986 33966 15988 34018
rect 15932 33460 15988 33966
rect 16044 34020 16100 34078
rect 16044 33954 16100 33964
rect 16156 34130 16212 37774
rect 16380 37268 16436 38892
rect 16604 38724 16660 38762
rect 16604 38658 16660 38668
rect 16940 38612 16996 39228
rect 16940 38546 16996 38556
rect 17276 39284 17332 39294
rect 16716 37828 16772 37838
rect 16604 37826 16772 37828
rect 16604 37774 16718 37826
rect 16770 37774 16772 37826
rect 16604 37772 16772 37774
rect 16604 37380 16660 37772
rect 16716 37762 16772 37772
rect 17164 37826 17220 37838
rect 17164 37774 17166 37826
rect 17218 37774 17220 37826
rect 16268 37212 16436 37268
rect 16492 37268 16548 37278
rect 16268 35812 16324 37212
rect 16492 37174 16548 37212
rect 16380 37042 16436 37054
rect 16380 36990 16382 37042
rect 16434 36990 16436 37042
rect 16380 36820 16436 36990
rect 16380 36754 16436 36764
rect 16604 36596 16660 37324
rect 17164 37268 17220 37774
rect 17164 37202 17220 37212
rect 16716 37042 16772 37054
rect 16716 36990 16718 37042
rect 16770 36990 16772 37042
rect 16716 36932 16772 36990
rect 16828 37044 16884 37054
rect 16828 36950 16884 36988
rect 16716 36866 16772 36876
rect 16716 36708 16772 36746
rect 16716 36642 16772 36652
rect 16268 35680 16324 35756
rect 16380 36540 16660 36596
rect 16156 34078 16158 34130
rect 16210 34078 16212 34130
rect 16156 33572 16212 34078
rect 16044 33460 16100 33470
rect 15932 33458 16100 33460
rect 15932 33406 16046 33458
rect 16098 33406 16100 33458
rect 15932 33404 16100 33406
rect 16044 33394 16100 33404
rect 15820 33346 15876 33358
rect 15820 33294 15822 33346
rect 15874 33294 15876 33346
rect 15820 32788 15876 33294
rect 15820 32694 15876 32732
rect 16044 33236 16100 33246
rect 15484 31938 15540 31948
rect 15596 31892 15764 31948
rect 15820 32452 15876 32462
rect 15484 31666 15540 31678
rect 15484 31614 15486 31666
rect 15538 31614 15540 31666
rect 15484 31444 15540 31614
rect 15484 31378 15540 31388
rect 15596 31556 15652 31892
rect 15372 30942 15374 30994
rect 15426 30942 15428 30994
rect 15372 30930 15428 30942
rect 15596 30772 15652 31500
rect 15820 31778 15876 32396
rect 15820 31726 15822 31778
rect 15874 31726 15876 31778
rect 15372 30716 15652 30772
rect 15708 30770 15764 30782
rect 15708 30718 15710 30770
rect 15762 30718 15764 30770
rect 15260 30324 15316 30334
rect 15148 30322 15316 30324
rect 15148 30270 15262 30322
rect 15314 30270 15316 30322
rect 15148 30268 15316 30270
rect 15260 30258 15316 30268
rect 15036 29810 15092 29820
rect 15260 29652 15316 29662
rect 15372 29652 15428 30716
rect 15708 30324 15764 30718
rect 15708 30258 15764 30268
rect 15820 30100 15876 31726
rect 16044 30884 16100 33180
rect 16156 32452 16212 33516
rect 16268 33460 16324 33470
rect 16268 33346 16324 33404
rect 16268 33294 16270 33346
rect 16322 33294 16324 33346
rect 16268 33282 16324 33294
rect 16380 33348 16436 36540
rect 16716 36484 16772 36494
rect 16716 36370 16772 36428
rect 16716 36318 16718 36370
rect 16770 36318 16772 36370
rect 16716 36306 16772 36318
rect 16828 36372 16884 36382
rect 16828 36278 16884 36316
rect 17052 36372 17108 36382
rect 16940 35924 16996 35934
rect 16940 35830 16996 35868
rect 16492 35812 16548 35822
rect 16492 34914 16548 35756
rect 16604 35700 16660 35710
rect 16828 35700 16884 35710
rect 16660 35644 16772 35700
rect 16604 35606 16660 35644
rect 16716 35364 16772 35644
rect 16828 35606 16884 35644
rect 16940 35476 16996 35486
rect 16716 35308 16884 35364
rect 16492 34862 16494 34914
rect 16546 34862 16548 34914
rect 16492 34850 16548 34862
rect 16604 35140 16660 35150
rect 16380 33282 16436 33292
rect 16380 33124 16436 33134
rect 16268 33122 16436 33124
rect 16268 33070 16382 33122
rect 16434 33070 16436 33122
rect 16268 33068 16436 33070
rect 16268 32564 16324 33068
rect 16380 33058 16436 33068
rect 16492 33122 16548 33134
rect 16492 33070 16494 33122
rect 16546 33070 16548 33122
rect 16380 32676 16436 32686
rect 16492 32676 16548 33070
rect 16380 32674 16548 32676
rect 16380 32622 16382 32674
rect 16434 32622 16548 32674
rect 16380 32620 16548 32622
rect 16380 32610 16436 32620
rect 16268 32498 16324 32508
rect 16156 32386 16212 32396
rect 16492 32452 16548 32462
rect 16492 32358 16548 32396
rect 16156 31554 16212 31566
rect 16156 31502 16158 31554
rect 16210 31502 16212 31554
rect 16156 30996 16212 31502
rect 16492 31108 16548 31118
rect 16492 31014 16548 31052
rect 16156 30930 16212 30940
rect 16044 30818 16100 30828
rect 16604 30772 16660 35084
rect 16828 35138 16884 35308
rect 16828 35086 16830 35138
rect 16882 35086 16884 35138
rect 16828 35074 16884 35086
rect 16716 34690 16772 34702
rect 16716 34638 16718 34690
rect 16770 34638 16772 34690
rect 16716 33348 16772 34638
rect 16828 34244 16884 34254
rect 16828 33796 16884 34188
rect 16940 34020 16996 35420
rect 17052 34804 17108 36316
rect 17052 34738 17108 34748
rect 17164 35924 17220 35934
rect 16940 34018 17108 34020
rect 16940 33966 16942 34018
rect 16994 33966 17108 34018
rect 16940 33964 17108 33966
rect 16940 33954 16996 33964
rect 16940 33796 16996 33806
rect 16828 33740 16940 33796
rect 16716 33292 16884 33348
rect 16716 33124 16772 33134
rect 16716 32562 16772 33068
rect 16716 32510 16718 32562
rect 16770 32510 16772 32562
rect 16716 32498 16772 32510
rect 16828 32340 16884 33292
rect 16940 32562 16996 33740
rect 17052 33124 17108 33964
rect 17052 33058 17108 33068
rect 16940 32510 16942 32562
rect 16994 32510 16996 32562
rect 16940 32498 16996 32510
rect 16828 32274 16884 32284
rect 16828 32004 16884 32014
rect 16828 31890 16884 31948
rect 16828 31838 16830 31890
rect 16882 31838 16884 31890
rect 16828 31826 16884 31838
rect 17052 31780 17108 31790
rect 17052 31218 17108 31724
rect 17052 31166 17054 31218
rect 17106 31166 17108 31218
rect 17052 31154 17108 31166
rect 16492 30716 16660 30772
rect 16716 31108 16772 31118
rect 16380 30212 16436 30222
rect 16380 30118 16436 30156
rect 15260 29650 15428 29652
rect 15260 29598 15262 29650
rect 15314 29598 15428 29650
rect 15260 29596 15428 29598
rect 15260 29586 15316 29596
rect 14924 29484 15204 29540
rect 14924 29428 14980 29484
rect 14924 29362 14980 29372
rect 15148 29426 15204 29484
rect 15148 29374 15150 29426
rect 15202 29374 15204 29426
rect 14812 29138 14868 29148
rect 15148 28980 15204 29374
rect 15260 29428 15316 29438
rect 15260 29202 15316 29372
rect 15260 29150 15262 29202
rect 15314 29150 15316 29202
rect 15260 29138 15316 29150
rect 15148 28924 15316 28980
rect 14924 28756 14980 28794
rect 14924 28690 14980 28700
rect 15036 28644 15092 28654
rect 14924 28532 14980 28542
rect 14924 28438 14980 28476
rect 14588 28364 14756 28420
rect 14588 28308 14644 28364
rect 14252 26796 14420 26852
rect 14476 28252 14644 28308
rect 14028 26628 14084 26638
rect 14028 26402 14084 26572
rect 14028 26350 14030 26402
rect 14082 26350 14084 26402
rect 14028 26338 14084 26350
rect 14140 26404 14196 26414
rect 14140 26290 14196 26348
rect 14140 26238 14142 26290
rect 14194 26238 14196 26290
rect 14140 26226 14196 26238
rect 13916 26114 13972 26124
rect 14252 26068 14308 26796
rect 14476 26516 14532 28252
rect 14700 27970 14756 27982
rect 14700 27918 14702 27970
rect 14754 27918 14756 27970
rect 14476 26450 14532 26460
rect 14588 27636 14644 27646
rect 14588 27298 14644 27580
rect 14588 27246 14590 27298
rect 14642 27246 14644 27298
rect 13804 25620 13860 25630
rect 13692 25618 13860 25620
rect 13692 25566 13806 25618
rect 13858 25566 13860 25618
rect 13692 25564 13860 25566
rect 13804 25554 13860 25564
rect 14140 25620 14196 25630
rect 14252 25620 14308 26012
rect 14140 25618 14308 25620
rect 14140 25566 14142 25618
rect 14194 25566 14308 25618
rect 14140 25564 14308 25566
rect 14028 25508 14084 25518
rect 14028 24724 14084 25452
rect 14140 24948 14196 25564
rect 14588 25396 14644 27246
rect 14700 27188 14756 27918
rect 14700 27122 14756 27132
rect 14140 24882 14196 24892
rect 14252 25340 14644 25396
rect 14700 26628 14756 26638
rect 14140 24724 14196 24734
rect 13580 23314 13636 23324
rect 13916 24722 14196 24724
rect 13916 24670 14142 24722
rect 14194 24670 14196 24722
rect 13916 24668 14196 24670
rect 13916 23938 13972 24668
rect 14140 24658 14196 24668
rect 13916 23886 13918 23938
rect 13970 23886 13972 23938
rect 13916 23604 13972 23886
rect 12796 23268 12852 23278
rect 12796 23174 12852 23212
rect 13804 23268 13860 23278
rect 12908 23154 12964 23166
rect 12908 23102 12910 23154
rect 12962 23102 12964 23154
rect 12796 22930 12852 22942
rect 12796 22878 12798 22930
rect 12850 22878 12852 22930
rect 12796 22370 12852 22878
rect 12796 22318 12798 22370
rect 12850 22318 12852 22370
rect 12796 22306 12852 22318
rect 12908 22148 12964 23102
rect 12684 22082 12740 22092
rect 12796 22092 12964 22148
rect 13020 23156 13076 23166
rect 12572 21476 12628 21486
rect 12796 21476 12852 22092
rect 12572 21474 12852 21476
rect 12572 21422 12574 21474
rect 12626 21422 12852 21474
rect 12572 21420 12852 21422
rect 12908 21586 12964 21598
rect 12908 21534 12910 21586
rect 12962 21534 12964 21586
rect 12572 21364 12628 21420
rect 12572 21298 12628 21308
rect 12908 21026 12964 21534
rect 12908 20974 12910 21026
rect 12962 20974 12964 21026
rect 12908 20962 12964 20974
rect 12796 20690 12852 20702
rect 12796 20638 12798 20690
rect 12850 20638 12852 20690
rect 12460 20132 12740 20188
rect 12572 20020 12628 20030
rect 12572 19926 12628 19964
rect 12124 19346 12404 19348
rect 12124 19294 12126 19346
rect 12178 19294 12404 19346
rect 12124 19292 12404 19294
rect 12572 19348 12628 19358
rect 12124 19282 12180 19292
rect 12572 19254 12628 19292
rect 12124 19124 12180 19134
rect 12124 18564 12180 19068
rect 12124 18450 12180 18508
rect 12124 18398 12126 18450
rect 12178 18398 12180 18450
rect 12124 18386 12180 18398
rect 12572 18452 12628 18462
rect 12572 18358 12628 18396
rect 12236 17442 12292 17454
rect 12236 17390 12238 17442
rect 12290 17390 12292 17442
rect 12012 17042 12068 17052
rect 12124 17108 12180 17118
rect 12236 17108 12292 17390
rect 12124 17106 12292 17108
rect 12124 17054 12126 17106
rect 12178 17054 12292 17106
rect 12124 17052 12292 17054
rect 12124 17042 12180 17052
rect 12236 16884 12292 17052
rect 12236 16818 12292 16828
rect 11788 16270 11790 16322
rect 11842 16270 11844 16322
rect 11788 16258 11844 16270
rect 12572 16212 12628 16222
rect 12684 16212 12740 20132
rect 12796 19458 12852 20638
rect 13020 20188 13076 23100
rect 13804 22258 13860 23212
rect 13916 22372 13972 23548
rect 14028 24500 14084 24510
rect 14028 23378 14084 24444
rect 14028 23326 14030 23378
rect 14082 23326 14084 23378
rect 14028 23314 14084 23326
rect 13916 22370 14084 22372
rect 13916 22318 13918 22370
rect 13970 22318 14084 22370
rect 13916 22316 14084 22318
rect 13916 22306 13972 22316
rect 13804 22206 13806 22258
rect 13858 22206 13860 22258
rect 13132 22148 13188 22158
rect 13580 22148 13636 22158
rect 13132 21252 13188 22092
rect 13468 22146 13636 22148
rect 13468 22094 13582 22146
rect 13634 22094 13636 22146
rect 13468 22092 13636 22094
rect 13244 21588 13300 21598
rect 13468 21588 13524 22092
rect 13580 22082 13636 22092
rect 13244 21586 13524 21588
rect 13244 21534 13246 21586
rect 13298 21534 13524 21586
rect 13244 21532 13524 21534
rect 13244 21522 13300 21532
rect 13132 21186 13188 21196
rect 13468 21028 13524 21532
rect 13468 20962 13524 20972
rect 13692 21364 13748 21374
rect 13692 21026 13748 21308
rect 13692 20974 13694 21026
rect 13746 20974 13748 21026
rect 13692 20962 13748 20974
rect 13804 20804 13860 22206
rect 13692 20748 13860 20804
rect 13916 21028 13972 21038
rect 12796 19406 12798 19458
rect 12850 19406 12852 19458
rect 12796 19394 12852 19406
rect 12908 20132 13076 20188
rect 13356 20580 13412 20590
rect 12908 19236 12964 20132
rect 13244 20018 13300 20030
rect 13244 19966 13246 20018
rect 13298 19966 13300 20018
rect 13132 19460 13188 19470
rect 13244 19460 13300 19966
rect 13356 19906 13412 20524
rect 13356 19854 13358 19906
rect 13410 19854 13412 19906
rect 13356 19842 13412 19854
rect 13132 19458 13300 19460
rect 13132 19406 13134 19458
rect 13186 19406 13300 19458
rect 13132 19404 13300 19406
rect 13132 19394 13188 19404
rect 12908 19180 13076 19236
rect 12908 19012 12964 19022
rect 12908 18918 12964 18956
rect 13020 17890 13076 19180
rect 13020 17838 13022 17890
rect 13074 17838 13076 17890
rect 13020 17826 13076 17838
rect 12572 16210 12740 16212
rect 12572 16158 12574 16210
rect 12626 16158 12740 16210
rect 12572 16156 12740 16158
rect 13020 16212 13076 16222
rect 12572 16146 12628 16156
rect 13020 16118 13076 16156
rect 11788 15316 11844 15326
rect 11788 15222 11844 15260
rect 11564 15138 11620 15148
rect 13020 14756 13076 14766
rect 13244 14756 13300 19404
rect 13580 19010 13636 19022
rect 13580 18958 13582 19010
rect 13634 18958 13636 19010
rect 13580 18788 13636 18958
rect 13356 18732 13636 18788
rect 13356 18452 13412 18732
rect 13356 18386 13412 18396
rect 13468 18564 13524 18574
rect 13468 17668 13524 18508
rect 13580 18450 13636 18462
rect 13580 18398 13582 18450
rect 13634 18398 13636 18450
rect 13580 17890 13636 18398
rect 13580 17838 13582 17890
rect 13634 17838 13636 17890
rect 13580 17826 13636 17838
rect 13580 17668 13636 17678
rect 13468 17666 13636 17668
rect 13468 17614 13582 17666
rect 13634 17614 13636 17666
rect 13468 17612 13636 17614
rect 13580 17602 13636 17612
rect 13580 16322 13636 16334
rect 13580 16270 13582 16322
rect 13634 16270 13636 16322
rect 13020 14754 13300 14756
rect 13020 14702 13022 14754
rect 13074 14702 13300 14754
rect 13020 14700 13300 14702
rect 13468 15876 13524 15886
rect 13020 14690 13076 14700
rect 12460 14306 12516 14318
rect 12460 14254 12462 14306
rect 12514 14254 12516 14306
rect 11228 13748 11284 13758
rect 11228 13654 11284 13692
rect 11116 13346 11172 13356
rect 11900 13412 11956 13422
rect 10892 13022 10894 13074
rect 10946 13022 10948 13074
rect 10892 13010 10948 13022
rect 11340 13188 11396 13198
rect 11340 13074 11396 13132
rect 11340 13022 11342 13074
rect 11394 13022 11396 13074
rect 10668 12350 10670 12402
rect 10722 12350 10724 12402
rect 9100 12126 9102 12178
rect 9154 12126 9156 12178
rect 9100 10834 9156 12126
rect 10668 11620 10724 12350
rect 11116 12964 11172 12974
rect 10892 11620 10948 11630
rect 10668 11618 10948 11620
rect 10668 11566 10894 11618
rect 10946 11566 10948 11618
rect 10668 11564 10948 11566
rect 10556 11508 10612 11518
rect 10668 11508 10724 11564
rect 10892 11554 10948 11564
rect 10556 11506 10724 11508
rect 10556 11454 10558 11506
rect 10610 11454 10724 11506
rect 10556 11452 10724 11454
rect 11116 11506 11172 12908
rect 11340 12964 11396 13022
rect 11340 12898 11396 12908
rect 11900 12964 11956 13356
rect 12348 13076 12404 13086
rect 12460 13076 12516 14254
rect 12348 13074 12516 13076
rect 12348 13022 12350 13074
rect 12402 13022 12516 13074
rect 12348 13020 12516 13022
rect 12348 13010 12404 13020
rect 11900 12870 11956 12908
rect 12460 12964 12516 13020
rect 12460 12898 12516 12908
rect 12908 12964 12964 12974
rect 12908 12870 12964 12908
rect 13468 12852 13524 15820
rect 13580 15876 13636 16270
rect 13692 16212 13748 20748
rect 13916 20690 13972 20972
rect 13916 20638 13918 20690
rect 13970 20638 13972 20690
rect 13916 20626 13972 20638
rect 13804 20580 13860 20590
rect 13804 20486 13860 20524
rect 14028 20188 14084 22316
rect 13916 20132 14084 20188
rect 14140 20916 14196 20926
rect 13916 19012 13972 20132
rect 13916 18946 13972 18956
rect 14028 19908 14084 19918
rect 14028 18450 14084 19852
rect 14028 18398 14030 18450
rect 14082 18398 14084 18450
rect 14028 18386 14084 18398
rect 14140 17778 14196 20860
rect 14252 20188 14308 25340
rect 14700 25284 14756 26572
rect 14364 25228 14756 25284
rect 14364 21812 14420 25228
rect 14924 24948 14980 24958
rect 14700 24724 14756 24734
rect 14588 24722 14756 24724
rect 14588 24670 14702 24722
rect 14754 24670 14756 24722
rect 14588 24668 14756 24670
rect 14588 23938 14644 24668
rect 14700 24658 14756 24668
rect 14588 23886 14590 23938
rect 14642 23886 14644 23938
rect 14476 23380 14532 23390
rect 14476 23286 14532 23324
rect 14476 21812 14532 21822
rect 14364 21810 14532 21812
rect 14364 21758 14478 21810
rect 14530 21758 14532 21810
rect 14364 21756 14532 21758
rect 14476 21746 14532 21756
rect 14588 21252 14644 23886
rect 14924 23378 14980 24892
rect 14924 23326 14926 23378
rect 14978 23326 14980 23378
rect 14924 23314 14980 23326
rect 14812 22484 14868 22494
rect 15036 22484 15092 28588
rect 15148 27972 15204 27982
rect 15148 27858 15204 27916
rect 15148 27806 15150 27858
rect 15202 27806 15204 27858
rect 15148 27794 15204 27806
rect 15260 26908 15316 28924
rect 15372 28642 15428 29596
rect 15372 28590 15374 28642
rect 15426 28590 15428 28642
rect 15372 27748 15428 28590
rect 15372 27682 15428 27692
rect 15484 30044 15876 30100
rect 15372 27076 15428 27086
rect 15372 26982 15428 27020
rect 15148 26852 15316 26908
rect 15148 24050 15204 26852
rect 15372 26290 15428 26302
rect 15372 26238 15374 26290
rect 15426 26238 15428 26290
rect 15148 23998 15150 24050
rect 15202 23998 15204 24050
rect 15148 23492 15204 23998
rect 15148 23426 15204 23436
rect 15260 26178 15316 26190
rect 15260 26126 15262 26178
rect 15314 26126 15316 26178
rect 15260 25618 15316 26126
rect 15260 25566 15262 25618
rect 15314 25566 15316 25618
rect 14812 22482 15092 22484
rect 14812 22430 14814 22482
rect 14866 22430 15092 22482
rect 14812 22428 15092 22430
rect 14812 22418 14868 22428
rect 15148 22148 15204 22158
rect 15148 22054 15204 22092
rect 14924 21476 14980 21486
rect 14924 21474 15204 21476
rect 14924 21422 14926 21474
rect 14978 21422 15204 21474
rect 14924 21420 15204 21422
rect 14924 21410 14980 21420
rect 14588 21196 15092 21252
rect 14812 20578 14868 20590
rect 14812 20526 14814 20578
rect 14866 20526 14868 20578
rect 14252 20132 14532 20188
rect 14476 20130 14532 20132
rect 14476 20078 14478 20130
rect 14530 20078 14532 20130
rect 14476 20066 14532 20078
rect 14364 19348 14420 19358
rect 14364 19254 14420 19292
rect 14140 17726 14142 17778
rect 14194 17726 14196 17778
rect 13692 16146 13748 16156
rect 13916 16884 13972 16894
rect 13580 15874 13748 15876
rect 13580 15822 13582 15874
rect 13634 15822 13748 15874
rect 13580 15820 13748 15822
rect 13580 15810 13636 15820
rect 13692 14642 13748 15820
rect 13916 14644 13972 16828
rect 14028 16772 14084 16782
rect 14028 15876 14084 16716
rect 14028 15782 14084 15820
rect 14140 14756 14196 17726
rect 14700 19012 14756 19022
rect 14588 17444 14644 17454
rect 14700 17444 14756 18956
rect 14364 17442 14756 17444
rect 14364 17390 14590 17442
rect 14642 17390 14756 17442
rect 14364 17388 14756 17390
rect 14364 16322 14420 17388
rect 14588 17378 14644 17388
rect 14476 16884 14532 16894
rect 14812 16884 14868 20526
rect 15036 17442 15092 21196
rect 15148 20802 15204 21420
rect 15260 20916 15316 25566
rect 15372 25508 15428 26238
rect 15372 25414 15428 25452
rect 15484 23380 15540 30044
rect 15820 29540 15876 29550
rect 16492 29540 16548 30716
rect 16604 30324 16660 30334
rect 16604 30230 16660 30268
rect 15708 28084 15764 28094
rect 15708 27990 15764 28028
rect 15596 27858 15652 27870
rect 15820 27860 15876 29484
rect 16380 29484 16548 29540
rect 16604 29652 16660 29662
rect 16156 29428 16212 29438
rect 16156 29334 16212 29372
rect 16156 28308 16212 28318
rect 15596 27806 15598 27858
rect 15650 27806 15652 27858
rect 15596 27636 15652 27806
rect 15596 27570 15652 27580
rect 15708 27804 15876 27860
rect 15932 28084 15988 28094
rect 15708 26852 15764 27804
rect 15820 26964 15876 27002
rect 15820 26898 15876 26908
rect 15708 26786 15764 26796
rect 15708 24948 15764 24958
rect 15708 24854 15764 24892
rect 15484 23314 15540 23324
rect 15596 23492 15652 23502
rect 15484 23156 15540 23166
rect 15484 23062 15540 23100
rect 15596 22482 15652 23436
rect 15596 22430 15598 22482
rect 15650 22430 15652 22482
rect 15596 22418 15652 22430
rect 15820 21812 15876 21822
rect 15596 21588 15652 21598
rect 15596 21494 15652 21532
rect 15820 21586 15876 21756
rect 15820 21534 15822 21586
rect 15874 21534 15876 21586
rect 15820 21476 15876 21534
rect 15820 21410 15876 21420
rect 15260 20850 15316 20860
rect 15820 20916 15876 20926
rect 15932 20916 15988 28028
rect 16156 27972 16212 28252
rect 16380 28084 16436 29484
rect 16380 28018 16436 28028
rect 16492 29316 16548 29326
rect 16604 29316 16660 29596
rect 16492 29314 16660 29316
rect 16492 29262 16494 29314
rect 16546 29262 16660 29314
rect 16492 29260 16660 29262
rect 16156 27906 16212 27916
rect 16492 27972 16548 29260
rect 16604 28420 16660 28430
rect 16604 28082 16660 28364
rect 16604 28030 16606 28082
rect 16658 28030 16660 28082
rect 16604 28018 16660 28030
rect 16268 27748 16324 27758
rect 16268 25394 16324 27692
rect 16380 26962 16436 26974
rect 16380 26910 16382 26962
rect 16434 26910 16436 26962
rect 16380 26068 16436 26910
rect 16492 26908 16548 27916
rect 16716 27860 16772 31052
rect 16828 30996 16884 31006
rect 16828 30434 16884 30940
rect 16828 30382 16830 30434
rect 16882 30382 16884 30434
rect 16828 30370 16884 30382
rect 16940 30436 16996 30446
rect 16940 29540 16996 30380
rect 17164 30324 17220 35868
rect 17276 35028 17332 39228
rect 17388 38836 17444 39454
rect 17388 38770 17444 38780
rect 17500 39394 17556 39406
rect 17500 39342 17502 39394
rect 17554 39342 17556 39394
rect 17388 37044 17444 37054
rect 17388 36706 17444 36988
rect 17388 36654 17390 36706
rect 17442 36654 17444 36706
rect 17388 36642 17444 36654
rect 17500 35252 17556 39342
rect 17724 39284 17780 39294
rect 17836 39284 17892 39564
rect 17948 39508 18004 40124
rect 18844 40068 18900 40348
rect 18844 40002 18900 40012
rect 17948 39442 18004 39452
rect 18060 39844 18116 39854
rect 17836 39228 18004 39284
rect 17724 38946 17780 39228
rect 17724 38894 17726 38946
rect 17778 38894 17780 38946
rect 17724 38882 17780 38894
rect 17948 38946 18004 39228
rect 17948 38894 17950 38946
rect 18002 38894 18004 38946
rect 17948 38882 18004 38894
rect 17836 38836 17892 38846
rect 17836 38668 17892 38780
rect 17612 38612 17668 38622
rect 17836 38612 18004 38668
rect 17612 38162 17668 38556
rect 17612 38110 17614 38162
rect 17666 38110 17668 38162
rect 17612 38098 17668 38110
rect 17836 37716 17892 37726
rect 17836 37490 17892 37660
rect 17836 37438 17838 37490
rect 17890 37438 17892 37490
rect 17724 37156 17780 37166
rect 17612 36482 17668 36494
rect 17612 36430 17614 36482
rect 17666 36430 17668 36482
rect 17612 35700 17668 36430
rect 17724 35810 17780 37100
rect 17836 36820 17892 37438
rect 17948 37490 18004 38612
rect 17948 37438 17950 37490
rect 18002 37438 18004 37490
rect 17948 37426 18004 37438
rect 18060 37378 18116 39788
rect 18620 39732 18676 39770
rect 18620 39666 18676 39676
rect 18284 39620 18340 39630
rect 18284 39284 18340 39564
rect 18732 39620 18788 39630
rect 18620 39508 18676 39518
rect 18284 39218 18340 39228
rect 18396 39396 18452 39406
rect 18284 38948 18340 38958
rect 18284 38854 18340 38892
rect 18172 38724 18228 38762
rect 18172 38658 18228 38668
rect 18172 38164 18228 38174
rect 18172 38070 18228 38108
rect 18060 37326 18062 37378
rect 18114 37326 18116 37378
rect 18060 36932 18116 37326
rect 18172 37604 18228 37614
rect 18172 37378 18228 37548
rect 18172 37326 18174 37378
rect 18226 37326 18228 37378
rect 18172 37314 18228 37326
rect 18396 37378 18452 39340
rect 18508 39394 18564 39406
rect 18508 39342 18510 39394
rect 18562 39342 18564 39394
rect 18508 39060 18564 39342
rect 18620 39172 18676 39452
rect 18732 39506 18788 39564
rect 18732 39454 18734 39506
rect 18786 39454 18788 39506
rect 18732 39442 18788 39454
rect 18844 39396 18900 39406
rect 18844 39302 18900 39340
rect 19068 39396 19124 39406
rect 18620 39116 18788 39172
rect 18508 38994 18564 39004
rect 18508 38274 18564 38286
rect 18508 38222 18510 38274
rect 18562 38222 18564 38274
rect 18508 38162 18564 38222
rect 18508 38110 18510 38162
rect 18562 38110 18564 38162
rect 18508 38098 18564 38110
rect 18396 37326 18398 37378
rect 18450 37326 18452 37378
rect 18396 37314 18452 37326
rect 18060 36866 18116 36876
rect 18508 37268 18564 37278
rect 17836 36764 18004 36820
rect 17836 36596 17892 36606
rect 17836 36502 17892 36540
rect 17724 35758 17726 35810
rect 17778 35758 17780 35810
rect 17724 35746 17780 35758
rect 17836 36036 17892 36046
rect 17612 35634 17668 35644
rect 17500 35186 17556 35196
rect 17500 35028 17556 35038
rect 17276 35026 17556 35028
rect 17276 34974 17502 35026
rect 17554 34974 17556 35026
rect 17276 34972 17556 34974
rect 17500 34916 17556 34972
rect 17500 34850 17556 34860
rect 17276 34692 17332 34702
rect 17276 31780 17332 34636
rect 17836 34468 17892 35980
rect 17948 35924 18004 36764
rect 18284 36596 18340 36606
rect 18172 36484 18228 36494
rect 18172 36390 18228 36428
rect 18284 36482 18340 36540
rect 18284 36430 18286 36482
rect 18338 36430 18340 36482
rect 18060 36258 18116 36270
rect 18060 36206 18062 36258
rect 18114 36206 18116 36258
rect 18060 36148 18116 36206
rect 18060 36082 18116 36092
rect 18284 35924 18340 36430
rect 17948 35868 18116 35924
rect 17948 35698 18004 35710
rect 17948 35646 17950 35698
rect 18002 35646 18004 35698
rect 17948 35028 18004 35646
rect 17948 34962 18004 34972
rect 17948 34692 18004 34702
rect 17948 34598 18004 34636
rect 17724 34412 18004 34468
rect 17612 34130 17668 34142
rect 17612 34078 17614 34130
rect 17666 34078 17668 34130
rect 17276 31714 17332 31724
rect 17388 34020 17444 34030
rect 17388 33234 17444 33964
rect 17612 33572 17668 34078
rect 17612 33506 17668 33516
rect 17724 33348 17780 34412
rect 17836 34242 17892 34254
rect 17836 34190 17838 34242
rect 17890 34190 17892 34242
rect 17836 34020 17892 34190
rect 17948 34242 18004 34412
rect 17948 34190 17950 34242
rect 18002 34190 18004 34242
rect 17948 34178 18004 34190
rect 17836 33954 17892 33964
rect 17388 33182 17390 33234
rect 17442 33182 17444 33234
rect 17388 32788 17444 33182
rect 17612 33292 17780 33348
rect 17836 33348 17892 33358
rect 17612 33234 17668 33292
rect 17836 33254 17892 33292
rect 17948 33348 18004 33358
rect 18060 33348 18116 35868
rect 18284 35858 18340 35868
rect 18284 35700 18340 35710
rect 18508 35700 18564 37212
rect 18620 36820 18676 36830
rect 18620 35922 18676 36764
rect 18620 35870 18622 35922
rect 18674 35870 18676 35922
rect 18620 35858 18676 35870
rect 18508 35644 18676 35700
rect 18284 35606 18340 35644
rect 18508 35474 18564 35486
rect 18508 35422 18510 35474
rect 18562 35422 18564 35474
rect 18508 35140 18564 35422
rect 18508 35074 18564 35084
rect 18396 35028 18452 35038
rect 18396 33796 18452 34972
rect 18620 34468 18676 35644
rect 18620 34402 18676 34412
rect 18732 34244 18788 39116
rect 18956 39060 19012 39070
rect 18956 38668 19012 39004
rect 18844 38612 19012 38668
rect 18844 37268 18900 38612
rect 19068 38052 19124 39340
rect 19180 38948 19236 38958
rect 19180 38834 19236 38892
rect 19180 38782 19182 38834
rect 19234 38782 19236 38834
rect 19180 38770 19236 38782
rect 19292 38612 19348 40572
rect 19628 40534 19684 40572
rect 20188 40516 20244 41246
rect 20748 41300 20804 41310
rect 19964 40460 20244 40516
rect 20412 41076 20468 41086
rect 19516 40178 19572 40190
rect 19516 40126 19518 40178
rect 19570 40126 19572 40178
rect 19404 39732 19460 39742
rect 19404 39618 19460 39676
rect 19404 39566 19406 39618
rect 19458 39566 19460 39618
rect 19404 39554 19460 39566
rect 19516 38946 19572 40126
rect 19964 40178 20020 40460
rect 20076 40292 20132 40302
rect 20076 40290 20244 40292
rect 20076 40238 20078 40290
rect 20130 40238 20244 40290
rect 20076 40236 20244 40238
rect 20076 40226 20132 40236
rect 19964 40126 19966 40178
rect 20018 40126 20020 40178
rect 19964 40114 20020 40126
rect 20188 40180 20244 40236
rect 19964 39732 20020 39742
rect 19964 39638 20020 39676
rect 19852 39508 19908 39518
rect 19852 39414 19908 39452
rect 20076 39396 20132 39434
rect 20076 39330 20132 39340
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19516 38894 19518 38946
rect 19570 38894 19572 38946
rect 19516 38882 19572 38894
rect 20188 38948 20244 40124
rect 20188 38882 20244 38892
rect 19404 38836 19460 38846
rect 19404 38742 19460 38780
rect 19292 38546 19348 38556
rect 19628 38612 19684 38622
rect 19404 38500 19460 38510
rect 18844 37202 18900 37212
rect 18956 37996 19124 38052
rect 19292 38274 19348 38286
rect 19292 38222 19294 38274
rect 19346 38222 19348 38274
rect 18956 36820 19012 37996
rect 19068 37828 19124 37838
rect 19292 37828 19348 38222
rect 19404 38050 19460 38444
rect 19404 37998 19406 38050
rect 19458 37998 19460 38050
rect 19404 37986 19460 37998
rect 19292 37772 19460 37828
rect 19068 37734 19124 37772
rect 19292 37268 19348 37278
rect 18956 36754 19012 36764
rect 19180 36932 19236 36942
rect 18956 36482 19012 36494
rect 18956 36430 18958 36482
rect 19010 36430 19012 36482
rect 18956 36036 19012 36430
rect 19180 36482 19236 36876
rect 19292 36708 19348 37212
rect 19404 37154 19460 37772
rect 19404 37102 19406 37154
rect 19458 37102 19460 37154
rect 19404 37042 19460 37102
rect 19404 36990 19406 37042
rect 19458 36990 19460 37042
rect 19404 36978 19460 36990
rect 19516 37044 19572 37054
rect 19404 36708 19460 36718
rect 19292 36706 19460 36708
rect 19292 36654 19406 36706
rect 19458 36654 19460 36706
rect 19292 36652 19460 36654
rect 19404 36642 19460 36652
rect 19180 36430 19182 36482
rect 19234 36430 19236 36482
rect 18956 35970 19012 35980
rect 19068 36258 19124 36270
rect 19068 36206 19070 36258
rect 19122 36206 19124 36258
rect 19068 35700 19124 36206
rect 19068 35634 19124 35644
rect 19180 35476 19236 36430
rect 19404 35924 19460 35934
rect 19404 35830 19460 35868
rect 19180 35410 19236 35420
rect 18396 33730 18452 33740
rect 18620 34188 18788 34244
rect 18844 35252 18900 35262
rect 18620 33460 18676 34188
rect 18732 34020 18788 34030
rect 18732 33926 18788 33964
rect 18620 33404 18788 33460
rect 17948 33346 18116 33348
rect 17948 33294 17950 33346
rect 18002 33294 18116 33346
rect 17948 33292 18116 33294
rect 17948 33282 18004 33292
rect 17612 33182 17614 33234
rect 17666 33182 17668 33234
rect 17612 33170 17668 33182
rect 17724 33124 17780 33134
rect 17724 33030 17780 33068
rect 17276 31556 17332 31566
rect 17388 31556 17444 32732
rect 17948 32452 18004 32462
rect 17948 32358 18004 32396
rect 17724 32340 17780 32350
rect 17724 32246 17780 32284
rect 18060 32340 18116 33292
rect 18396 33348 18452 33358
rect 18396 33254 18452 33292
rect 18620 33236 18676 33246
rect 18620 33142 18676 33180
rect 18284 33124 18340 33134
rect 17724 31892 17780 31902
rect 17724 31798 17780 31836
rect 17276 31554 17388 31556
rect 17276 31502 17278 31554
rect 17330 31502 17388 31554
rect 17276 31500 17388 31502
rect 17276 31332 17332 31500
rect 17388 31424 17444 31500
rect 18060 31444 18116 32284
rect 18172 32450 18228 32462
rect 18172 32398 18174 32450
rect 18226 32398 18228 32450
rect 18172 31668 18228 32398
rect 18284 31890 18340 33068
rect 18396 32788 18452 32798
rect 18396 32694 18452 32732
rect 18620 32562 18676 32574
rect 18620 32510 18622 32562
rect 18674 32510 18676 32562
rect 18508 32450 18564 32462
rect 18508 32398 18510 32450
rect 18562 32398 18564 32450
rect 18508 32002 18564 32398
rect 18620 32340 18676 32510
rect 18620 32274 18676 32284
rect 18732 32228 18788 33404
rect 18844 33346 18900 35196
rect 19292 35140 19348 35150
rect 18956 34916 19012 34926
rect 18956 34822 19012 34860
rect 19180 34804 19236 34814
rect 19180 34710 19236 34748
rect 19068 34690 19124 34702
rect 19068 34638 19070 34690
rect 19122 34638 19124 34690
rect 19068 33572 19124 34638
rect 19180 34356 19236 34366
rect 19292 34356 19348 35084
rect 19404 34692 19460 34702
rect 19404 34598 19460 34636
rect 19516 34468 19572 36988
rect 19180 34354 19348 34356
rect 19180 34302 19182 34354
rect 19234 34302 19348 34354
rect 19180 34300 19348 34302
rect 19404 34412 19572 34468
rect 19628 34916 19684 38556
rect 19964 38610 20020 38622
rect 19964 38558 19966 38610
rect 20018 38558 20020 38610
rect 19964 38052 20020 38558
rect 19964 37986 20020 37996
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19964 37492 20020 37502
rect 19964 37398 20020 37436
rect 19964 37042 20020 37054
rect 19964 36990 19966 37042
rect 20018 36990 20020 37042
rect 19964 36372 20020 36990
rect 20412 36820 20468 41020
rect 20636 40964 20692 40974
rect 20524 40516 20580 40526
rect 20524 38834 20580 40460
rect 20524 38782 20526 38834
rect 20578 38782 20580 38834
rect 20524 38770 20580 38782
rect 20636 38946 20692 40908
rect 20748 40740 20804 41244
rect 20860 41300 20916 41310
rect 20972 41300 21028 41916
rect 21084 41878 21140 41916
rect 21420 41748 21476 43260
rect 21532 41860 21588 44942
rect 21644 44322 21700 45164
rect 21756 45106 21812 48190
rect 21980 47572 22036 47582
rect 21756 45054 21758 45106
rect 21810 45054 21812 45106
rect 21756 44548 21812 45054
rect 21756 44482 21812 44492
rect 21868 47236 21924 47246
rect 21644 44270 21646 44322
rect 21698 44270 21700 44322
rect 21644 44258 21700 44270
rect 21868 44322 21924 47180
rect 21980 45668 22036 47516
rect 22092 46676 22148 49868
rect 22092 46610 22148 46620
rect 22204 49812 22260 49822
rect 22092 45668 22148 45678
rect 21980 45666 22148 45668
rect 21980 45614 22094 45666
rect 22146 45614 22148 45666
rect 21980 45612 22148 45614
rect 22092 44660 22148 45612
rect 22092 44594 22148 44604
rect 22204 44548 22260 49756
rect 22316 47572 22372 50652
rect 22316 47506 22372 47516
rect 22428 47234 22484 51100
rect 22540 50036 22596 50046
rect 22540 49698 22596 49980
rect 22540 49646 22542 49698
rect 22594 49646 22596 49698
rect 22540 48916 22596 49646
rect 22540 48850 22596 48860
rect 22652 49138 22708 51884
rect 22876 51492 22932 53116
rect 22988 53060 23044 53070
rect 22988 52162 23044 53004
rect 23324 52946 23380 52958
rect 23324 52894 23326 52946
rect 23378 52894 23380 52946
rect 23324 52836 23380 52894
rect 22988 52110 22990 52162
rect 23042 52110 23044 52162
rect 22988 52098 23044 52110
rect 23100 52612 23156 52622
rect 23100 52164 23156 52556
rect 23212 52164 23268 52174
rect 23100 52162 23268 52164
rect 23100 52110 23214 52162
rect 23266 52110 23268 52162
rect 23100 52108 23268 52110
rect 23212 52098 23268 52108
rect 23324 52164 23380 52780
rect 23436 52724 23492 53564
rect 23436 52658 23492 52668
rect 23548 53730 23716 53732
rect 23548 53678 23662 53730
rect 23714 53678 23716 53730
rect 23548 53676 23716 53678
rect 23548 52946 23604 53676
rect 23660 53666 23716 53676
rect 23996 53732 24052 53742
rect 24108 53732 24164 55244
rect 24220 55076 24276 55086
rect 24220 54982 24276 55020
rect 24444 54740 24500 54750
rect 24444 54646 24500 54684
rect 23996 53730 24164 53732
rect 23996 53678 23998 53730
rect 24050 53678 24164 53730
rect 23996 53676 24164 53678
rect 24220 53732 24276 53742
rect 23996 53666 24052 53676
rect 24220 53638 24276 53676
rect 23772 53508 23828 53518
rect 23772 53058 23828 53452
rect 23884 53506 23940 53518
rect 23884 53454 23886 53506
rect 23938 53454 23940 53506
rect 23884 53172 23940 53454
rect 24108 53508 24164 53518
rect 24108 53506 24500 53508
rect 24108 53454 24110 53506
rect 24162 53454 24500 53506
rect 24108 53452 24500 53454
rect 24108 53442 24164 53452
rect 23884 53116 24388 53172
rect 23772 53006 23774 53058
rect 23826 53006 23828 53058
rect 23548 52894 23550 52946
rect 23602 52894 23604 52946
rect 23324 52098 23380 52108
rect 23100 51940 23156 51950
rect 23100 51846 23156 51884
rect 23212 51828 23268 51838
rect 22988 51492 23044 51502
rect 22876 51490 23044 51492
rect 22876 51438 22990 51490
rect 23042 51438 23044 51490
rect 22876 51436 23044 51438
rect 22876 50708 22932 51436
rect 22988 51426 23044 51436
rect 23212 51378 23268 51772
rect 23548 51602 23604 52894
rect 23660 52948 23716 52958
rect 23660 51940 23716 52892
rect 23772 52388 23828 53006
rect 23996 52946 24052 52958
rect 23996 52894 23998 52946
rect 24050 52894 24052 52946
rect 23884 52836 23940 52846
rect 23884 52742 23940 52780
rect 23996 52724 24052 52894
rect 23996 52658 24052 52668
rect 24220 52948 24276 52958
rect 23772 52332 23940 52388
rect 23772 52164 23828 52174
rect 23772 52070 23828 52108
rect 23660 51884 23828 51940
rect 23548 51550 23550 51602
rect 23602 51550 23604 51602
rect 23548 51538 23604 51550
rect 23212 51326 23214 51378
rect 23266 51326 23268 51378
rect 23212 51314 23268 51326
rect 22876 50642 22932 50652
rect 23212 50932 23268 50942
rect 22876 50484 22932 50494
rect 22764 50370 22820 50382
rect 22764 50318 22766 50370
rect 22818 50318 22820 50370
rect 22764 50036 22820 50318
rect 22764 49970 22820 49980
rect 22876 49250 22932 50428
rect 22876 49198 22878 49250
rect 22930 49198 22932 49250
rect 22876 49186 22932 49198
rect 23100 50260 23156 50270
rect 22652 49086 22654 49138
rect 22706 49086 22708 49138
rect 22652 48466 22708 49086
rect 23100 49140 23156 50204
rect 23100 49026 23156 49084
rect 23100 48974 23102 49026
rect 23154 48974 23156 49026
rect 23100 48692 23156 48974
rect 22652 48414 22654 48466
rect 22706 48414 22708 48466
rect 22652 48356 22708 48414
rect 22652 48290 22708 48300
rect 22876 48636 23100 48692
rect 22428 47182 22430 47234
rect 22482 47182 22484 47234
rect 22428 45892 22484 47182
rect 22764 47796 22820 47806
rect 22540 46562 22596 46574
rect 22540 46510 22542 46562
rect 22594 46510 22596 46562
rect 22540 46452 22596 46510
rect 22540 46386 22596 46396
rect 22652 45892 22708 45902
rect 22428 45890 22708 45892
rect 22428 45838 22654 45890
rect 22706 45838 22708 45890
rect 22428 45836 22708 45838
rect 22540 45556 22596 45566
rect 22540 44660 22596 45500
rect 22652 45108 22708 45836
rect 22764 45220 22820 47740
rect 22876 47570 22932 48636
rect 23100 48626 23156 48636
rect 23212 49588 23268 50876
rect 23660 50818 23716 50830
rect 23660 50766 23662 50818
rect 23714 50766 23716 50818
rect 23660 50706 23716 50766
rect 23660 50654 23662 50706
rect 23714 50654 23716 50706
rect 23324 50594 23380 50606
rect 23324 50542 23326 50594
rect 23378 50542 23380 50594
rect 23324 50372 23380 50542
rect 23324 50306 23380 50316
rect 23548 49812 23604 49822
rect 23436 49810 23604 49812
rect 23436 49758 23550 49810
rect 23602 49758 23604 49810
rect 23436 49756 23604 49758
rect 23436 49588 23492 49756
rect 23548 49746 23604 49756
rect 23212 49532 23492 49588
rect 22876 47518 22878 47570
rect 22930 47518 22932 47570
rect 22876 46002 22932 47518
rect 22988 48356 23044 48366
rect 22988 46898 23044 48300
rect 22988 46846 22990 46898
rect 23042 46846 23044 46898
rect 22988 46834 23044 46846
rect 23212 46676 23268 49532
rect 23660 49476 23716 50654
rect 23772 50596 23828 51884
rect 23772 49698 23828 50540
rect 23772 49646 23774 49698
rect 23826 49646 23828 49698
rect 23772 49634 23828 49646
rect 23884 49476 23940 52332
rect 24220 52162 24276 52892
rect 24332 52274 24388 53116
rect 24332 52222 24334 52274
rect 24386 52222 24388 52274
rect 24332 52210 24388 52222
rect 24220 52110 24222 52162
rect 24274 52110 24276 52162
rect 24220 52098 24276 52110
rect 24444 52164 24500 53452
rect 24556 52834 24612 56028
rect 24668 55972 24724 55982
rect 24780 55972 24836 57484
rect 24668 55970 24836 55972
rect 24668 55918 24670 55970
rect 24722 55918 24836 55970
rect 24668 55916 24836 55918
rect 24668 55906 24724 55916
rect 24668 55300 24724 55310
rect 24668 55206 24724 55244
rect 24780 54852 24836 55916
rect 25004 56980 25060 56990
rect 25004 56866 25060 56924
rect 25004 56814 25006 56866
rect 25058 56814 25060 56866
rect 25004 55860 25060 56814
rect 25116 56868 25172 56878
rect 25116 56774 25172 56812
rect 25228 56644 25284 56654
rect 25228 56550 25284 56588
rect 25060 55804 25172 55860
rect 25004 55794 25060 55804
rect 24668 54796 24836 54852
rect 24668 53508 24724 54796
rect 25004 54404 25060 54414
rect 25004 54310 25060 54348
rect 24892 53508 24948 53518
rect 24668 53442 24724 53452
rect 24780 53506 24948 53508
rect 24780 53454 24894 53506
rect 24946 53454 24948 53506
rect 24780 53452 24948 53454
rect 24668 53060 24724 53070
rect 24668 52966 24724 53004
rect 24556 52782 24558 52834
rect 24610 52782 24612 52834
rect 24556 52770 24612 52782
rect 24668 52164 24724 52174
rect 24444 52162 24724 52164
rect 24444 52110 24670 52162
rect 24722 52110 24724 52162
rect 24444 52108 24724 52110
rect 24668 52098 24724 52108
rect 24332 52052 24388 52062
rect 23660 49420 23940 49476
rect 23772 49026 23828 49038
rect 23772 48974 23774 49026
rect 23826 48974 23828 49026
rect 23660 48804 23716 48814
rect 23436 48468 23492 48478
rect 23436 48374 23492 48412
rect 23324 48356 23380 48366
rect 23324 48262 23380 48300
rect 23548 48244 23604 48254
rect 23660 48244 23716 48748
rect 23548 48242 23716 48244
rect 23548 48190 23550 48242
rect 23602 48190 23716 48242
rect 23548 48188 23716 48190
rect 23548 48178 23604 48188
rect 23548 48020 23604 48030
rect 23324 47460 23380 47470
rect 23324 47366 23380 47404
rect 23548 46900 23604 47964
rect 23436 46844 23604 46900
rect 23660 47236 23716 48188
rect 23772 48130 23828 48974
rect 23772 48078 23774 48130
rect 23826 48078 23828 48130
rect 23772 47460 23828 48078
rect 23884 47460 23940 49420
rect 24108 51828 24164 51838
rect 24108 50372 24164 51772
rect 24108 48804 24164 50316
rect 24332 51378 24388 51996
rect 24444 51940 24500 51950
rect 24444 51846 24500 51884
rect 24780 51828 24836 53452
rect 24892 53442 24948 53452
rect 24892 53172 24948 53182
rect 24892 53058 24948 53116
rect 24892 53006 24894 53058
rect 24946 53006 24948 53058
rect 24892 52994 24948 53006
rect 25004 52836 25060 52846
rect 25004 52386 25060 52780
rect 25004 52334 25006 52386
rect 25058 52334 25060 52386
rect 25004 52322 25060 52334
rect 24780 51762 24836 51772
rect 24892 52162 24948 52174
rect 25116 52164 25172 55804
rect 25340 54740 25396 60844
rect 30156 60116 30212 63181
rect 35196 60396 35460 60406
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35196 60330 35460 60340
rect 30156 60050 30212 60060
rect 31052 60116 31108 60126
rect 31052 60022 31108 60060
rect 50204 60116 50260 63181
rect 50204 60050 50260 60060
rect 51100 60116 51156 60126
rect 51100 60022 51156 60060
rect 30380 60002 30436 60014
rect 30380 59950 30382 60002
rect 30434 59950 30436 60002
rect 26908 59890 26964 59902
rect 26908 59838 26910 59890
rect 26962 59838 26964 59890
rect 25676 59668 25732 59678
rect 25676 59442 25732 59612
rect 25676 59390 25678 59442
rect 25730 59390 25732 59442
rect 25676 59378 25732 59390
rect 26684 59332 26740 59342
rect 26684 59218 26740 59276
rect 26908 59332 26964 59838
rect 27020 59780 27076 59790
rect 29820 59780 29876 59790
rect 27020 59778 27972 59780
rect 27020 59726 27022 59778
rect 27074 59726 27972 59778
rect 27020 59724 27972 59726
rect 27020 59714 27076 59724
rect 27916 59442 27972 59724
rect 29820 59686 29876 59724
rect 30380 59780 30436 59950
rect 33964 60004 34020 60014
rect 33964 60002 34244 60004
rect 33964 59950 33966 60002
rect 34018 59950 34244 60002
rect 33964 59948 34244 59950
rect 33964 59938 34020 59948
rect 33628 59890 33684 59902
rect 33628 59838 33630 59890
rect 33682 59838 33684 59890
rect 30380 59714 30436 59724
rect 33180 59780 33236 59790
rect 33628 59780 33684 59838
rect 33180 59778 33684 59780
rect 33180 59726 33182 59778
rect 33234 59726 33684 59778
rect 33180 59724 33684 59726
rect 33180 59714 33236 59724
rect 27916 59390 27918 59442
rect 27970 59390 27972 59442
rect 27916 59378 27972 59390
rect 26908 59266 26964 59276
rect 29932 59332 29988 59342
rect 30156 59332 30212 59342
rect 29932 59330 30100 59332
rect 29932 59278 29934 59330
rect 29986 59278 30100 59330
rect 29932 59276 30100 59278
rect 29932 59266 29988 59276
rect 26684 59166 26686 59218
rect 26738 59166 26740 59218
rect 26684 59154 26740 59166
rect 28028 59220 28084 59230
rect 28028 59126 28084 59164
rect 28140 59218 28196 59230
rect 28140 59166 28142 59218
rect 28194 59166 28196 59218
rect 26796 59106 26852 59118
rect 26796 59054 26798 59106
rect 26850 59054 26852 59106
rect 26796 58548 26852 59054
rect 27244 59106 27300 59118
rect 27244 59054 27246 59106
rect 27298 59054 27300 59106
rect 27244 58772 27300 59054
rect 27244 58706 27300 58716
rect 27692 58884 27748 58894
rect 26796 58482 26852 58492
rect 26908 58660 26964 58670
rect 25452 58434 25508 58446
rect 25452 58382 25454 58434
rect 25506 58382 25508 58434
rect 25452 58324 25508 58382
rect 25900 58436 25956 58446
rect 25900 58342 25956 58380
rect 26460 58436 26516 58446
rect 25452 58258 25508 58268
rect 26348 58324 26404 58334
rect 26348 58230 26404 58268
rect 25564 57540 25620 57550
rect 26012 57540 26068 57550
rect 25564 57446 25620 57484
rect 25900 57538 26068 57540
rect 25900 57486 26014 57538
rect 26066 57486 26068 57538
rect 25900 57484 26068 57486
rect 25788 56980 25844 56990
rect 25788 56886 25844 56924
rect 25564 55972 25620 55982
rect 25452 55970 25620 55972
rect 25452 55918 25566 55970
rect 25618 55918 25620 55970
rect 25452 55916 25620 55918
rect 25452 55636 25508 55916
rect 25564 55906 25620 55916
rect 25452 54964 25508 55580
rect 25564 55412 25620 55422
rect 25564 55318 25620 55356
rect 25900 55188 25956 57484
rect 26012 57474 26068 57484
rect 26348 57204 26404 57214
rect 26124 57092 26180 57102
rect 26124 56978 26180 57036
rect 26124 56926 26126 56978
rect 26178 56926 26180 56978
rect 26124 56914 26180 56926
rect 26236 56082 26292 56094
rect 26236 56030 26238 56082
rect 26290 56030 26292 56082
rect 26236 55412 26292 56030
rect 26236 55346 26292 55356
rect 25452 54898 25508 54908
rect 25564 55132 25956 55188
rect 26012 55298 26068 55310
rect 26012 55246 26014 55298
rect 26066 55246 26068 55298
rect 25340 54684 25508 54740
rect 24892 52110 24894 52162
rect 24946 52110 24948 52162
rect 24332 51326 24334 51378
rect 24386 51326 24388 51378
rect 24220 49026 24276 49038
rect 24220 48974 24222 49026
rect 24274 48974 24276 49026
rect 24220 48916 24276 48974
rect 24220 48850 24276 48860
rect 24108 48738 24164 48748
rect 23996 48692 24052 48702
rect 23996 48242 24052 48636
rect 23996 48190 23998 48242
rect 24050 48190 24052 48242
rect 23996 48178 24052 48190
rect 24332 48132 24388 51326
rect 24556 51380 24612 51390
rect 24612 51324 24724 51380
rect 24556 51286 24612 51324
rect 24444 51266 24500 51278
rect 24444 51214 24446 51266
rect 24498 51214 24500 51266
rect 24444 50596 24500 51214
rect 24556 50596 24612 50606
rect 24444 50594 24612 50596
rect 24444 50542 24558 50594
rect 24610 50542 24612 50594
rect 24444 50540 24612 50542
rect 24556 50530 24612 50540
rect 24668 49252 24724 51324
rect 24892 51156 24948 52110
rect 25004 52108 25172 52164
rect 25340 53506 25396 53518
rect 25340 53454 25342 53506
rect 25394 53454 25396 53506
rect 25340 52388 25396 53454
rect 25004 51604 25060 52108
rect 25004 51538 25060 51548
rect 25116 51938 25172 51950
rect 25116 51886 25118 51938
rect 25170 51886 25172 51938
rect 25004 51380 25060 51390
rect 25116 51380 25172 51886
rect 25228 51940 25284 51950
rect 25228 51846 25284 51884
rect 25340 51716 25396 52332
rect 25004 51378 25172 51380
rect 25004 51326 25006 51378
rect 25058 51326 25172 51378
rect 25004 51324 25172 51326
rect 25228 51660 25396 51716
rect 25004 51314 25060 51324
rect 24892 51100 25060 51156
rect 24892 50594 24948 50606
rect 24892 50542 24894 50594
rect 24946 50542 24948 50594
rect 24780 49700 24836 49710
rect 24780 49606 24836 49644
rect 24668 49186 24724 49196
rect 24892 49138 24948 50542
rect 25004 50370 25060 51100
rect 25116 50484 25172 50522
rect 25116 50418 25172 50428
rect 25004 50318 25006 50370
rect 25058 50318 25060 50370
rect 25004 50306 25060 50318
rect 24892 49086 24894 49138
rect 24946 49086 24948 49138
rect 24892 49074 24948 49086
rect 25004 49252 25060 49262
rect 25228 49252 25284 51660
rect 25452 50428 25508 54684
rect 24780 49026 24836 49038
rect 24780 48974 24782 49026
rect 24834 48974 24836 49026
rect 24444 48132 24500 48142
rect 24332 48076 24444 48132
rect 24444 48038 24500 48076
rect 24780 48132 24836 48974
rect 25004 49026 25060 49196
rect 25004 48974 25006 49026
rect 25058 48974 25060 49026
rect 25004 48962 25060 48974
rect 25116 49196 25284 49252
rect 25340 50372 25508 50428
rect 25564 54180 25620 55132
rect 26012 55076 26068 55246
rect 25676 54404 25732 54414
rect 25676 54402 25844 54404
rect 25676 54350 25678 54402
rect 25730 54350 25844 54402
rect 25676 54348 25844 54350
rect 25676 54338 25732 54348
rect 25564 50428 25620 54124
rect 25676 53506 25732 53518
rect 25676 53454 25678 53506
rect 25730 53454 25732 53506
rect 25676 53396 25732 53454
rect 25676 53330 25732 53340
rect 25676 53060 25732 53070
rect 25788 53060 25844 54348
rect 26012 53844 26068 55020
rect 26012 53778 26068 53788
rect 26124 54402 26180 54414
rect 26124 54350 26126 54402
rect 26178 54350 26180 54402
rect 25732 53004 25844 53060
rect 25900 53396 25956 53406
rect 25676 52834 25732 53004
rect 25676 52782 25678 52834
rect 25730 52782 25732 52834
rect 25676 52164 25732 52782
rect 25676 52098 25732 52108
rect 25900 51490 25956 53340
rect 26124 52612 26180 54350
rect 26236 53732 26292 53742
rect 26348 53732 26404 57148
rect 26460 56306 26516 58380
rect 26908 58434 26964 58604
rect 27356 58548 27412 58558
rect 27356 58454 27412 58492
rect 26908 58382 26910 58434
rect 26962 58382 26964 58434
rect 26908 58370 26964 58382
rect 27132 58322 27188 58334
rect 27132 58270 27134 58322
rect 27186 58270 27188 58322
rect 27132 57988 27188 58270
rect 27468 58324 27524 58334
rect 27468 58230 27524 58268
rect 27132 57922 27188 57932
rect 26572 57092 26628 57102
rect 26572 56978 26628 57036
rect 26572 56926 26574 56978
rect 26626 56926 26628 56978
rect 26572 56914 26628 56926
rect 26460 56254 26462 56306
rect 26514 56254 26516 56306
rect 26460 56242 26516 56254
rect 27020 56642 27076 56654
rect 27020 56590 27022 56642
rect 27074 56590 27076 56642
rect 27020 56532 27076 56590
rect 26572 56082 26628 56094
rect 26572 56030 26574 56082
rect 26626 56030 26628 56082
rect 26460 55300 26516 55310
rect 26460 55206 26516 55244
rect 26572 55076 26628 56030
rect 26572 55010 26628 55020
rect 26796 56082 26852 56094
rect 26796 56030 26798 56082
rect 26850 56030 26852 56082
rect 26684 54740 26740 54750
rect 26796 54740 26852 56030
rect 27020 55748 27076 56476
rect 27692 56308 27748 58828
rect 28140 58548 28196 59166
rect 28700 59220 28756 59230
rect 27804 58324 27860 58334
rect 27804 57762 27860 58268
rect 27916 57988 27972 57998
rect 27916 57874 27972 57932
rect 27916 57822 27918 57874
rect 27970 57822 27972 57874
rect 27916 57810 27972 57822
rect 28140 57874 28196 58492
rect 28140 57822 28142 57874
rect 28194 57822 28196 57874
rect 28140 57810 28196 57822
rect 28364 59106 28420 59118
rect 28364 59054 28366 59106
rect 28418 59054 28420 59106
rect 28364 58772 28420 59054
rect 27804 57710 27806 57762
rect 27858 57710 27860 57762
rect 27804 57698 27860 57710
rect 28364 57764 28420 58716
rect 28588 58994 28644 59006
rect 28588 58942 28590 58994
rect 28642 58942 28644 58994
rect 28588 58660 28644 58942
rect 28588 58594 28644 58604
rect 28700 58546 28756 59164
rect 29820 59218 29876 59230
rect 29820 59166 29822 59218
rect 29874 59166 29876 59218
rect 29372 59108 29428 59118
rect 29820 59108 29876 59166
rect 29372 59106 29876 59108
rect 29372 59054 29374 59106
rect 29426 59054 29876 59106
rect 29372 59052 29876 59054
rect 29372 59042 29428 59052
rect 28700 58494 28702 58546
rect 28754 58494 28756 58546
rect 28700 58482 28756 58494
rect 28812 58324 28868 58334
rect 28812 58230 28868 58268
rect 29148 58324 29204 58334
rect 28588 58210 28644 58222
rect 28588 58158 28590 58210
rect 28642 58158 28644 58210
rect 28588 57988 28644 58158
rect 28644 57932 28868 57988
rect 28588 57922 28644 57932
rect 28588 57764 28644 57774
rect 28364 57762 28644 57764
rect 28364 57710 28590 57762
rect 28642 57710 28644 57762
rect 28364 57708 28644 57710
rect 28588 57698 28644 57708
rect 28700 57652 28756 57662
rect 28700 57558 28756 57596
rect 28812 57428 28868 57932
rect 29148 57650 29204 58268
rect 29148 57598 29150 57650
rect 29202 57598 29204 57650
rect 29148 57586 29204 57598
rect 29484 58212 29540 59052
rect 29932 58996 29988 59006
rect 29484 57874 29540 58156
rect 29484 57822 29486 57874
rect 29538 57822 29540 57874
rect 28700 57372 28868 57428
rect 27916 57316 27972 57326
rect 27804 56308 27860 56318
rect 27692 56306 27860 56308
rect 27692 56254 27806 56306
rect 27858 56254 27860 56306
rect 27692 56252 27860 56254
rect 27356 55972 27412 55982
rect 27356 55878 27412 55916
rect 27020 55682 27076 55692
rect 26684 54738 26852 54740
rect 26684 54686 26686 54738
rect 26738 54686 26852 54738
rect 26684 54684 26852 54686
rect 27132 55300 27188 55310
rect 26684 54674 26740 54684
rect 27132 54626 27188 55244
rect 27132 54574 27134 54626
rect 27186 54574 27188 54626
rect 27132 54562 27188 54574
rect 27580 55298 27636 55310
rect 27580 55246 27582 55298
rect 27634 55246 27636 55298
rect 27244 54516 27300 54526
rect 27244 53732 27300 54460
rect 27468 54514 27524 54526
rect 27468 54462 27470 54514
rect 27522 54462 27524 54514
rect 27468 53732 27524 54462
rect 26236 53730 26404 53732
rect 26236 53678 26238 53730
rect 26290 53678 26404 53730
rect 26236 53676 26404 53678
rect 26236 53666 26292 53676
rect 26348 52948 26404 53676
rect 26908 53730 27300 53732
rect 26908 53678 27246 53730
rect 27298 53678 27300 53730
rect 26908 53676 27300 53678
rect 26796 53508 26852 53518
rect 26684 53506 26852 53508
rect 26684 53454 26798 53506
rect 26850 53454 26852 53506
rect 26684 53452 26852 53454
rect 26348 52882 26404 52892
rect 26460 52948 26516 52958
rect 26684 52948 26740 53452
rect 26796 53442 26852 53452
rect 26908 53170 26964 53676
rect 27244 53666 27300 53676
rect 27356 53676 27468 53732
rect 27356 53618 27412 53676
rect 27468 53666 27524 53676
rect 27580 53730 27636 55246
rect 27580 53678 27582 53730
rect 27634 53678 27636 53730
rect 27580 53666 27636 53678
rect 27692 55188 27748 56252
rect 27804 56242 27860 56252
rect 27356 53566 27358 53618
rect 27410 53566 27412 53618
rect 27356 53554 27412 53566
rect 26908 53118 26910 53170
rect 26962 53118 26964 53170
rect 26908 53106 26964 53118
rect 26460 52946 26740 52948
rect 26460 52894 26462 52946
rect 26514 52894 26740 52946
rect 26460 52892 26740 52894
rect 26796 52946 26852 52958
rect 26796 52894 26798 52946
rect 26850 52894 26852 52946
rect 26124 52546 26180 52556
rect 26348 52388 26404 52398
rect 26348 52274 26404 52332
rect 26348 52222 26350 52274
rect 26402 52222 26404 52274
rect 26348 52210 26404 52222
rect 25900 51438 25902 51490
rect 25954 51438 25956 51490
rect 25900 51426 25956 51438
rect 26012 51938 26068 51950
rect 26012 51886 26014 51938
rect 26066 51886 26068 51938
rect 25788 50482 25844 50494
rect 25788 50430 25790 50482
rect 25842 50430 25844 50482
rect 25564 50372 25732 50428
rect 24780 48066 24836 48076
rect 24892 48916 24948 48926
rect 24892 48130 24948 48860
rect 24892 48078 24894 48130
rect 24946 48078 24948 48130
rect 24668 47908 24724 47918
rect 23884 47404 24052 47460
rect 23772 47394 23828 47404
rect 23772 47236 23828 47246
rect 23660 47180 23772 47236
rect 22876 45950 22878 46002
rect 22930 45950 22932 46002
rect 22876 45444 22932 45950
rect 22876 45378 22932 45388
rect 22988 46620 23268 46676
rect 23324 46788 23380 46798
rect 22764 45164 22932 45220
rect 22652 45042 22708 45052
rect 22764 44994 22820 45006
rect 22764 44942 22766 44994
rect 22818 44942 22820 44994
rect 22540 44604 22708 44660
rect 22204 44492 22596 44548
rect 21868 44270 21870 44322
rect 21922 44270 21924 44322
rect 21868 44258 21924 44270
rect 22092 44324 22148 44362
rect 22092 44258 22148 44268
rect 22204 44322 22260 44334
rect 22204 44270 22206 44322
rect 22258 44270 22260 44322
rect 21756 44212 21812 44222
rect 21644 43540 21700 43550
rect 21644 43446 21700 43484
rect 21644 42642 21700 42654
rect 21644 42590 21646 42642
rect 21698 42590 21700 42642
rect 21644 42196 21700 42590
rect 21644 42130 21700 42140
rect 21756 42082 21812 44156
rect 22204 44212 22260 44270
rect 22204 44146 22260 44156
rect 22316 44324 22372 44334
rect 22092 44098 22148 44110
rect 22092 44046 22094 44098
rect 22146 44046 22148 44098
rect 21980 43540 22036 43550
rect 21980 42754 22036 43484
rect 22092 42978 22148 44046
rect 22092 42926 22094 42978
rect 22146 42926 22148 42978
rect 22092 42914 22148 42926
rect 21980 42702 21982 42754
rect 22034 42702 22036 42754
rect 21980 42196 22036 42702
rect 22204 42756 22260 42766
rect 22204 42662 22260 42700
rect 21980 42130 22036 42140
rect 22092 42644 22148 42654
rect 21756 42030 21758 42082
rect 21810 42030 21812 42082
rect 21532 41804 21700 41860
rect 21420 41692 21588 41748
rect 20860 41298 21028 41300
rect 20860 41246 20862 41298
rect 20914 41246 21028 41298
rect 20860 41244 21028 41246
rect 20860 41234 20916 41244
rect 20748 40402 20804 40684
rect 20972 40516 21028 41244
rect 21420 41076 21476 41086
rect 21308 40628 21364 40638
rect 21308 40534 21364 40572
rect 21420 40626 21476 41020
rect 21420 40574 21422 40626
rect 21474 40574 21476 40626
rect 21420 40562 21476 40574
rect 21532 40962 21588 41692
rect 21532 40910 21534 40962
rect 21586 40910 21588 40962
rect 20972 40450 21028 40460
rect 20748 40350 20750 40402
rect 20802 40350 20804 40402
rect 20748 40338 20804 40350
rect 21196 40404 21252 40414
rect 21196 40310 21252 40348
rect 21532 40404 21588 40910
rect 21532 40338 21588 40348
rect 21644 39844 21700 41804
rect 21756 41188 21812 42030
rect 21868 42084 21924 42094
rect 21868 41970 21924 42028
rect 21868 41918 21870 41970
rect 21922 41918 21924 41970
rect 21868 41906 21924 41918
rect 21980 41970 22036 41982
rect 21980 41918 21982 41970
rect 22034 41918 22036 41970
rect 21756 41122 21812 41132
rect 21308 39788 21700 39844
rect 21756 40740 21812 40750
rect 20972 39620 21028 39630
rect 20972 39526 21028 39564
rect 20636 38894 20638 38946
rect 20690 38894 20692 38946
rect 20524 38050 20580 38062
rect 20524 37998 20526 38050
rect 20578 37998 20580 38050
rect 20524 37044 20580 37998
rect 20524 36950 20580 36988
rect 20636 37938 20692 38894
rect 20636 37886 20638 37938
rect 20690 37886 20692 37938
rect 20412 36764 20580 36820
rect 19964 36278 20020 36316
rect 20188 36706 20244 36718
rect 20188 36654 20190 36706
rect 20242 36654 20244 36706
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 20076 35810 20132 35822
rect 20076 35758 20078 35810
rect 20130 35758 20132 35810
rect 20076 35588 20132 35758
rect 20076 35140 20132 35532
rect 20076 35074 20132 35084
rect 19180 34020 19236 34300
rect 19180 33954 19236 33964
rect 19068 33506 19124 33516
rect 18844 33294 18846 33346
rect 18898 33294 18900 33346
rect 18844 33282 18900 33294
rect 18956 33346 19012 33358
rect 18956 33294 18958 33346
rect 19010 33294 19012 33346
rect 18956 33124 19012 33294
rect 18956 32788 19012 33068
rect 18956 32722 19012 32732
rect 19404 33012 19460 34412
rect 19628 34020 19684 34860
rect 20076 34916 20132 34926
rect 20076 34822 20132 34860
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19740 34020 19796 34030
rect 19628 33964 19740 34020
rect 19740 33926 19796 33964
rect 20188 34018 20244 36654
rect 20524 36706 20580 36764
rect 20524 36654 20526 36706
rect 20578 36654 20580 36706
rect 20524 36642 20580 36654
rect 20412 36258 20468 36270
rect 20412 36206 20414 36258
rect 20466 36206 20468 36258
rect 20412 36036 20468 36206
rect 20636 36148 20692 37886
rect 20748 38724 20804 38734
rect 20748 38050 20804 38668
rect 20748 37998 20750 38050
rect 20802 37998 20804 38050
rect 20748 37716 20804 37998
rect 21196 38722 21252 38734
rect 21196 38670 21198 38722
rect 21250 38670 21252 38722
rect 20748 37660 20916 37716
rect 20748 37380 20804 37390
rect 20748 37266 20804 37324
rect 20748 37214 20750 37266
rect 20802 37214 20804 37266
rect 20748 37202 20804 37214
rect 20748 36708 20804 36718
rect 20748 36260 20804 36652
rect 20860 36484 20916 37660
rect 20972 37380 21028 37390
rect 20972 37286 21028 37324
rect 21084 37268 21140 37278
rect 21084 37174 21140 37212
rect 21196 36708 21252 38670
rect 21308 38722 21364 39788
rect 21756 39618 21812 40684
rect 21980 40628 22036 41918
rect 22092 40628 22148 42588
rect 22316 42644 22372 44268
rect 22316 42578 22372 42588
rect 22428 42756 22484 42766
rect 22428 42530 22484 42700
rect 22428 42478 22430 42530
rect 22482 42478 22484 42530
rect 22428 42466 22484 42478
rect 22316 42196 22372 42206
rect 22316 41748 22372 42140
rect 22428 41972 22484 41982
rect 22428 41878 22484 41916
rect 22316 41692 22484 41748
rect 22316 40962 22372 40974
rect 22316 40910 22318 40962
rect 22370 40910 22372 40962
rect 22316 40852 22372 40910
rect 22316 40786 22372 40796
rect 22204 40628 22260 40638
rect 22092 40572 22204 40628
rect 21980 40562 22036 40572
rect 22204 40534 22260 40572
rect 22316 40516 22372 40526
rect 21756 39566 21758 39618
rect 21810 39566 21812 39618
rect 21756 39554 21812 39566
rect 21868 40404 21924 40414
rect 21868 39506 21924 40348
rect 22316 39618 22372 40460
rect 22316 39566 22318 39618
rect 22370 39566 22372 39618
rect 22316 39554 22372 39566
rect 21868 39454 21870 39506
rect 21922 39454 21924 39506
rect 21532 38836 21588 38846
rect 21308 38670 21310 38722
rect 21362 38670 21364 38722
rect 21308 38658 21364 38670
rect 21420 38780 21532 38836
rect 21308 37380 21364 37390
rect 21420 37380 21476 38780
rect 21532 38742 21588 38780
rect 21868 38668 21924 39454
rect 21756 38612 21924 38668
rect 22092 39394 22148 39406
rect 22092 39342 22094 39394
rect 22146 39342 22148 39394
rect 21308 37378 21476 37380
rect 21308 37326 21310 37378
rect 21362 37326 21476 37378
rect 21308 37324 21476 37326
rect 21644 38050 21700 38062
rect 21644 37998 21646 38050
rect 21698 37998 21700 38050
rect 21644 37380 21700 37998
rect 21308 37314 21364 37324
rect 21644 37314 21700 37324
rect 21756 36708 21812 38612
rect 21868 38052 21924 38062
rect 21868 37958 21924 37996
rect 21868 37492 21924 37502
rect 21868 37398 21924 37436
rect 22092 37492 22148 39342
rect 22092 37360 22148 37436
rect 22428 37940 22484 41692
rect 22540 39060 22596 44492
rect 22652 41300 22708 44604
rect 22764 43764 22820 44942
rect 22764 43698 22820 43708
rect 22764 43426 22820 43438
rect 22764 43374 22766 43426
rect 22818 43374 22820 43426
rect 22764 42868 22820 43374
rect 22764 42802 22820 42812
rect 22876 41970 22932 45164
rect 22988 44324 23044 46620
rect 23324 45890 23380 46732
rect 23436 46452 23492 46844
rect 23548 46676 23604 46686
rect 23548 46582 23604 46620
rect 23436 46396 23604 46452
rect 23324 45838 23326 45890
rect 23378 45838 23380 45890
rect 23324 45826 23380 45838
rect 23100 45666 23156 45678
rect 23100 45614 23102 45666
rect 23154 45614 23156 45666
rect 23100 45556 23156 45614
rect 23212 45668 23268 45678
rect 23212 45574 23268 45612
rect 23100 45490 23156 45500
rect 22988 44258 23044 44268
rect 23212 44994 23268 45006
rect 23212 44942 23214 44994
rect 23266 44942 23268 44994
rect 23212 44212 23268 44942
rect 23548 44660 23604 46396
rect 23660 44884 23716 47180
rect 23772 47104 23828 47180
rect 23772 46788 23828 46798
rect 23772 46694 23828 46732
rect 23996 46674 24052 47404
rect 24556 47348 24612 47358
rect 24556 47254 24612 47292
rect 24332 47236 24388 47246
rect 24332 47142 24388 47180
rect 24444 47234 24500 47246
rect 24444 47182 24446 47234
rect 24498 47182 24500 47234
rect 23996 46622 23998 46674
rect 24050 46622 24052 46674
rect 23884 46562 23940 46574
rect 23884 46510 23886 46562
rect 23938 46510 23940 46562
rect 23884 46004 23940 46510
rect 23996 46228 24052 46622
rect 24220 46674 24276 46686
rect 24220 46622 24222 46674
rect 24274 46622 24276 46674
rect 24220 46452 24276 46622
rect 24444 46676 24500 47182
rect 24444 46610 24500 46620
rect 24220 46386 24276 46396
rect 23996 46172 24500 46228
rect 23884 45948 24388 46004
rect 24332 45890 24388 45948
rect 24332 45838 24334 45890
rect 24386 45838 24388 45890
rect 24220 45780 24276 45790
rect 23996 45444 24052 45454
rect 23996 45330 24052 45388
rect 23996 45278 23998 45330
rect 24050 45278 24052 45330
rect 23996 45266 24052 45278
rect 24108 45332 24164 45342
rect 24220 45332 24276 45724
rect 24332 45444 24388 45838
rect 24332 45378 24388 45388
rect 24444 45668 24500 46172
rect 24668 46116 24724 47852
rect 24668 46050 24724 46060
rect 24780 47234 24836 47246
rect 24780 47182 24782 47234
rect 24834 47182 24836 47234
rect 24780 46004 24836 47182
rect 24892 46788 24948 48078
rect 25116 47460 25172 49196
rect 25228 49028 25284 49038
rect 25228 48934 25284 48972
rect 25116 47394 25172 47404
rect 24892 46722 24948 46732
rect 25228 47236 25284 47246
rect 25004 46564 25060 46574
rect 25004 46562 25172 46564
rect 25004 46510 25006 46562
rect 25058 46510 25172 46562
rect 25004 46508 25172 46510
rect 25004 46498 25060 46508
rect 24780 45938 24836 45948
rect 24892 46452 24948 46462
rect 24780 45780 24836 45790
rect 24892 45780 24948 46396
rect 24780 45778 24948 45780
rect 24780 45726 24782 45778
rect 24834 45726 24948 45778
rect 24780 45724 24948 45726
rect 24780 45714 24836 45724
rect 24556 45668 24612 45678
rect 24444 45666 24612 45668
rect 24444 45614 24558 45666
rect 24610 45614 24612 45666
rect 24444 45612 24612 45614
rect 24108 45330 24276 45332
rect 24108 45278 24110 45330
rect 24162 45278 24276 45330
rect 24108 45276 24276 45278
rect 24108 45266 24164 45276
rect 23660 44818 23716 44828
rect 23772 45108 23828 45118
rect 23548 44604 23716 44660
rect 22988 44100 23044 44110
rect 22988 44098 23156 44100
rect 22988 44046 22990 44098
rect 23042 44046 23156 44098
rect 22988 44044 23156 44046
rect 22988 44034 23044 44044
rect 23100 43426 23156 44044
rect 23100 43374 23102 43426
rect 23154 43374 23156 43426
rect 23100 43204 23156 43374
rect 23100 43138 23156 43148
rect 23100 42644 23156 42654
rect 23100 42550 23156 42588
rect 23212 42420 23268 44156
rect 23548 44100 23604 44110
rect 23548 44006 23604 44044
rect 23660 43876 23716 44604
rect 23772 43988 23828 45052
rect 24220 45108 24276 45118
rect 23884 44996 23940 45006
rect 23884 44100 23940 44940
rect 24220 44660 24276 45052
rect 24332 45106 24388 45118
rect 24332 45054 24334 45106
rect 24386 45054 24388 45106
rect 24332 44884 24388 45054
rect 24332 44818 24388 44828
rect 24220 44594 24276 44604
rect 23884 44006 23940 44044
rect 23772 43922 23828 43932
rect 22876 41918 22878 41970
rect 22930 41918 22932 41970
rect 22876 41524 22932 41918
rect 22876 41458 22932 41468
rect 23100 42364 23268 42420
rect 23548 43820 23716 43876
rect 22652 41244 23044 41300
rect 22876 41076 22932 41086
rect 22764 40964 22820 40974
rect 22652 40962 22820 40964
rect 22652 40910 22766 40962
rect 22818 40910 22820 40962
rect 22652 40908 22820 40910
rect 22652 40516 22708 40908
rect 22764 40898 22820 40908
rect 22652 40422 22708 40460
rect 22876 40404 22932 41020
rect 22876 40338 22932 40348
rect 22988 40068 23044 41244
rect 23100 40516 23156 42364
rect 23436 41636 23492 41646
rect 23212 41300 23268 41310
rect 23212 41206 23268 41244
rect 23100 40460 23268 40516
rect 22876 39732 22932 39742
rect 22988 39732 23044 40012
rect 22876 39730 23044 39732
rect 22876 39678 22878 39730
rect 22930 39678 23044 39730
rect 22876 39676 23044 39678
rect 22876 39666 22932 39676
rect 23100 39172 23156 39182
rect 22652 39060 22708 39070
rect 22540 39058 23044 39060
rect 22540 39006 22654 39058
rect 22706 39006 23044 39058
rect 22540 39004 23044 39006
rect 22652 38994 22708 39004
rect 22988 38724 23044 39004
rect 23100 39058 23156 39116
rect 23100 39006 23102 39058
rect 23154 39006 23156 39058
rect 23100 38948 23156 39006
rect 23100 38882 23156 38892
rect 22988 38612 23156 38668
rect 22876 38500 22932 38510
rect 22652 38164 22708 38174
rect 22652 38070 22708 38108
rect 22764 38050 22820 38062
rect 22764 37998 22766 38050
rect 22818 37998 22820 38050
rect 22764 37940 22820 37998
rect 22428 37884 22820 37940
rect 21980 37268 22036 37278
rect 21980 37174 22036 37212
rect 22428 37266 22484 37884
rect 22876 37828 22932 38444
rect 22428 37214 22430 37266
rect 22482 37214 22484 37266
rect 21196 36652 21700 36708
rect 21756 36652 22260 36708
rect 21532 36484 21588 36494
rect 20860 36482 21588 36484
rect 20860 36430 21534 36482
rect 21586 36430 21588 36482
rect 20860 36428 21588 36430
rect 21532 36418 21588 36428
rect 20860 36260 20916 36270
rect 20748 36204 20860 36260
rect 20636 36092 20804 36148
rect 20860 36128 20916 36204
rect 20412 35970 20468 35980
rect 20300 35924 20356 35934
rect 20300 35830 20356 35868
rect 20636 35924 20692 35934
rect 20524 35700 20580 35710
rect 20524 35606 20580 35644
rect 20412 35588 20468 35598
rect 20412 35494 20468 35532
rect 20524 35028 20580 35038
rect 20524 34934 20580 34972
rect 20300 34914 20356 34926
rect 20300 34862 20302 34914
rect 20354 34862 20356 34914
rect 20300 34804 20356 34862
rect 20300 34738 20356 34748
rect 20636 34356 20692 35868
rect 20188 33966 20190 34018
rect 20242 33966 20244 34018
rect 19404 32786 19460 32956
rect 19404 32734 19406 32786
rect 19458 32734 19460 32786
rect 19404 32452 19460 32734
rect 19404 32386 19460 32396
rect 19516 33908 19572 33918
rect 18732 32172 19124 32228
rect 18508 31950 18510 32002
rect 18562 31950 18564 32002
rect 18508 31938 18564 31950
rect 18844 32004 18900 32014
rect 18284 31838 18286 31890
rect 18338 31838 18340 31890
rect 18284 31826 18340 31838
rect 18732 31780 18788 31790
rect 18732 31686 18788 31724
rect 18172 31602 18228 31612
rect 18060 31378 18116 31388
rect 17276 31266 17332 31276
rect 16716 27794 16772 27804
rect 16828 29484 16996 29540
rect 17052 30268 17220 30324
rect 17388 31220 17444 31230
rect 17052 29540 17108 30268
rect 17276 30212 17332 30222
rect 17276 30118 17332 30156
rect 16492 26852 16660 26908
rect 16492 26068 16548 26078
rect 16380 26012 16492 26068
rect 16492 25974 16548 26012
rect 16268 25342 16270 25394
rect 16322 25342 16324 25394
rect 16268 25172 16324 25342
rect 16604 25172 16660 26852
rect 16268 25106 16324 25116
rect 16492 25116 16660 25172
rect 16156 24610 16212 24622
rect 16156 24558 16158 24610
rect 16210 24558 16212 24610
rect 16156 23940 16212 24558
rect 16156 23874 16212 23884
rect 15820 20914 15988 20916
rect 15820 20862 15822 20914
rect 15874 20862 15988 20914
rect 15820 20860 15988 20862
rect 16044 23716 16100 23726
rect 16044 23042 16100 23660
rect 16044 22990 16046 23042
rect 16098 22990 16100 23042
rect 15820 20850 15876 20860
rect 15148 20750 15150 20802
rect 15202 20750 15204 20802
rect 15148 20738 15204 20750
rect 15596 20020 15652 20030
rect 15260 19906 15316 19918
rect 15260 19854 15262 19906
rect 15314 19854 15316 19906
rect 15260 19684 15316 19854
rect 15260 19618 15316 19628
rect 15596 19906 15652 19964
rect 15596 19854 15598 19906
rect 15650 19854 15652 19906
rect 15036 17390 15038 17442
rect 15090 17390 15092 17442
rect 14476 16882 14868 16884
rect 14476 16830 14478 16882
rect 14530 16830 14868 16882
rect 14476 16828 14868 16830
rect 14924 17108 14980 17118
rect 15036 17108 15092 17390
rect 15372 19234 15428 19246
rect 15372 19182 15374 19234
rect 15426 19182 15428 19234
rect 15372 17890 15428 19182
rect 15596 19012 15652 19854
rect 16044 19906 16100 22990
rect 16380 23714 16436 23726
rect 16380 23662 16382 23714
rect 16434 23662 16436 23714
rect 16380 22820 16436 23662
rect 16492 23716 16548 25116
rect 16604 24948 16660 24958
rect 16828 24948 16884 29484
rect 17052 29474 17108 29484
rect 17164 29876 17220 29886
rect 16940 29314 16996 29326
rect 16940 29262 16942 29314
rect 16994 29262 16996 29314
rect 16940 29204 16996 29262
rect 16940 29138 16996 29148
rect 16940 28754 16996 28766
rect 16940 28702 16942 28754
rect 16994 28702 16996 28754
rect 16940 28644 16996 28702
rect 16940 28578 16996 28588
rect 17164 28642 17220 29820
rect 17164 28590 17166 28642
rect 17218 28590 17220 28642
rect 17164 28578 17220 28590
rect 17388 28420 17444 31164
rect 17836 31220 17892 31230
rect 17836 31126 17892 31164
rect 18844 31218 18900 31948
rect 18844 31166 18846 31218
rect 18898 31166 18900 31218
rect 18844 31154 18900 31166
rect 19068 31892 19124 32172
rect 19068 31220 19124 31836
rect 19068 31154 19124 31164
rect 19180 32116 19236 32126
rect 18284 30884 18340 30894
rect 18172 30882 18340 30884
rect 18172 30830 18286 30882
rect 18338 30830 18340 30882
rect 18172 30828 18340 30830
rect 17500 30770 17556 30782
rect 17500 30718 17502 30770
rect 17554 30718 17556 30770
rect 17500 29652 17556 30718
rect 18172 30770 18228 30828
rect 18284 30818 18340 30828
rect 18172 30718 18174 30770
rect 18226 30718 18228 30770
rect 18172 30706 18228 30718
rect 18396 30548 18452 30558
rect 18172 30436 18228 30446
rect 18172 30210 18228 30380
rect 18172 30158 18174 30210
rect 18226 30158 18228 30210
rect 17724 30098 17780 30110
rect 17724 30046 17726 30098
rect 17778 30046 17780 30098
rect 17724 29876 17780 30046
rect 17948 29988 18004 29998
rect 17724 29810 17780 29820
rect 17836 29986 18004 29988
rect 17836 29934 17950 29986
rect 18002 29934 18004 29986
rect 17836 29932 18004 29934
rect 17500 29586 17556 29596
rect 17500 28868 17556 28878
rect 17500 28642 17556 28812
rect 17836 28756 17892 29932
rect 17948 29922 18004 29932
rect 18060 29986 18116 29998
rect 18060 29934 18062 29986
rect 18114 29934 18116 29986
rect 17948 29540 18004 29550
rect 18060 29540 18116 29934
rect 18172 29764 18228 30158
rect 18172 29698 18228 29708
rect 18396 30210 18452 30492
rect 19068 30436 19124 30446
rect 18396 30158 18398 30210
rect 18450 30158 18452 30210
rect 17948 29538 18116 29540
rect 17948 29486 17950 29538
rect 18002 29486 18116 29538
rect 17948 29484 18116 29486
rect 18172 29540 18228 29550
rect 17948 29474 18004 29484
rect 18172 29446 18228 29484
rect 18284 29202 18340 29214
rect 18284 29150 18286 29202
rect 18338 29150 18340 29202
rect 18284 28868 18340 29150
rect 18284 28802 18340 28812
rect 17836 28690 17892 28700
rect 17500 28590 17502 28642
rect 17554 28590 17556 28642
rect 17500 28578 17556 28590
rect 18172 28644 18228 28654
rect 16940 28364 17444 28420
rect 17836 28420 17892 28430
rect 17836 28418 18004 28420
rect 17836 28366 17838 28418
rect 17890 28366 18004 28418
rect 17836 28364 18004 28366
rect 16940 27524 16996 28364
rect 17836 28354 17892 28364
rect 17052 27748 17108 27758
rect 17052 27746 17220 27748
rect 17052 27694 17054 27746
rect 17106 27694 17220 27746
rect 17052 27692 17220 27694
rect 17052 27682 17108 27692
rect 16940 27468 17108 27524
rect 16940 26964 16996 26974
rect 16940 25618 16996 26908
rect 16940 25566 16942 25618
rect 16994 25566 16996 25618
rect 16940 25554 16996 25566
rect 16660 24892 16884 24948
rect 17052 24946 17108 27468
rect 17052 24894 17054 24946
rect 17106 24894 17108 24946
rect 16604 24816 16660 24892
rect 17052 24882 17108 24894
rect 17164 24164 17220 27692
rect 17948 27074 18004 28364
rect 18060 27746 18116 27758
rect 18060 27694 18062 27746
rect 18114 27694 18116 27746
rect 18060 27412 18116 27694
rect 18060 27346 18116 27356
rect 17948 27022 17950 27074
rect 18002 27022 18004 27074
rect 17948 27010 18004 27022
rect 18172 26964 18228 28588
rect 18396 28196 18452 30158
rect 18732 30324 18788 30334
rect 18396 28130 18452 28140
rect 18508 28868 18564 28878
rect 18508 27970 18564 28812
rect 18620 28644 18676 28654
rect 18620 28530 18676 28588
rect 18620 28478 18622 28530
rect 18674 28478 18676 28530
rect 18620 28466 18676 28478
rect 18732 28308 18788 30268
rect 18844 29316 18900 29326
rect 18844 29314 19012 29316
rect 18844 29262 18846 29314
rect 18898 29262 19012 29314
rect 18844 29260 19012 29262
rect 18844 29250 18900 29260
rect 18844 28868 18900 28878
rect 18844 28774 18900 28812
rect 18732 28242 18788 28252
rect 18844 28532 18900 28542
rect 18508 27918 18510 27970
rect 18562 27918 18564 27970
rect 18508 27906 18564 27918
rect 18620 28084 18676 28094
rect 18508 27076 18564 27086
rect 18620 27076 18676 28028
rect 18844 27746 18900 28476
rect 18844 27694 18846 27746
rect 18898 27694 18900 27746
rect 18844 27682 18900 27694
rect 18956 27524 19012 29260
rect 19068 28868 19124 30380
rect 19180 30324 19236 32060
rect 19292 32002 19348 32014
rect 19292 31950 19294 32002
rect 19346 31950 19348 32002
rect 19292 30994 19348 31950
rect 19516 31780 19572 33852
rect 20188 33908 20244 33966
rect 20188 33842 20244 33852
rect 20300 34300 20692 34356
rect 20748 34356 20804 36092
rect 20860 36036 20916 36046
rect 20860 34692 20916 35980
rect 21084 35698 21140 35710
rect 21308 35700 21364 35710
rect 21084 35646 21086 35698
rect 21138 35646 21140 35698
rect 21084 35588 21140 35646
rect 21084 35522 21140 35532
rect 21196 35698 21364 35700
rect 21196 35646 21310 35698
rect 21362 35646 21364 35698
rect 21196 35644 21364 35646
rect 20972 35140 21028 35150
rect 21196 35140 21252 35644
rect 21308 35634 21364 35644
rect 21420 35700 21476 35710
rect 20972 35138 21252 35140
rect 20972 35086 20974 35138
rect 21026 35086 21252 35138
rect 20972 35084 21252 35086
rect 20972 35074 21028 35084
rect 21420 35028 21476 35644
rect 21532 35588 21588 35598
rect 21532 35494 21588 35532
rect 21532 35028 21588 35038
rect 21420 35026 21588 35028
rect 21420 34974 21534 35026
rect 21586 34974 21588 35026
rect 21420 34972 21588 34974
rect 21532 34962 21588 34972
rect 21644 34804 21700 36652
rect 21868 36482 21924 36494
rect 21868 36430 21870 36482
rect 21922 36430 21924 36482
rect 21868 36372 21924 36430
rect 21756 36258 21812 36270
rect 21756 36206 21758 36258
rect 21810 36206 21812 36258
rect 21756 35698 21812 36206
rect 21756 35646 21758 35698
rect 21810 35646 21812 35698
rect 21756 35634 21812 35646
rect 21644 34738 21700 34748
rect 20860 34626 20916 34636
rect 21420 34692 21476 34702
rect 20748 34300 21252 34356
rect 19628 33460 19684 33470
rect 20300 33460 20356 34300
rect 20636 34132 20692 34142
rect 21084 34132 21140 34142
rect 20524 34020 20580 34030
rect 19628 33366 19684 33404
rect 19964 33404 20356 33460
rect 20412 33460 20468 33470
rect 19964 33346 20020 33404
rect 19964 33294 19966 33346
rect 20018 33294 20020 33346
rect 19964 33282 20020 33294
rect 19740 33124 19796 33162
rect 19740 33058 19796 33068
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 20188 32564 20244 33404
rect 20412 33366 20468 33404
rect 20300 32676 20356 32686
rect 20300 32582 20356 32620
rect 20076 32562 20244 32564
rect 20076 32510 20190 32562
rect 20242 32510 20244 32562
rect 20076 32508 20244 32510
rect 19964 32450 20020 32462
rect 19964 32398 19966 32450
rect 20018 32398 20020 32450
rect 19964 32340 20020 32398
rect 19964 32274 20020 32284
rect 20076 32004 20132 32508
rect 20188 32498 20244 32508
rect 20524 32452 20580 33964
rect 20636 34018 20692 34076
rect 20636 33966 20638 34018
rect 20690 33966 20692 34018
rect 20636 33124 20692 33966
rect 20972 34130 21140 34132
rect 20972 34078 21086 34130
rect 21138 34078 21140 34130
rect 20972 34076 21140 34078
rect 20860 33124 20916 33134
rect 20636 33122 20916 33124
rect 20636 33070 20862 33122
rect 20914 33070 20916 33122
rect 20636 33068 20916 33070
rect 20300 32396 20580 32452
rect 20636 32900 20692 32910
rect 20076 31938 20132 31948
rect 20188 32116 20244 32126
rect 20188 31890 20244 32060
rect 20188 31838 20190 31890
rect 20242 31838 20244 31890
rect 20188 31826 20244 31838
rect 19964 31780 20020 31790
rect 19516 31778 20020 31780
rect 19516 31726 19966 31778
rect 20018 31726 20020 31778
rect 19516 31724 20020 31726
rect 19964 31714 20020 31724
rect 19292 30942 19294 30994
rect 19346 30942 19348 30994
rect 19292 30930 19348 30942
rect 19404 31556 19460 31566
rect 19404 31106 19460 31500
rect 19516 31556 19572 31566
rect 19628 31556 19684 31566
rect 19516 31554 19628 31556
rect 19516 31502 19518 31554
rect 19570 31502 19628 31554
rect 19516 31500 19628 31502
rect 19516 31490 19572 31500
rect 19404 31054 19406 31106
rect 19458 31054 19460 31106
rect 19404 30996 19460 31054
rect 19404 30930 19460 30940
rect 19516 31220 19572 31230
rect 19180 30210 19236 30268
rect 19180 30158 19182 30210
rect 19234 30158 19236 30210
rect 19180 30146 19236 30158
rect 19292 30660 19348 30670
rect 19292 29988 19348 30604
rect 19404 30548 19460 30558
rect 19404 30210 19460 30492
rect 19404 30158 19406 30210
rect 19458 30158 19460 30210
rect 19404 30146 19460 30158
rect 19180 29932 19348 29988
rect 19180 29316 19236 29932
rect 19292 29764 19348 29774
rect 19292 29538 19348 29708
rect 19516 29650 19572 31164
rect 19628 30660 19684 31500
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 20300 30994 20356 32396
rect 20524 32004 20580 32014
rect 20524 31778 20580 31948
rect 20524 31726 20526 31778
rect 20578 31726 20580 31778
rect 20524 31714 20580 31726
rect 20412 31668 20468 31678
rect 20412 31574 20468 31612
rect 20300 30942 20302 30994
rect 20354 30942 20356 30994
rect 19628 30594 19684 30604
rect 19852 30882 19908 30894
rect 19852 30830 19854 30882
rect 19906 30830 19908 30882
rect 19628 30436 19684 30446
rect 19628 30342 19684 30380
rect 19740 30210 19796 30222
rect 19740 30158 19742 30210
rect 19794 30158 19796 30210
rect 19740 30100 19796 30158
rect 19740 30034 19796 30044
rect 19852 29988 19908 30830
rect 20076 30882 20132 30894
rect 20076 30830 20078 30882
rect 20130 30830 20132 30882
rect 19852 29922 19908 29932
rect 19964 29988 20020 29998
rect 20076 29988 20132 30830
rect 20300 30772 20356 30942
rect 20300 30706 20356 30716
rect 19964 29986 20132 29988
rect 19964 29934 19966 29986
rect 20018 29934 20132 29986
rect 19964 29932 20132 29934
rect 20412 29988 20468 29998
rect 19964 29922 20020 29932
rect 20412 29894 20468 29932
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19516 29598 19518 29650
rect 19570 29598 19572 29650
rect 19516 29586 19572 29598
rect 19292 29486 19294 29538
rect 19346 29486 19348 29538
rect 19292 29474 19348 29486
rect 20412 29538 20468 29550
rect 20412 29486 20414 29538
rect 20466 29486 20468 29538
rect 20300 29426 20356 29438
rect 20300 29374 20302 29426
rect 20354 29374 20356 29426
rect 19628 29316 19684 29326
rect 19180 29260 19460 29316
rect 19068 28812 19236 28868
rect 19068 28642 19124 28654
rect 19068 28590 19070 28642
rect 19122 28590 19124 28642
rect 19068 28532 19124 28590
rect 19068 28466 19124 28476
rect 18508 27074 18676 27076
rect 18508 27022 18510 27074
rect 18562 27022 18676 27074
rect 18508 27020 18676 27022
rect 18732 27468 19012 27524
rect 18508 27010 18564 27020
rect 18172 25732 18228 26908
rect 18732 26516 18788 27468
rect 19180 27300 19236 28812
rect 19292 28642 19348 28654
rect 19292 28590 19294 28642
rect 19346 28590 19348 28642
rect 19292 27860 19348 28590
rect 19292 27794 19348 27804
rect 18732 26450 18788 26460
rect 18844 27244 19236 27300
rect 18732 26292 18788 26302
rect 18732 26198 18788 26236
rect 18620 26178 18676 26190
rect 18620 26126 18622 26178
rect 18674 26126 18676 26178
rect 18172 25676 18564 25732
rect 18172 25506 18228 25676
rect 18172 25454 18174 25506
rect 18226 25454 18228 25506
rect 18172 25442 18228 25454
rect 18396 25508 18452 25518
rect 17164 24098 17220 24108
rect 18060 24722 18116 24734
rect 18060 24670 18062 24722
rect 18114 24670 18116 24722
rect 17612 23828 17668 23838
rect 16492 23650 16548 23660
rect 16828 23716 16884 23726
rect 16828 23622 16884 23660
rect 17612 23380 17668 23772
rect 18060 23716 18116 24670
rect 18396 24610 18452 25452
rect 18396 24558 18398 24610
rect 18450 24558 18452 24610
rect 18396 24546 18452 24558
rect 18284 24052 18340 24062
rect 18284 23958 18340 23996
rect 18060 23650 18116 23660
rect 17612 23314 17668 23324
rect 17948 23380 18004 23390
rect 17948 23378 18340 23380
rect 17948 23326 17950 23378
rect 18002 23326 18340 23378
rect 17948 23324 18340 23326
rect 17948 23314 18004 23324
rect 16380 22754 16436 22764
rect 16716 23154 16772 23166
rect 16716 23102 16718 23154
rect 16770 23102 16772 23154
rect 16380 22258 16436 22270
rect 16380 22206 16382 22258
rect 16434 22206 16436 22258
rect 16044 19854 16046 19906
rect 16098 19854 16100 19906
rect 16044 19794 16100 19854
rect 16044 19742 16046 19794
rect 16098 19742 16100 19794
rect 16044 19730 16100 19742
rect 16156 21028 16212 21038
rect 16044 19236 16100 19246
rect 16156 19236 16212 20972
rect 16380 20804 16436 22206
rect 16604 21698 16660 21710
rect 16604 21646 16606 21698
rect 16658 21646 16660 21698
rect 16492 20804 16548 20814
rect 16380 20802 16548 20804
rect 16380 20750 16494 20802
rect 16546 20750 16548 20802
rect 16380 20748 16548 20750
rect 16492 20738 16548 20748
rect 16268 20578 16324 20590
rect 16268 20526 16270 20578
rect 16322 20526 16324 20578
rect 16268 19908 16324 20526
rect 16492 20020 16548 20030
rect 16492 19926 16548 19964
rect 16268 19842 16324 19852
rect 16044 19234 16212 19236
rect 16044 19182 16046 19234
rect 16098 19182 16212 19234
rect 16044 19180 16212 19182
rect 16044 19170 16100 19180
rect 15596 18946 15652 18956
rect 16268 18562 16324 18574
rect 16268 18510 16270 18562
rect 16322 18510 16324 18562
rect 16156 18452 16212 18462
rect 15372 17838 15374 17890
rect 15426 17838 15428 17890
rect 15372 17668 15428 17838
rect 15708 18340 15764 18350
rect 15484 17668 15540 17678
rect 15372 17666 15540 17668
rect 15372 17614 15486 17666
rect 15538 17614 15540 17666
rect 15372 17612 15540 17614
rect 15036 17052 15204 17108
rect 14476 16818 14532 16828
rect 14364 16270 14366 16322
rect 14418 16270 14420 16322
rect 14364 16258 14420 16270
rect 14588 16212 14644 16222
rect 14588 16118 14644 16156
rect 14924 15876 14980 17052
rect 15036 16882 15092 16894
rect 15036 16830 15038 16882
rect 15090 16830 15092 16882
rect 15036 16100 15092 16830
rect 15148 16772 15204 17052
rect 15148 16706 15204 16716
rect 15372 16100 15428 17612
rect 15484 17602 15540 17612
rect 15708 17108 15764 18284
rect 16156 17666 16212 18396
rect 16156 17614 16158 17666
rect 16210 17614 16212 17666
rect 16156 17602 16212 17614
rect 16268 17444 16324 18510
rect 16604 18452 16660 21646
rect 16716 20132 16772 23102
rect 16940 23156 16996 23166
rect 17836 23156 17892 23166
rect 16940 23062 16996 23100
rect 17276 23154 17892 23156
rect 17276 23102 17838 23154
rect 17890 23102 17892 23154
rect 17276 23100 17892 23102
rect 17276 22482 17332 23100
rect 17276 22430 17278 22482
rect 17330 22430 17332 22482
rect 17276 22418 17332 22430
rect 17612 22820 17668 22830
rect 17052 22370 17108 22382
rect 17052 22318 17054 22370
rect 17106 22318 17108 22370
rect 16716 20066 16772 20076
rect 16828 21812 16884 21822
rect 16156 17108 16212 17118
rect 15708 17106 16212 17108
rect 15708 17054 15710 17106
rect 15762 17054 16158 17106
rect 16210 17054 16212 17106
rect 15708 17052 16212 17054
rect 15708 17042 15764 17052
rect 16156 17042 16212 17052
rect 16268 16884 16324 17388
rect 16268 16818 16324 16828
rect 16380 18396 16660 18452
rect 16716 19794 16772 19806
rect 16716 19742 16718 19794
rect 16770 19742 16772 19794
rect 15036 16098 15428 16100
rect 15036 16046 15374 16098
rect 15426 16046 15428 16098
rect 15036 16044 15428 16046
rect 15036 15876 15092 15886
rect 14924 15874 15092 15876
rect 14924 15822 15038 15874
rect 15090 15822 15092 15874
rect 14924 15820 15092 15822
rect 15036 15810 15092 15820
rect 15372 15428 15428 16044
rect 16044 16100 16100 16110
rect 16380 16100 16436 18396
rect 16604 17108 16660 17118
rect 16716 17108 16772 19742
rect 16604 17106 16772 17108
rect 16604 17054 16606 17106
rect 16658 17054 16772 17106
rect 16604 17052 16772 17054
rect 16828 17108 16884 21756
rect 16940 21700 16996 21710
rect 16940 21606 16996 21644
rect 17052 21476 17108 22318
rect 17164 21476 17220 21486
rect 17052 21420 17164 21476
rect 17164 20914 17220 21420
rect 17164 20862 17166 20914
rect 17218 20862 17220 20914
rect 17164 20850 17220 20862
rect 17052 19908 17108 19918
rect 17052 18674 17108 19852
rect 17052 18622 17054 18674
rect 17106 18622 17108 18674
rect 17052 18610 17108 18622
rect 17612 18452 17668 22764
rect 17836 22484 17892 23100
rect 18172 23156 18228 23166
rect 17948 22932 18004 22942
rect 17948 22838 18004 22876
rect 17836 22428 18116 22484
rect 17948 22260 18004 22270
rect 17724 22258 18004 22260
rect 17724 22206 17950 22258
rect 18002 22206 18004 22258
rect 17724 22204 18004 22206
rect 17724 21700 17780 22204
rect 17948 22194 18004 22204
rect 17724 21634 17780 21644
rect 17836 22036 17892 22046
rect 17836 21810 17892 21980
rect 17836 21758 17838 21810
rect 17890 21758 17892 21810
rect 17836 21588 17892 21758
rect 17948 21812 18004 21822
rect 18060 21812 18116 22428
rect 18172 22036 18228 23100
rect 18172 21970 18228 21980
rect 17948 21810 18116 21812
rect 17948 21758 17950 21810
rect 18002 21758 18116 21810
rect 17948 21756 18116 21758
rect 18172 21812 18228 21822
rect 17948 21746 18004 21756
rect 17724 20804 17780 20814
rect 17724 20710 17780 20748
rect 17836 20244 17892 21532
rect 18060 21588 18116 21598
rect 18172 21588 18228 21756
rect 18060 21586 18228 21588
rect 18060 21534 18062 21586
rect 18114 21534 18228 21586
rect 18060 21532 18228 21534
rect 18284 21588 18340 23324
rect 18508 23268 18564 25676
rect 18620 25620 18676 26126
rect 18620 25554 18676 25564
rect 18732 24948 18788 24958
rect 18732 24834 18788 24892
rect 18732 24782 18734 24834
rect 18786 24782 18788 24834
rect 18732 24770 18788 24782
rect 18732 24052 18788 24062
rect 18844 24052 18900 27244
rect 19404 27076 19460 29260
rect 19628 29222 19684 29260
rect 20300 29316 20356 29374
rect 20300 29250 20356 29260
rect 20300 28532 20356 28542
rect 19740 28420 19796 28430
rect 19292 27020 19460 27076
rect 19516 28418 19796 28420
rect 19516 28366 19742 28418
rect 19794 28366 19796 28418
rect 19516 28364 19796 28366
rect 18956 26962 19012 26974
rect 18956 26910 18958 26962
rect 19010 26910 19012 26962
rect 18956 26628 19012 26910
rect 18956 26562 19012 26572
rect 19180 26964 19236 26974
rect 19068 26292 19124 26302
rect 19068 25618 19124 26236
rect 19068 25566 19070 25618
rect 19122 25566 19124 25618
rect 18732 24050 18900 24052
rect 18732 23998 18734 24050
rect 18786 23998 18900 24050
rect 18732 23996 18900 23998
rect 18956 25060 19012 25070
rect 18732 23986 18788 23996
rect 18956 23828 19012 25004
rect 18508 23174 18564 23212
rect 18732 23772 19012 23828
rect 19068 24052 19124 25566
rect 18732 23156 18788 23772
rect 18620 23100 18788 23156
rect 18956 23268 19012 23278
rect 18620 23044 18676 23100
rect 18508 22988 18676 23044
rect 18956 23042 19012 23212
rect 18956 22990 18958 23042
rect 19010 22990 19012 23042
rect 18396 22820 18452 22830
rect 18396 22370 18452 22764
rect 18396 22318 18398 22370
rect 18450 22318 18452 22370
rect 18396 22306 18452 22318
rect 18508 21588 18564 22988
rect 18732 22932 18788 22942
rect 18732 22482 18788 22876
rect 18732 22430 18734 22482
rect 18786 22430 18788 22482
rect 18620 21812 18676 21822
rect 18732 21812 18788 22430
rect 18620 21810 18788 21812
rect 18620 21758 18622 21810
rect 18674 21758 18788 21810
rect 18620 21756 18788 21758
rect 18620 21746 18676 21756
rect 18844 21700 18900 21710
rect 18340 21532 18452 21588
rect 18508 21532 18676 21588
rect 18060 21522 18116 21532
rect 18284 21522 18340 21532
rect 18284 21140 18340 21150
rect 18060 20916 18116 20926
rect 18060 20822 18116 20860
rect 18284 20580 18340 21084
rect 17836 20242 18004 20244
rect 17836 20190 17838 20242
rect 17890 20190 18004 20242
rect 17836 20188 18004 20190
rect 17836 20178 17892 20188
rect 17836 18452 17892 18462
rect 17612 18450 17892 18452
rect 17612 18398 17838 18450
rect 17890 18398 17892 18450
rect 17612 18396 17892 18398
rect 17836 18386 17892 18396
rect 17948 18340 18004 20188
rect 18284 20130 18340 20524
rect 18284 20078 18286 20130
rect 18338 20078 18340 20130
rect 18284 20066 18340 20078
rect 18396 19684 18452 21532
rect 18508 20578 18564 20590
rect 18508 20526 18510 20578
rect 18562 20526 18564 20578
rect 18508 19908 18564 20526
rect 18508 19842 18564 19852
rect 17948 18274 18004 18284
rect 18284 19010 18340 19022
rect 18284 18958 18286 19010
rect 18338 18958 18340 19010
rect 16604 17042 16660 17052
rect 16828 17042 16884 17052
rect 17724 18226 17780 18238
rect 17724 18174 17726 18226
rect 17778 18174 17780 18226
rect 17724 17106 17780 18174
rect 17724 17054 17726 17106
rect 17778 17054 17780 17106
rect 17724 17042 17780 17054
rect 18060 17108 18116 17118
rect 18060 17014 18116 17052
rect 17052 16996 17108 17006
rect 17052 16902 17108 16940
rect 16044 16098 16436 16100
rect 16044 16046 16046 16098
rect 16098 16046 16436 16098
rect 16044 16044 16436 16046
rect 17948 16884 18004 16894
rect 16044 16034 16100 16044
rect 15260 15316 15316 15326
rect 15260 15148 15316 15260
rect 14140 14690 14196 14700
rect 15148 15092 15316 15148
rect 14028 14644 14084 14654
rect 13692 14590 13694 14642
rect 13746 14590 13748 14642
rect 13692 14578 13748 14590
rect 13804 14642 14084 14644
rect 13804 14590 14030 14642
rect 14082 14590 14084 14642
rect 13804 14588 14084 14590
rect 13692 13972 13748 13982
rect 13804 13972 13860 14588
rect 14028 14578 14084 14588
rect 14476 14308 14532 14318
rect 14924 14308 14980 14318
rect 14476 14306 14980 14308
rect 14476 14254 14478 14306
rect 14530 14254 14926 14306
rect 14978 14254 14980 14306
rect 14476 14252 14980 14254
rect 14476 14242 14532 14252
rect 13692 13970 13860 13972
rect 13692 13918 13694 13970
rect 13746 13918 13860 13970
rect 13692 13916 13860 13918
rect 13580 13076 13636 13086
rect 13692 13076 13748 13916
rect 14924 13634 14980 14252
rect 14924 13582 14926 13634
rect 14978 13582 14980 13634
rect 14252 13524 14308 13534
rect 14252 13430 14308 13468
rect 13580 13074 13692 13076
rect 13580 13022 13582 13074
rect 13634 13022 13692 13074
rect 13580 13020 13692 13022
rect 13580 13010 13636 13020
rect 13692 12944 13748 13020
rect 13916 13076 13972 13086
rect 13468 12796 13860 12852
rect 11116 11454 11118 11506
rect 11170 11454 11172 11506
rect 10556 11442 10612 11452
rect 10332 11396 10388 11406
rect 10332 11302 10388 11340
rect 11116 11396 11172 11454
rect 11116 11330 11172 11340
rect 11228 12180 11284 12190
rect 11676 12180 11732 12190
rect 11228 12178 11732 12180
rect 11228 12126 11230 12178
rect 11282 12126 11678 12178
rect 11730 12126 11732 12178
rect 11228 12124 11732 12126
rect 9100 10782 9102 10834
rect 9154 10782 9156 10834
rect 9100 10770 9156 10782
rect 9660 11282 9716 11294
rect 9660 11230 9662 11282
rect 9714 11230 9716 11282
rect 9660 10724 9716 11230
rect 9660 10658 9716 10668
rect 9996 10722 10052 10734
rect 9996 10670 9998 10722
rect 10050 10670 10052 10722
rect 8428 9938 8708 9940
rect 8428 9886 8430 9938
rect 8482 9886 8708 9938
rect 8428 9884 8708 9886
rect 8316 9266 8372 9278
rect 8316 9214 8318 9266
rect 8370 9214 8372 9266
rect 8316 9156 8372 9214
rect 8428 9268 8484 9884
rect 9548 9826 9604 9838
rect 9548 9774 9550 9826
rect 9602 9774 9604 9826
rect 8876 9602 8932 9614
rect 8876 9550 8878 9602
rect 8930 9550 8932 9602
rect 8876 9268 8932 9550
rect 8988 9268 9044 9278
rect 8876 9266 9044 9268
rect 8876 9214 8990 9266
rect 9042 9214 9044 9266
rect 8876 9212 9044 9214
rect 8428 9202 8484 9212
rect 8988 9202 9044 9212
rect 8316 9090 8372 9100
rect 9548 9044 9604 9774
rect 9884 9828 9940 9838
rect 9884 9734 9940 9772
rect 8988 8708 9044 8718
rect 7756 8372 7812 8382
rect 7756 8258 7812 8316
rect 7756 8206 7758 8258
rect 7810 8206 7812 8258
rect 7756 8194 7812 8206
rect 8092 8370 8148 8382
rect 8204 8372 8372 8428
rect 8092 8318 8094 8370
rect 8146 8318 8148 8370
rect 7980 8036 8036 8046
rect 7980 7942 8036 7980
rect 8092 7362 8148 8318
rect 8316 8260 8372 8372
rect 8204 8204 8484 8260
rect 8204 8146 8260 8204
rect 8204 8094 8206 8146
rect 8258 8094 8260 8146
rect 8204 8082 8260 8094
rect 8428 8036 8484 8204
rect 8652 8036 8708 8046
rect 8428 8034 8708 8036
rect 8428 7982 8654 8034
rect 8706 7982 8708 8034
rect 8428 7980 8708 7982
rect 8092 7310 8094 7362
rect 8146 7310 8148 7362
rect 8092 7298 8148 7310
rect 8316 7474 8372 7486
rect 8316 7422 8318 7474
rect 8370 7422 8372 7474
rect 8316 7252 8372 7422
rect 8316 7186 8372 7196
rect 8540 7252 8596 7262
rect 7644 6560 7700 6636
rect 8316 6692 8372 6702
rect 7196 6514 7252 6524
rect 7980 6468 8036 6478
rect 7980 6374 8036 6412
rect 6076 4338 6356 4340
rect 6076 4286 6078 4338
rect 6130 4286 6356 4338
rect 6076 4284 6356 4286
rect 6636 4844 6804 4900
rect 7308 6132 7364 6142
rect 6076 4274 6132 4284
rect 5740 3714 5796 3724
rect 6636 3668 6692 4844
rect 6748 3668 6804 3678
rect 6636 3666 6804 3668
rect 6636 3614 6750 3666
rect 6802 3614 6804 3666
rect 6636 3612 6804 3614
rect 6748 3602 6804 3612
rect 7308 3666 7364 6076
rect 8316 6130 8372 6636
rect 8540 6690 8596 7196
rect 8540 6638 8542 6690
rect 8594 6638 8596 6690
rect 8540 6626 8596 6638
rect 8316 6078 8318 6130
rect 8370 6078 8372 6130
rect 8316 6020 8372 6078
rect 8652 6132 8708 7980
rect 8988 7586 9044 8652
rect 8988 7534 8990 7586
rect 9042 7534 9044 7586
rect 8988 7522 9044 7534
rect 9548 8258 9604 8988
rect 9772 9042 9828 9054
rect 9772 8990 9774 9042
rect 9826 8990 9828 9042
rect 9772 8708 9828 8990
rect 9772 8642 9828 8652
rect 9996 8428 10052 10670
rect 10332 10724 10388 10734
rect 10332 10630 10388 10668
rect 9548 8206 9550 8258
rect 9602 8206 9604 8258
rect 9548 7476 9604 8206
rect 9884 8372 10052 8428
rect 10108 9154 10164 9166
rect 10108 9102 10110 9154
rect 10162 9102 10164 9154
rect 10108 8428 10164 9102
rect 11004 9156 11060 9166
rect 11004 9062 11060 9100
rect 10556 9044 10612 9054
rect 10556 8950 10612 8988
rect 10108 8372 10276 8428
rect 9884 8258 9940 8372
rect 9884 8206 9886 8258
rect 9938 8206 9940 8258
rect 9884 8194 9940 8206
rect 9660 7476 9716 7486
rect 9548 7474 9716 7476
rect 9548 7422 9662 7474
rect 9714 7422 9716 7474
rect 9548 7420 9716 7422
rect 8876 6692 8932 6702
rect 8876 6598 8932 6636
rect 9548 6692 9604 6702
rect 9660 6692 9716 7420
rect 10220 7474 10276 8372
rect 10220 7422 10222 7474
rect 10274 7422 10276 7474
rect 10220 7410 10276 7422
rect 9604 6636 9716 6692
rect 9548 6560 9604 6636
rect 8652 6066 8708 6076
rect 9100 6132 9156 6142
rect 9100 6038 9156 6076
rect 8372 5964 8484 6020
rect 8316 5888 8372 5964
rect 8316 5124 8372 5134
rect 8316 5030 8372 5068
rect 8428 4562 8484 5964
rect 8428 4510 8430 4562
rect 8482 4510 8484 4562
rect 8428 4498 8484 4510
rect 9660 5796 9716 6636
rect 9996 6692 10052 6702
rect 9996 6598 10052 6636
rect 10220 6132 10276 6142
rect 10108 5906 10164 5918
rect 10108 5854 10110 5906
rect 10162 5854 10164 5906
rect 10108 5796 10164 5854
rect 9660 5794 10164 5796
rect 9660 5742 9662 5794
rect 9714 5742 10164 5794
rect 9660 5740 10164 5742
rect 9660 5234 9716 5740
rect 10220 5684 10276 6076
rect 9660 5182 9662 5234
rect 9714 5182 9716 5234
rect 9100 4340 9156 4350
rect 9100 4246 9156 4284
rect 7308 3614 7310 3666
rect 7362 3614 7364 3666
rect 7308 3602 7364 3614
rect 7644 4228 7700 4238
rect 7644 3666 7700 4172
rect 7644 3614 7646 3666
rect 7698 3614 7700 3666
rect 5852 3556 5908 3566
rect 5068 3554 5908 3556
rect 5068 3502 5070 3554
rect 5122 3502 5854 3554
rect 5906 3502 5908 3554
rect 5068 3500 5908 3502
rect 5068 3490 5124 3500
rect 5852 3490 5908 3500
rect 6300 3556 6356 3566
rect 6300 3462 6356 3500
rect 7644 3556 7700 3614
rect 9660 3666 9716 5182
rect 10108 5628 10276 5684
rect 10780 5906 10836 5918
rect 10780 5854 10782 5906
rect 10834 5854 10836 5906
rect 10780 5684 10836 5854
rect 9772 4340 9828 4350
rect 9772 4246 9828 4284
rect 9660 3614 9662 3666
rect 9714 3614 9716 3666
rect 9660 3602 9716 3614
rect 10108 3666 10164 5628
rect 10780 5618 10836 5628
rect 10220 4228 10276 4238
rect 10220 4134 10276 4172
rect 11228 4116 11284 12124
rect 11676 12114 11732 12124
rect 13132 11732 13188 11742
rect 11676 11618 11732 11630
rect 11676 11566 11678 11618
rect 11730 11566 11732 11618
rect 11676 11506 11732 11566
rect 11676 11454 11678 11506
rect 11730 11454 11732 11506
rect 11676 11442 11732 11454
rect 12908 11396 12964 11406
rect 12460 9604 12516 9614
rect 12460 9510 12516 9548
rect 12908 8372 12964 11340
rect 13020 10052 13076 10062
rect 13020 9958 13076 9996
rect 13132 9828 13188 11676
rect 13580 10612 13636 10622
rect 13580 10518 13636 10556
rect 13020 9268 13076 9278
rect 13132 9268 13188 9772
rect 13020 9266 13188 9268
rect 13020 9214 13022 9266
rect 13074 9214 13188 9266
rect 13020 9212 13188 9214
rect 13580 9602 13636 9614
rect 13580 9550 13582 9602
rect 13634 9550 13636 9602
rect 13020 9202 13076 9212
rect 13580 9044 13636 9550
rect 13356 8932 13412 8942
rect 13356 8838 13412 8876
rect 13020 8372 13076 8382
rect 12908 8370 13076 8372
rect 12908 8318 13022 8370
rect 13074 8318 13076 8370
rect 12908 8316 13076 8318
rect 13020 8306 13076 8316
rect 12460 8034 12516 8046
rect 12460 7982 12462 8034
rect 12514 7982 12516 8034
rect 12460 7700 12516 7982
rect 13580 8034 13636 8988
rect 13580 7982 13582 8034
rect 13634 7982 13636 8034
rect 12796 7700 12852 7710
rect 12460 7698 12852 7700
rect 12460 7646 12798 7698
rect 12850 7646 12852 7698
rect 12460 7644 12852 7646
rect 12460 6468 12516 6478
rect 12796 6468 12852 7644
rect 13356 7700 13412 7710
rect 13356 7252 13412 7644
rect 13356 7186 13412 7196
rect 13580 6802 13636 7982
rect 13804 7700 13860 12796
rect 13916 9940 13972 13020
rect 14588 13076 14644 13086
rect 14588 12982 14644 13020
rect 14140 12740 14196 12750
rect 14028 10610 14084 10622
rect 14028 10558 14030 10610
rect 14082 10558 14084 10610
rect 14028 10500 14084 10558
rect 14140 10612 14196 12684
rect 14924 12740 14980 13582
rect 14924 12674 14980 12684
rect 15148 12290 15204 15092
rect 15372 14530 15428 15372
rect 16604 15428 16660 15438
rect 16604 15334 16660 15372
rect 17612 15428 17668 15438
rect 17612 15334 17668 15372
rect 15372 14478 15374 14530
rect 15426 14478 15428 14530
rect 15372 13636 15428 14478
rect 16044 14532 16100 14570
rect 16044 14466 16100 14476
rect 17948 14532 18004 16828
rect 18284 16212 18340 18958
rect 18396 18788 18452 19628
rect 18396 18732 18564 18788
rect 18396 18338 18452 18350
rect 18396 18286 18398 18338
rect 18450 18286 18452 18338
rect 18396 16324 18452 18286
rect 18508 18228 18564 18732
rect 18508 18096 18564 18172
rect 18396 16258 18452 16268
rect 18508 17444 18564 17454
rect 18284 15986 18340 16156
rect 18284 15934 18286 15986
rect 18338 15934 18340 15986
rect 18284 15922 18340 15934
rect 18508 15764 18564 17388
rect 18620 16660 18676 21532
rect 18844 21586 18900 21644
rect 18844 21534 18846 21586
rect 18898 21534 18900 21586
rect 18732 21474 18788 21486
rect 18732 21422 18734 21474
rect 18786 21422 18788 21474
rect 18732 21028 18788 21422
rect 18732 20962 18788 20972
rect 18844 20356 18900 21534
rect 18732 20300 18900 20356
rect 18732 19908 18788 20300
rect 18956 20244 19012 22990
rect 19068 20914 19124 23996
rect 19180 24050 19236 26908
rect 19292 24836 19348 27020
rect 19516 26964 19572 28364
rect 19740 28354 19796 28364
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19404 26908 19572 26964
rect 19852 27860 19908 27870
rect 19404 25060 19460 26908
rect 19852 26850 19908 27804
rect 20300 27858 20356 28476
rect 20412 28420 20468 29486
rect 20524 29314 20580 29326
rect 20524 29262 20526 29314
rect 20578 29262 20580 29314
rect 20524 28868 20580 29262
rect 20636 28980 20692 32844
rect 20860 32788 20916 33068
rect 20860 32722 20916 32732
rect 20748 32674 20804 32686
rect 20748 32622 20750 32674
rect 20802 32622 20804 32674
rect 20748 31892 20804 32622
rect 20972 32116 21028 34076
rect 21084 34066 21140 34076
rect 21084 33572 21140 33582
rect 21084 32562 21140 33516
rect 21084 32510 21086 32562
rect 21138 32510 21140 32562
rect 21084 32498 21140 32510
rect 20972 32050 21028 32060
rect 20748 31826 20804 31836
rect 20860 30324 20916 30334
rect 20860 29986 20916 30268
rect 20860 29934 20862 29986
rect 20914 29934 20916 29986
rect 20860 29092 20916 29934
rect 21084 29316 21140 29326
rect 21084 29222 21140 29260
rect 20860 29036 21140 29092
rect 20636 28924 20916 28980
rect 20524 28812 20692 28868
rect 20524 28644 20580 28654
rect 20524 28550 20580 28588
rect 20412 28354 20468 28364
rect 20300 27806 20302 27858
rect 20354 27806 20356 27858
rect 20300 27794 20356 27806
rect 19964 27746 20020 27758
rect 19964 27694 19966 27746
rect 20018 27694 20020 27746
rect 19964 27636 20020 27694
rect 19964 27570 20020 27580
rect 20636 26908 20692 28812
rect 20860 28084 20916 28924
rect 20972 28642 21028 28654
rect 20972 28590 20974 28642
rect 21026 28590 21028 28642
rect 20972 28420 21028 28590
rect 20972 28354 21028 28364
rect 20860 28082 21028 28084
rect 20860 28030 20862 28082
rect 20914 28030 21028 28082
rect 20860 28028 21028 28030
rect 20860 28018 20916 28028
rect 20860 27188 20916 27198
rect 20860 26964 20916 27132
rect 20636 26852 20804 26908
rect 20860 26898 20916 26908
rect 19852 26798 19854 26850
rect 19906 26798 19908 26850
rect 19852 26786 19908 26798
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19964 26516 20020 26526
rect 19404 24994 19460 25004
rect 19628 25732 19684 25742
rect 19628 24948 19684 25676
rect 19964 25620 20020 26460
rect 20076 26180 20132 26190
rect 20076 26086 20132 26124
rect 20076 25620 20132 25630
rect 19964 25618 20132 25620
rect 19964 25566 20078 25618
rect 20130 25566 20132 25618
rect 19964 25564 20132 25566
rect 20076 25284 20132 25564
rect 20076 25228 20244 25284
rect 20188 25172 20244 25228
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20188 25106 20244 25116
rect 20524 25282 20580 25294
rect 20524 25230 20526 25282
rect 20578 25230 20580 25282
rect 19836 25050 20100 25060
rect 19852 24948 19908 24958
rect 19628 24946 19908 24948
rect 19628 24894 19854 24946
rect 19906 24894 19908 24946
rect 19628 24892 19908 24894
rect 19852 24882 19908 24892
rect 19292 24780 19460 24836
rect 19180 23998 19182 24050
rect 19234 23998 19236 24050
rect 19180 23986 19236 23998
rect 19292 24612 19348 24622
rect 19292 23828 19348 24556
rect 19068 20862 19070 20914
rect 19122 20862 19124 20914
rect 19068 20850 19124 20862
rect 19180 23772 19348 23828
rect 19404 23828 19460 24780
rect 20524 24612 20580 25230
rect 20748 25284 20804 26852
rect 20748 25218 20804 25228
rect 20860 26516 20916 26526
rect 20860 24948 20916 26460
rect 20972 26292 21028 28028
rect 20972 26226 21028 26236
rect 20860 24882 20916 24892
rect 20524 24546 20580 24556
rect 20860 24722 20916 24734
rect 20860 24670 20862 24722
rect 20914 24670 20916 24722
rect 19516 24500 19572 24510
rect 19516 24498 19684 24500
rect 19516 24446 19518 24498
rect 19570 24446 19684 24498
rect 19516 24444 19684 24446
rect 19516 24434 19572 24444
rect 19516 24052 19572 24062
rect 19516 23958 19572 23996
rect 19180 20692 19236 23772
rect 19404 23762 19460 23772
rect 19628 23716 19684 24444
rect 20524 24052 20580 24062
rect 19628 23650 19684 23660
rect 20188 23940 20244 23950
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19852 23380 19908 23390
rect 20188 23380 20244 23884
rect 19852 23378 20244 23380
rect 19852 23326 19854 23378
rect 19906 23326 20244 23378
rect 19852 23324 20244 23326
rect 19852 23314 19908 23324
rect 19516 23042 19572 23054
rect 19516 22990 19518 23042
rect 19570 22990 19572 23042
rect 19516 22372 19572 22990
rect 19516 22306 19572 22316
rect 20188 22484 20244 23324
rect 20188 22370 20244 22428
rect 20188 22318 20190 22370
rect 20242 22318 20244 22370
rect 19516 22146 19572 22158
rect 19516 22094 19518 22146
rect 19570 22094 19572 22146
rect 19516 21812 19572 22094
rect 19516 21746 19572 21756
rect 19628 22146 19684 22158
rect 19628 22094 19630 22146
rect 19682 22094 19684 22146
rect 19292 21588 19348 21598
rect 19628 21588 19684 22094
rect 19740 22148 19796 22186
rect 19740 22082 19796 22092
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19292 21586 19684 21588
rect 19292 21534 19294 21586
rect 19346 21534 19684 21586
rect 19292 21532 19684 21534
rect 20076 21588 20132 21598
rect 19292 21522 19348 21532
rect 20076 21494 20132 21532
rect 20188 20916 20244 22318
rect 20412 23042 20468 23054
rect 20412 22990 20414 23042
rect 20466 22990 20468 23042
rect 20412 21700 20468 22990
rect 20524 22146 20580 23996
rect 20636 23938 20692 23950
rect 20636 23886 20638 23938
rect 20690 23886 20692 23938
rect 20636 23156 20692 23886
rect 20748 23716 20804 23726
rect 20748 23622 20804 23660
rect 20636 23090 20692 23100
rect 20748 23042 20804 23054
rect 20748 22990 20750 23042
rect 20802 22990 20804 23042
rect 20748 22932 20804 22990
rect 20748 22866 20804 22876
rect 20860 22596 20916 24670
rect 20748 22540 20916 22596
rect 20524 22094 20526 22146
rect 20578 22094 20580 22146
rect 20524 21924 20580 22094
rect 20524 21858 20580 21868
rect 20636 22148 20692 22158
rect 20524 21700 20580 21710
rect 20412 21644 20524 21700
rect 19516 20804 19572 20814
rect 18844 20188 19012 20244
rect 19068 20636 19236 20692
rect 19292 20802 19572 20804
rect 19292 20750 19518 20802
rect 19570 20750 19572 20802
rect 19292 20748 19572 20750
rect 18844 20130 18900 20188
rect 18844 20078 18846 20130
rect 18898 20078 18900 20130
rect 18844 20066 18900 20078
rect 19068 19908 19124 20636
rect 18732 19852 19012 19908
rect 18732 18338 18788 18350
rect 18732 18286 18734 18338
rect 18786 18286 18788 18338
rect 18732 18226 18788 18286
rect 18732 18174 18734 18226
rect 18786 18174 18788 18226
rect 18732 18162 18788 18174
rect 18844 16996 18900 17006
rect 18844 16902 18900 16940
rect 18620 16594 18676 16604
rect 18956 16658 19012 19852
rect 19068 19842 19124 19852
rect 19180 20132 19236 20142
rect 19180 19906 19236 20076
rect 19180 19854 19182 19906
rect 19234 19854 19236 19906
rect 19068 19684 19124 19694
rect 19068 19458 19124 19628
rect 19068 19406 19070 19458
rect 19122 19406 19124 19458
rect 19068 19394 19124 19406
rect 19180 19460 19236 19854
rect 19292 19684 19348 20748
rect 19516 20738 19572 20748
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20188 20244 20244 20860
rect 19740 20020 19796 20030
rect 19516 20018 19796 20020
rect 19516 19966 19742 20018
rect 19794 19966 19796 20018
rect 19516 19964 19796 19966
rect 19292 19618 19348 19628
rect 19404 19908 19460 19918
rect 19292 19460 19348 19470
rect 19180 19458 19348 19460
rect 19180 19406 19294 19458
rect 19346 19406 19348 19458
rect 19180 19404 19348 19406
rect 19292 19394 19348 19404
rect 19404 19346 19460 19852
rect 19404 19294 19406 19346
rect 19458 19294 19460 19346
rect 19404 19282 19460 19294
rect 19180 18340 19236 18350
rect 19180 18246 19236 18284
rect 19516 17892 19572 19964
rect 19740 19954 19796 19964
rect 20188 19348 20244 20188
rect 20300 21586 20356 21598
rect 20300 21534 20302 21586
rect 20354 21534 20356 21586
rect 20300 19796 20356 21534
rect 20524 20242 20580 21644
rect 20524 20190 20526 20242
rect 20578 20190 20580 20242
rect 20524 20178 20580 20190
rect 20636 21362 20692 22092
rect 20748 22146 20804 22540
rect 20860 22372 20916 22382
rect 20860 22278 20916 22316
rect 20748 22094 20750 22146
rect 20802 22094 20804 22146
rect 20748 21700 20804 22094
rect 21084 22036 21140 29036
rect 21196 28308 21252 34300
rect 21308 34020 21364 34030
rect 21308 33926 21364 33964
rect 21308 33124 21364 33134
rect 21308 32676 21364 33068
rect 21308 32610 21364 32620
rect 21420 31218 21476 34636
rect 21420 31166 21422 31218
rect 21474 31166 21476 31218
rect 21420 31154 21476 31166
rect 21532 34130 21588 34142
rect 21532 34078 21534 34130
rect 21586 34078 21588 34130
rect 21308 30996 21364 31006
rect 21308 29426 21364 30940
rect 21532 30882 21588 34078
rect 21644 34132 21700 34142
rect 21868 34132 21924 36316
rect 22092 36484 22148 36494
rect 21980 34692 22036 34702
rect 21980 34598 22036 34636
rect 21700 34076 21924 34132
rect 21644 34038 21700 34076
rect 21644 33908 21700 33918
rect 21644 33346 21700 33852
rect 22092 33684 22148 36428
rect 22204 36370 22260 36652
rect 22204 36318 22206 36370
rect 22258 36318 22260 36370
rect 22204 36148 22260 36318
rect 22428 36372 22484 37214
rect 22428 36306 22484 36316
rect 22652 37772 22932 37828
rect 22988 37938 23044 37950
rect 22988 37886 22990 37938
rect 23042 37886 23044 37938
rect 22204 36082 22260 36092
rect 22204 35924 22260 35934
rect 22652 35924 22708 37772
rect 22764 37492 22820 37502
rect 22764 36482 22820 37436
rect 22988 37492 23044 37886
rect 22988 37426 23044 37436
rect 23100 37490 23156 38612
rect 23100 37438 23102 37490
rect 23154 37438 23156 37490
rect 23100 37426 23156 37438
rect 22764 36430 22766 36482
rect 22818 36430 22820 36482
rect 22764 36418 22820 36430
rect 22876 36260 22932 36270
rect 23100 36260 23156 36270
rect 22876 36166 22932 36204
rect 22988 36258 23156 36260
rect 22988 36206 23102 36258
rect 23154 36206 23156 36258
rect 22988 36204 23156 36206
rect 22652 35868 22820 35924
rect 22204 35830 22260 35868
rect 22652 35588 22708 35598
rect 22652 35494 22708 35532
rect 22652 35138 22708 35150
rect 22652 35086 22654 35138
rect 22706 35086 22708 35138
rect 22652 35028 22708 35086
rect 22428 35026 22708 35028
rect 22428 34974 22654 35026
rect 22706 34974 22708 35026
rect 22428 34972 22708 34974
rect 22316 34018 22372 34030
rect 22316 33966 22318 34018
rect 22370 33966 22372 34018
rect 22316 33906 22372 33966
rect 22316 33854 22318 33906
rect 22370 33854 22372 33906
rect 22316 33842 22372 33854
rect 22428 33684 22484 34972
rect 22652 34962 22708 34972
rect 22764 34356 22820 35868
rect 22652 34300 22820 34356
rect 22652 34018 22708 34300
rect 22652 33966 22654 34018
rect 22706 33966 22708 34018
rect 22092 33628 22260 33684
rect 21644 33294 21646 33346
rect 21698 33294 21700 33346
rect 21644 33282 21700 33294
rect 22092 33460 22148 33470
rect 21980 33234 22036 33246
rect 21980 33182 21982 33234
rect 22034 33182 22036 33234
rect 21868 33122 21924 33134
rect 21868 33070 21870 33122
rect 21922 33070 21924 33122
rect 21756 32676 21812 32686
rect 21756 32562 21812 32620
rect 21756 32510 21758 32562
rect 21810 32510 21812 32562
rect 21756 32498 21812 32510
rect 21868 32452 21924 33070
rect 21868 32386 21924 32396
rect 21980 32228 22036 33182
rect 22092 33234 22148 33404
rect 22092 33182 22094 33234
rect 22146 33182 22148 33234
rect 22092 33170 22148 33182
rect 22092 32788 22148 32798
rect 22092 32452 22148 32732
rect 22092 32386 22148 32396
rect 21980 32172 22148 32228
rect 21756 31892 21812 31902
rect 21756 31778 21812 31836
rect 21756 31726 21758 31778
rect 21810 31726 21812 31778
rect 21756 31714 21812 31726
rect 21980 31780 22036 31790
rect 21980 31686 22036 31724
rect 21532 30830 21534 30882
rect 21586 30830 21588 30882
rect 21532 30818 21588 30830
rect 21644 31220 21700 31230
rect 21644 30548 21700 31164
rect 21868 31108 21924 31118
rect 21868 31014 21924 31052
rect 22092 30996 22148 32172
rect 22204 31892 22260 33628
rect 22204 31826 22260 31836
rect 22316 33628 22484 33684
rect 22540 33906 22596 33918
rect 22540 33854 22542 33906
rect 22594 33854 22596 33906
rect 22540 33684 22596 33854
rect 22652 33908 22708 33966
rect 22652 33842 22708 33852
rect 22764 34020 22820 34030
rect 22540 33628 22708 33684
rect 22204 31556 22260 31566
rect 22204 31462 22260 31500
rect 22092 30930 22148 30940
rect 21644 30482 21700 30492
rect 21756 30884 21812 30894
rect 21532 29988 21588 29998
rect 21532 29894 21588 29932
rect 21308 29374 21310 29426
rect 21362 29374 21364 29426
rect 21308 29362 21364 29374
rect 21196 28242 21252 28252
rect 21308 27748 21364 27758
rect 21756 27748 21812 30828
rect 21980 30100 22036 30110
rect 21980 29540 22036 30044
rect 22316 30100 22372 33628
rect 22428 33458 22484 33470
rect 22428 33406 22430 33458
rect 22482 33406 22484 33458
rect 22428 31778 22484 33406
rect 22428 31726 22430 31778
rect 22482 31726 22484 31778
rect 22428 31714 22484 31726
rect 22540 33460 22596 33470
rect 22316 30034 22372 30044
rect 22092 29986 22148 29998
rect 22092 29934 22094 29986
rect 22146 29934 22148 29986
rect 22092 29764 22148 29934
rect 22092 29698 22148 29708
rect 22428 29876 22484 29886
rect 21980 28642 22036 29484
rect 21980 28590 21982 28642
rect 22034 28590 22036 28642
rect 21980 28578 22036 28590
rect 22428 29650 22484 29820
rect 22428 29598 22430 29650
rect 22482 29598 22484 29650
rect 22428 28756 22484 29598
rect 22204 28532 22260 28542
rect 22204 28438 22260 28476
rect 22316 28084 22372 28094
rect 22428 28084 22484 28700
rect 22316 28082 22484 28084
rect 22316 28030 22318 28082
rect 22370 28030 22484 28082
rect 22316 28028 22484 28030
rect 22316 28018 22372 28028
rect 22540 27972 22596 33404
rect 22652 31108 22708 33628
rect 22764 32674 22820 33964
rect 22876 33348 22932 33358
rect 22876 33254 22932 33292
rect 22764 32622 22766 32674
rect 22818 32622 22820 32674
rect 22764 32610 22820 32622
rect 22876 33012 22932 33022
rect 22876 32452 22932 32956
rect 22988 32786 23044 36204
rect 23100 36194 23156 36204
rect 23100 34690 23156 34702
rect 23100 34638 23102 34690
rect 23154 34638 23156 34690
rect 23100 34020 23156 34638
rect 23100 33926 23156 33964
rect 23212 33684 23268 40460
rect 23324 40402 23380 40414
rect 23324 40350 23326 40402
rect 23378 40350 23380 40402
rect 23324 39732 23380 40350
rect 23324 39666 23380 39676
rect 23324 35924 23380 35934
rect 23324 35698 23380 35868
rect 23324 35646 23326 35698
rect 23378 35646 23380 35698
rect 23324 35634 23380 35646
rect 23212 33618 23268 33628
rect 23324 33906 23380 33918
rect 23324 33854 23326 33906
rect 23378 33854 23380 33906
rect 23212 33348 23268 33358
rect 23324 33348 23380 33854
rect 23212 33346 23380 33348
rect 23212 33294 23214 33346
rect 23266 33294 23380 33346
rect 23212 33292 23380 33294
rect 23212 33282 23268 33292
rect 23100 33124 23156 33134
rect 23100 33030 23156 33068
rect 23436 32900 23492 41580
rect 23548 39844 23604 43820
rect 23996 43764 24052 43774
rect 23996 43652 24052 43708
rect 23884 43650 24052 43652
rect 23884 43598 23998 43650
rect 24050 43598 24052 43650
rect 23884 43596 24052 43598
rect 23660 43426 23716 43438
rect 23660 43374 23662 43426
rect 23714 43374 23716 43426
rect 23660 43314 23716 43374
rect 23660 43262 23662 43314
rect 23714 43262 23716 43314
rect 23660 43250 23716 43262
rect 23660 42756 23716 42766
rect 23660 42662 23716 42700
rect 23660 42420 23716 42430
rect 23660 41970 23716 42364
rect 23660 41918 23662 41970
rect 23714 41918 23716 41970
rect 23660 40740 23716 41918
rect 23772 41860 23828 41870
rect 23772 41298 23828 41804
rect 23772 41246 23774 41298
rect 23826 41246 23828 41298
rect 23772 41234 23828 41246
rect 23660 40684 23828 40740
rect 23548 39778 23604 39788
rect 23660 40404 23716 40414
rect 23548 39618 23604 39630
rect 23548 39566 23550 39618
rect 23602 39566 23604 39618
rect 23548 39060 23604 39566
rect 23548 38994 23604 39004
rect 23548 38834 23604 38846
rect 23548 38782 23550 38834
rect 23602 38782 23604 38834
rect 23548 38500 23604 38782
rect 23548 38434 23604 38444
rect 23548 37940 23604 37950
rect 23548 37490 23604 37884
rect 23548 37438 23550 37490
rect 23602 37438 23604 37490
rect 23548 37426 23604 37438
rect 23660 36932 23716 40348
rect 23772 38500 23828 40684
rect 23884 40404 23940 43596
rect 23996 43586 24052 43596
rect 24108 43428 24164 43438
rect 23996 42754 24052 42766
rect 23996 42702 23998 42754
rect 24050 42702 24052 42754
rect 23996 40628 24052 42702
rect 24108 42084 24164 43372
rect 24108 41858 24164 42028
rect 24108 41806 24110 41858
rect 24162 41806 24164 41858
rect 24108 41794 24164 41806
rect 24220 41972 24276 41982
rect 24220 41412 24276 41916
rect 24444 41636 24500 45612
rect 24556 45602 24612 45612
rect 24668 45666 24724 45678
rect 24668 45614 24670 45666
rect 24722 45614 24724 45666
rect 24668 44996 24724 45614
rect 24556 44940 24724 44996
rect 24892 45556 24948 45566
rect 24556 44546 24612 44940
rect 24556 44494 24558 44546
rect 24610 44494 24612 44546
rect 24556 44482 24612 44494
rect 24668 44548 24724 44558
rect 24668 44454 24724 44492
rect 24892 44546 24948 45500
rect 25004 45332 25060 45342
rect 25004 45238 25060 45276
rect 24892 44494 24894 44546
rect 24946 44494 24948 44546
rect 24892 44482 24948 44494
rect 25004 44772 25060 44782
rect 25004 44546 25060 44716
rect 25004 44494 25006 44546
rect 25058 44494 25060 44546
rect 25004 44482 25060 44494
rect 25116 44324 25172 46508
rect 25228 45332 25284 47180
rect 25340 46228 25396 50372
rect 25676 50036 25732 50372
rect 25676 49904 25732 49980
rect 25564 49586 25620 49598
rect 25564 49534 25566 49586
rect 25618 49534 25620 49586
rect 25452 48916 25508 48926
rect 25452 48822 25508 48860
rect 25564 47236 25620 49534
rect 25788 49364 25844 50430
rect 25676 49308 25844 49364
rect 26012 50372 26068 51886
rect 26124 51380 26180 51390
rect 26124 51286 26180 51324
rect 26460 51154 26516 52892
rect 26796 52612 26852 52894
rect 27020 52948 27076 52958
rect 27020 52854 27076 52892
rect 26796 52546 26852 52556
rect 27244 52836 27300 52846
rect 27468 52836 27524 52846
rect 27300 52834 27524 52836
rect 27300 52782 27470 52834
rect 27522 52782 27524 52834
rect 27300 52780 27524 52782
rect 26908 52052 26964 52062
rect 26460 51102 26462 51154
rect 26514 51102 26516 51154
rect 26460 50932 26516 51102
rect 26460 50866 26516 50876
rect 26796 52050 26964 52052
rect 26796 51998 26910 52050
rect 26962 51998 26964 52050
rect 26796 51996 26964 51998
rect 25676 48692 25732 49308
rect 26012 49028 26068 50316
rect 26236 50484 26292 50494
rect 26124 49698 26180 49710
rect 26124 49646 26126 49698
rect 26178 49646 26180 49698
rect 26124 49586 26180 49646
rect 26124 49534 26126 49586
rect 26178 49534 26180 49586
rect 26124 49522 26180 49534
rect 25676 48020 25732 48636
rect 25900 48972 26012 49028
rect 25788 48580 25844 48590
rect 25788 48466 25844 48524
rect 25788 48414 25790 48466
rect 25842 48414 25844 48466
rect 25788 48402 25844 48414
rect 25676 47954 25732 47964
rect 25564 47170 25620 47180
rect 25676 47460 25732 47470
rect 25676 47234 25732 47404
rect 25676 47182 25678 47234
rect 25730 47182 25732 47234
rect 25676 46900 25732 47182
rect 25900 47124 25956 48972
rect 26012 48962 26068 48972
rect 26012 48802 26068 48814
rect 26012 48750 26014 48802
rect 26066 48750 26068 48802
rect 26012 47348 26068 48750
rect 26124 47682 26180 47694
rect 26124 47630 26126 47682
rect 26178 47630 26180 47682
rect 26124 47570 26180 47630
rect 26124 47518 26126 47570
rect 26178 47518 26180 47570
rect 26124 47506 26180 47518
rect 26012 47282 26068 47292
rect 25900 47068 26180 47124
rect 25676 46834 25732 46844
rect 25900 46900 25956 46910
rect 25788 46564 25844 46574
rect 25676 46508 25788 46564
rect 25676 46450 25732 46508
rect 25788 46498 25844 46508
rect 25676 46398 25678 46450
rect 25730 46398 25732 46450
rect 25676 46386 25732 46398
rect 25340 46162 25396 46172
rect 25452 45892 25508 45930
rect 25452 45826 25508 45836
rect 25564 45778 25620 45790
rect 25564 45726 25566 45778
rect 25618 45726 25620 45778
rect 25340 45668 25396 45678
rect 25340 45574 25396 45612
rect 25564 45668 25620 45726
rect 25788 45780 25844 45790
rect 25788 45686 25844 45724
rect 25564 45602 25620 45612
rect 25228 45266 25284 45276
rect 25676 45108 25732 45146
rect 25676 45042 25732 45052
rect 25676 44882 25732 44894
rect 25676 44830 25678 44882
rect 25730 44830 25732 44882
rect 24556 44268 25172 44324
rect 25228 44660 25284 44670
rect 24556 43650 24612 44268
rect 24556 43598 24558 43650
rect 24610 43598 24612 43650
rect 24556 43540 24612 43598
rect 24556 43474 24612 43484
rect 24780 43988 24836 43998
rect 24668 42084 24724 42094
rect 24556 41748 24612 41758
rect 24556 41654 24612 41692
rect 24444 41570 24500 41580
rect 24444 41412 24500 41422
rect 24220 41410 24500 41412
rect 24220 41358 24446 41410
rect 24498 41358 24500 41410
rect 24220 41356 24500 41358
rect 24444 41346 24500 41356
rect 24668 41410 24724 42028
rect 24668 41358 24670 41410
rect 24722 41358 24724 41410
rect 24668 41346 24724 41358
rect 24332 41186 24388 41198
rect 24780 41188 24836 43932
rect 25116 43764 25172 43774
rect 25004 43426 25060 43438
rect 25004 43374 25006 43426
rect 25058 43374 25060 43426
rect 24332 41134 24334 41186
rect 24386 41134 24388 41186
rect 24332 40852 24388 41134
rect 24332 40786 24388 40796
rect 24668 41132 24836 41188
rect 24892 42644 24948 42654
rect 23996 40562 24052 40572
rect 24444 40628 24500 40638
rect 23884 40348 24276 40404
rect 23772 38434 23828 38444
rect 23884 39620 23940 39630
rect 23548 36876 23716 36932
rect 23548 34692 23604 36876
rect 23660 36706 23716 36718
rect 23660 36654 23662 36706
rect 23714 36654 23716 36706
rect 23660 36594 23716 36654
rect 23660 36542 23662 36594
rect 23714 36542 23716 36594
rect 23660 36530 23716 36542
rect 23884 35698 23940 39564
rect 23996 38948 24052 38958
rect 23996 38854 24052 38892
rect 24108 38050 24164 38062
rect 24108 37998 24110 38050
rect 24162 37998 24164 38050
rect 23996 37940 24052 37950
rect 23996 37490 24052 37884
rect 24108 37828 24164 37998
rect 24108 37762 24164 37772
rect 23996 37438 23998 37490
rect 24050 37438 24052 37490
rect 23996 37426 24052 37438
rect 24108 37042 24164 37054
rect 24108 36990 24110 37042
rect 24162 36990 24164 37042
rect 23996 36258 24052 36270
rect 23996 36206 23998 36258
rect 24050 36206 24052 36258
rect 23996 36148 24052 36206
rect 23996 36082 24052 36092
rect 23884 35646 23886 35698
rect 23938 35646 23940 35698
rect 23884 35138 23940 35646
rect 23884 35086 23886 35138
rect 23938 35086 23940 35138
rect 23884 35074 23940 35086
rect 23548 34690 23716 34692
rect 23548 34638 23550 34690
rect 23602 34638 23716 34690
rect 23548 34636 23716 34638
rect 23548 34626 23604 34636
rect 23548 34468 23604 34478
rect 23548 34354 23604 34412
rect 23548 34302 23550 34354
rect 23602 34302 23604 34354
rect 23548 34290 23604 34302
rect 22988 32734 22990 32786
rect 23042 32734 23044 32786
rect 22988 32722 23044 32734
rect 23100 32844 23492 32900
rect 23660 33906 23716 34636
rect 23660 33854 23662 33906
rect 23714 33854 23716 33906
rect 22764 32396 22932 32452
rect 22764 31332 22820 32396
rect 23100 32116 23156 32844
rect 23324 32676 23380 32686
rect 23548 32676 23604 32686
rect 23324 32674 23548 32676
rect 23324 32622 23326 32674
rect 23378 32622 23548 32674
rect 23324 32620 23548 32622
rect 23324 32610 23380 32620
rect 23548 32610 23604 32620
rect 23212 32562 23268 32574
rect 23212 32510 23214 32562
rect 23266 32510 23268 32562
rect 23212 32452 23268 32510
rect 23212 32386 23268 32396
rect 23324 32452 23380 32462
rect 23324 32450 23604 32452
rect 23324 32398 23326 32450
rect 23378 32398 23604 32450
rect 23324 32396 23604 32398
rect 23324 32386 23380 32396
rect 22988 32060 23156 32116
rect 22876 31892 22932 31902
rect 22876 31798 22932 31836
rect 22988 31668 23044 32060
rect 22764 31266 22820 31276
rect 22876 31612 23044 31668
rect 23100 31892 23156 31902
rect 22652 31052 22820 31108
rect 22652 30884 22708 30894
rect 22652 30790 22708 30828
rect 22652 30212 22708 30222
rect 22652 30118 22708 30156
rect 22764 28980 22820 31052
rect 22764 28084 22820 28924
rect 21084 21970 21140 21980
rect 21196 27746 21812 27748
rect 21196 27694 21310 27746
rect 21362 27694 21812 27746
rect 21196 27692 21812 27694
rect 22428 27916 22596 27972
rect 22652 28028 22820 28084
rect 20748 21634 20804 21644
rect 21196 21588 21252 27692
rect 21308 27682 21364 27692
rect 21756 27132 22260 27188
rect 21756 26402 21812 27132
rect 22204 27074 22260 27132
rect 22204 27022 22206 27074
rect 22258 27022 22260 27074
rect 21868 26962 21924 26974
rect 21868 26910 21870 26962
rect 21922 26910 21924 26962
rect 21868 26908 21924 26910
rect 21868 26852 22036 26908
rect 21756 26350 21758 26402
rect 21810 26350 21812 26402
rect 21756 26338 21812 26350
rect 21980 26290 22036 26852
rect 21980 26238 21982 26290
rect 22034 26238 22036 26290
rect 21868 25732 21924 25742
rect 21868 25618 21924 25676
rect 21868 25566 21870 25618
rect 21922 25566 21924 25618
rect 21868 25554 21924 25566
rect 21420 25172 21476 25182
rect 21420 24722 21476 25116
rect 21980 24834 22036 26238
rect 21980 24782 21982 24834
rect 22034 24782 22036 24834
rect 21980 24770 22036 24782
rect 22092 26292 22148 26302
rect 22092 25730 22148 26236
rect 22092 25678 22094 25730
rect 22146 25678 22148 25730
rect 21420 24670 21422 24722
rect 21474 24670 21476 24722
rect 21420 23940 21476 24670
rect 21868 24612 21924 24622
rect 21420 23874 21476 23884
rect 21756 23938 21812 23950
rect 21756 23886 21758 23938
rect 21810 23886 21812 23938
rect 21308 23156 21364 23166
rect 21308 23062 21364 23100
rect 21644 22484 21700 22494
rect 21644 22390 21700 22428
rect 21420 22372 21476 22382
rect 21308 21588 21364 21598
rect 21196 21586 21364 21588
rect 21196 21534 21310 21586
rect 21362 21534 21364 21586
rect 21196 21532 21364 21534
rect 21308 21476 21364 21532
rect 21308 21410 21364 21420
rect 20636 21310 20638 21362
rect 20690 21310 20692 21362
rect 20636 20132 20692 21310
rect 21420 20242 21476 22316
rect 21644 22036 21700 22046
rect 21420 20190 21422 20242
rect 21474 20190 21476 20242
rect 21420 20178 21476 20190
rect 21532 21924 21588 21934
rect 21308 20132 21364 20142
rect 20636 20130 21364 20132
rect 20636 20078 21310 20130
rect 21362 20078 21364 20130
rect 20636 20076 21364 20078
rect 21308 20066 21364 20076
rect 20300 19740 20580 19796
rect 20524 19458 20580 19740
rect 20524 19406 20526 19458
rect 20578 19406 20580 19458
rect 20524 19394 20580 19406
rect 20860 19458 20916 19470
rect 20860 19406 20862 19458
rect 20914 19406 20916 19458
rect 20412 19348 20468 19358
rect 20188 19346 20468 19348
rect 20188 19294 20414 19346
rect 20466 19294 20468 19346
rect 20188 19292 20468 19294
rect 19964 19012 20020 19022
rect 19628 19010 20020 19012
rect 19628 18958 19966 19010
rect 20018 18958 20020 19010
rect 19628 18956 20020 18958
rect 19628 18676 19684 18956
rect 19964 18946 20020 18956
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19628 18620 19796 18676
rect 19628 18340 19684 18350
rect 19628 18246 19684 18284
rect 18956 16606 18958 16658
rect 19010 16606 19012 16658
rect 18956 16594 19012 16606
rect 19068 17836 19572 17892
rect 18060 15708 18564 15764
rect 18956 16324 19012 16334
rect 18060 15538 18116 15708
rect 18060 15486 18062 15538
rect 18114 15486 18116 15538
rect 18060 15474 18116 15486
rect 17948 14466 18004 14476
rect 18284 14418 18340 15708
rect 18508 15316 18564 15326
rect 18508 15222 18564 15260
rect 18956 15148 19012 16268
rect 19068 16322 19124 17836
rect 19628 17780 19684 17790
rect 19628 17686 19684 17724
rect 19180 17668 19236 17678
rect 19180 17574 19236 17612
rect 19740 17668 19796 18620
rect 20076 18338 20132 18350
rect 20076 18286 20078 18338
rect 20130 18286 20132 18338
rect 20076 18228 20132 18286
rect 19964 17780 20020 17790
rect 20076 17780 20132 18172
rect 19740 17602 19796 17612
rect 19852 17778 20132 17780
rect 19852 17726 19966 17778
rect 20018 17726 20132 17778
rect 19852 17724 20132 17726
rect 20188 18226 20244 19292
rect 20412 19282 20468 19292
rect 20188 18174 20190 18226
rect 20242 18174 20244 18226
rect 20188 17780 20244 18174
rect 20860 19010 20916 19406
rect 20860 18958 20862 19010
rect 20914 18958 20916 19010
rect 19852 17556 19908 17724
rect 19964 17714 20020 17724
rect 20188 17714 20244 17724
rect 20524 17780 20580 17790
rect 20524 17686 20580 17724
rect 19852 17444 19908 17500
rect 19628 17388 19908 17444
rect 20188 17444 20244 17454
rect 19180 17108 19236 17118
rect 19628 17108 19684 17388
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19852 17108 19908 17118
rect 19628 17106 19908 17108
rect 19628 17054 19854 17106
rect 19906 17054 19908 17106
rect 19628 17052 19908 17054
rect 19180 17014 19236 17052
rect 19852 17042 19908 17052
rect 19068 16270 19070 16322
rect 19122 16270 19124 16322
rect 19068 16258 19124 16270
rect 19516 16658 19572 16670
rect 19516 16606 19518 16658
rect 19570 16606 19572 16658
rect 19516 16210 19572 16606
rect 19516 16158 19518 16210
rect 19570 16158 19572 16210
rect 19516 16146 19572 16158
rect 19628 16212 19684 16222
rect 19628 15540 19684 16156
rect 19852 16212 19908 16222
rect 19852 16118 19908 16156
rect 20188 15988 20244 17388
rect 20860 17220 20916 18958
rect 21084 18674 21140 18686
rect 21084 18622 21086 18674
rect 21138 18622 21140 18674
rect 20972 17780 21028 17790
rect 20972 17686 21028 17724
rect 20860 17154 20916 17164
rect 20972 17556 21028 17566
rect 20524 17108 20580 17118
rect 20524 17014 20580 17052
rect 20972 17106 21028 17500
rect 20972 17054 20974 17106
rect 21026 17054 21028 17106
rect 20972 17042 21028 17054
rect 21084 16996 21140 18622
rect 21308 18450 21364 18462
rect 21308 18398 21310 18450
rect 21362 18398 21364 18450
rect 21308 17332 21364 18398
rect 21308 17266 21364 17276
rect 21420 17220 21476 17230
rect 21420 17106 21476 17164
rect 21420 17054 21422 17106
rect 21474 17054 21476 17106
rect 21420 17042 21476 17054
rect 21084 16930 21140 16940
rect 20412 16324 20468 16334
rect 20412 16210 20468 16268
rect 20412 16158 20414 16210
rect 20466 16158 20468 16210
rect 20412 16146 20468 16158
rect 20860 16324 20916 16334
rect 20860 16210 20916 16268
rect 20860 16158 20862 16210
rect 20914 16158 20916 16210
rect 20860 16146 20916 16158
rect 20188 15922 20244 15932
rect 21420 15988 21476 15998
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19740 15540 19796 15550
rect 19628 15538 19796 15540
rect 19628 15486 19742 15538
rect 19794 15486 19796 15538
rect 19628 15484 19796 15486
rect 19292 15202 19348 15214
rect 19292 15150 19294 15202
rect 19346 15150 19348 15202
rect 19292 15148 19348 15150
rect 18956 15092 19124 15148
rect 19068 14754 19124 15092
rect 19068 14702 19070 14754
rect 19122 14702 19124 14754
rect 19068 14690 19124 14702
rect 19180 15092 19348 15148
rect 18284 14366 18286 14418
rect 18338 14366 18340 14418
rect 16044 14308 16100 14318
rect 15820 13636 15876 13646
rect 15372 13634 15876 13636
rect 15372 13582 15374 13634
rect 15426 13582 15822 13634
rect 15874 13582 15876 13634
rect 15372 13580 15876 13582
rect 15372 12962 15428 13580
rect 15820 13570 15876 13580
rect 15372 12910 15374 12962
rect 15426 12910 15428 12962
rect 15372 12740 15428 12910
rect 16044 12962 16100 14252
rect 16268 13748 16324 13758
rect 16268 13654 16324 13692
rect 16044 12910 16046 12962
rect 16098 12910 16100 12962
rect 16044 12898 16100 12910
rect 18284 13412 18340 14366
rect 15372 12674 15428 12684
rect 18284 12850 18340 13356
rect 19180 14308 19236 15092
rect 19404 14308 19460 14318
rect 19180 14306 19460 14308
rect 19180 14254 19406 14306
rect 19458 14254 19460 14306
rect 19180 14252 19460 14254
rect 19180 13634 19236 14252
rect 19404 14242 19460 14252
rect 19180 13582 19182 13634
rect 19234 13582 19236 13634
rect 19180 13412 19236 13582
rect 19068 13188 19124 13198
rect 19068 13094 19124 13132
rect 18284 12798 18286 12850
rect 18338 12798 18340 12850
rect 17052 12404 17108 12414
rect 15148 12238 15150 12290
rect 15202 12238 15204 12290
rect 14924 11172 14980 11182
rect 14140 10546 14196 10556
rect 14812 11170 14980 11172
rect 14812 11118 14926 11170
rect 14978 11118 14980 11170
rect 14812 11116 14980 11118
rect 14028 10434 14084 10444
rect 14028 9940 14084 9950
rect 13916 9938 14084 9940
rect 13916 9886 14030 9938
rect 14082 9886 14084 9938
rect 13916 9884 14084 9886
rect 13916 9604 13972 9884
rect 14028 9874 14084 9884
rect 13916 9538 13972 9548
rect 14812 9602 14868 11116
rect 14924 11106 14980 11116
rect 14812 9550 14814 9602
rect 14866 9550 14868 9602
rect 13804 7634 13860 7644
rect 14028 9266 14084 9278
rect 14028 9214 14030 9266
rect 14082 9214 14084 9266
rect 14028 8034 14084 9214
rect 14812 9044 14868 9550
rect 15036 9044 15092 9054
rect 14812 8988 15036 9044
rect 14028 7982 14030 8034
rect 14082 7982 14084 8034
rect 13692 7364 13748 7374
rect 14028 7364 14084 7982
rect 13692 7362 14084 7364
rect 13692 7310 13694 7362
rect 13746 7310 14084 7362
rect 13692 7308 14084 7310
rect 13692 7298 13748 7308
rect 13580 6750 13582 6802
rect 13634 6750 13636 6802
rect 13580 6738 13636 6750
rect 12460 6466 12852 6468
rect 12460 6414 12462 6466
rect 12514 6414 12852 6466
rect 12460 6412 12852 6414
rect 12460 6402 12516 6412
rect 12796 6132 12852 6412
rect 13020 6468 13076 6478
rect 13020 6466 13188 6468
rect 13020 6414 13022 6466
rect 13074 6414 13188 6466
rect 13020 6412 13188 6414
rect 13020 6402 13076 6412
rect 12796 6066 12852 6076
rect 13132 5460 13188 6412
rect 14028 6466 14084 7308
rect 15036 8258 15092 8988
rect 15148 8428 15204 12238
rect 16044 12292 16100 12302
rect 15484 11394 15540 11406
rect 15484 11342 15486 11394
rect 15538 11342 15540 11394
rect 15484 9826 15540 11342
rect 16044 11394 16100 12236
rect 16044 11342 16046 11394
rect 16098 11342 16100 11394
rect 16044 11330 16100 11342
rect 16492 11956 16548 11966
rect 16492 10834 16548 11900
rect 16492 10782 16494 10834
rect 16546 10782 16548 10834
rect 16492 10770 16548 10782
rect 17052 10834 17108 12348
rect 18284 11956 18340 12798
rect 18732 13076 18788 13086
rect 18732 12178 18788 13020
rect 18732 12126 18734 12178
rect 18786 12126 18788 12178
rect 18732 12114 18788 12126
rect 19180 12068 19236 13356
rect 19628 13076 19684 15484
rect 19740 15474 19796 15484
rect 21196 15316 21252 15326
rect 21196 15222 21252 15260
rect 21420 15314 21476 15932
rect 21420 15262 21422 15314
rect 21474 15262 21476 15314
rect 21420 15250 21476 15262
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19180 11936 19236 12012
rect 19292 12964 19348 12974
rect 19628 12944 19684 13020
rect 19740 13634 19796 13646
rect 19740 13582 19742 13634
rect 19794 13582 19796 13634
rect 19740 12964 19796 13582
rect 18284 11284 18340 11900
rect 17052 10782 17054 10834
rect 17106 10782 17108 10834
rect 17052 10770 17108 10782
rect 18060 11282 18340 11284
rect 18060 11230 18286 11282
rect 18338 11230 18340 11282
rect 18060 11228 18340 11230
rect 18060 10834 18116 11228
rect 18284 11218 18340 11228
rect 18508 11620 18564 11630
rect 18060 10782 18062 10834
rect 18114 10782 18116 10834
rect 18060 10770 18116 10782
rect 15484 9774 15486 9826
rect 15538 9774 15540 9826
rect 15484 9044 15540 9774
rect 15932 10724 15988 10734
rect 15932 9826 15988 10668
rect 17612 10612 17668 10622
rect 17612 10518 17668 10556
rect 18508 10500 18564 11564
rect 19068 11508 19124 11518
rect 19068 11414 19124 11452
rect 18508 10406 18564 10444
rect 15932 9774 15934 9826
rect 15986 9774 15988 9826
rect 15932 9762 15988 9774
rect 19292 9938 19348 12908
rect 19740 12898 19796 12908
rect 20188 13076 20244 13086
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 20188 12402 20244 13020
rect 20524 12964 20580 12974
rect 20524 12870 20580 12908
rect 20188 12350 20190 12402
rect 20242 12350 20244 12402
rect 20188 12338 20244 12350
rect 21420 12292 21476 12302
rect 21420 12198 21476 12236
rect 19628 12068 19684 12078
rect 21532 12068 21588 21868
rect 21644 20130 21700 21980
rect 21756 21700 21812 23886
rect 21868 23938 21924 24556
rect 22092 24050 22148 25678
rect 22092 23998 22094 24050
rect 22146 23998 22148 24050
rect 22092 23986 22148 23998
rect 21868 23886 21870 23938
rect 21922 23886 21924 23938
rect 21868 23874 21924 23886
rect 22204 23938 22260 27022
rect 22428 25730 22484 27916
rect 22652 27860 22708 28028
rect 22540 27804 22708 27860
rect 22764 27860 22820 27870
rect 22540 26404 22596 27804
rect 22764 26908 22820 27804
rect 22540 26338 22596 26348
rect 22652 26852 22820 26908
rect 22428 25678 22430 25730
rect 22482 25678 22484 25730
rect 22428 25666 22484 25678
rect 22204 23886 22206 23938
rect 22258 23886 22260 23938
rect 22204 23716 22260 23886
rect 22204 23650 22260 23660
rect 22316 25284 22372 25294
rect 22316 23492 22372 25228
rect 22540 23828 22596 23838
rect 22204 23436 22372 23492
rect 22428 23492 22484 23502
rect 21980 23268 22036 23278
rect 21980 22482 22036 23212
rect 21980 22430 21982 22482
rect 22034 22430 22036 22482
rect 21980 22372 22036 22430
rect 21980 22306 22036 22316
rect 21756 21634 21812 21644
rect 22204 21588 22260 23436
rect 22316 23268 22372 23278
rect 22316 23174 22372 23212
rect 21868 21586 22260 21588
rect 21868 21534 22206 21586
rect 22258 21534 22260 21586
rect 21868 21532 22260 21534
rect 21644 20078 21646 20130
rect 21698 20078 21700 20130
rect 21644 20066 21700 20078
rect 21756 21476 21812 21486
rect 21756 20802 21812 21420
rect 21756 20750 21758 20802
rect 21810 20750 21812 20802
rect 21756 20580 21812 20750
rect 21756 19684 21812 20524
rect 21644 19628 21812 19684
rect 21868 21026 21924 21532
rect 22204 21522 22260 21532
rect 22316 21474 22372 21486
rect 22316 21422 22318 21474
rect 22370 21422 22372 21474
rect 22204 21364 22260 21374
rect 22204 21270 22260 21308
rect 21868 20974 21870 21026
rect 21922 20974 21924 21026
rect 21644 18340 21700 19628
rect 21868 18564 21924 20974
rect 21980 21252 22036 21262
rect 21980 20692 22036 21196
rect 22316 21140 22372 21422
rect 21980 20626 22036 20636
rect 22092 21084 22372 21140
rect 22428 21140 22484 23436
rect 22540 22482 22596 23772
rect 22540 22430 22542 22482
rect 22594 22430 22596 22482
rect 22540 22418 22596 22430
rect 22092 20804 22148 21084
rect 22428 21074 22484 21084
rect 22540 21812 22596 21822
rect 22092 20356 22148 20748
rect 22092 20290 22148 20300
rect 22540 20188 22596 21756
rect 22652 21252 22708 26852
rect 22764 26404 22820 26414
rect 22764 26310 22820 26348
rect 22764 25844 22820 25854
rect 22764 21476 22820 25788
rect 22876 21812 22932 31612
rect 22988 30210 23044 30222
rect 22988 30158 22990 30210
rect 23042 30158 23044 30210
rect 22988 30100 23044 30158
rect 22988 30034 23044 30044
rect 22988 27300 23044 27310
rect 23100 27300 23156 31836
rect 23548 31890 23604 32396
rect 23548 31838 23550 31890
rect 23602 31838 23604 31890
rect 23548 31826 23604 31838
rect 23660 31780 23716 33854
rect 23884 34468 23940 34478
rect 23772 31780 23828 31790
rect 23660 31778 23828 31780
rect 23660 31726 23774 31778
rect 23826 31726 23828 31778
rect 23660 31724 23828 31726
rect 23772 31668 23828 31724
rect 23212 30882 23268 30894
rect 23212 30830 23214 30882
rect 23266 30830 23268 30882
rect 23212 30212 23268 30830
rect 23660 30882 23716 30894
rect 23660 30830 23662 30882
rect 23714 30830 23716 30882
rect 23660 30660 23716 30830
rect 23660 30594 23716 30604
rect 23212 28082 23268 30156
rect 23436 30100 23492 30110
rect 23436 29426 23492 30044
rect 23436 29374 23438 29426
rect 23490 29374 23492 29426
rect 23436 29362 23492 29374
rect 23548 29314 23604 29326
rect 23548 29262 23550 29314
rect 23602 29262 23604 29314
rect 23548 29204 23604 29262
rect 23548 28754 23604 29148
rect 23772 29204 23828 31612
rect 23772 29138 23828 29148
rect 23884 28980 23940 34412
rect 23996 34356 24052 34366
rect 24108 34356 24164 36990
rect 24220 36260 24276 40348
rect 24332 38388 24388 38398
rect 24332 37492 24388 38332
rect 24444 38050 24500 40572
rect 24444 37998 24446 38050
rect 24498 37998 24500 38050
rect 24444 37716 24500 37998
rect 24556 38722 24612 38734
rect 24556 38670 24558 38722
rect 24610 38670 24612 38722
rect 24556 37940 24612 38670
rect 24556 37874 24612 37884
rect 24444 37660 24612 37716
rect 24444 37492 24500 37502
rect 24332 37490 24500 37492
rect 24332 37438 24446 37490
rect 24498 37438 24500 37490
rect 24332 37436 24500 37438
rect 24332 37044 24388 37436
rect 24444 37426 24500 37436
rect 24332 36706 24388 36988
rect 24332 36654 24334 36706
rect 24386 36654 24388 36706
rect 24332 36642 24388 36654
rect 24444 36260 24500 36270
rect 24220 36204 24444 36260
rect 24444 36166 24500 36204
rect 24556 35140 24612 37660
rect 24332 35084 24612 35140
rect 23996 34354 24108 34356
rect 23996 34302 23998 34354
rect 24050 34302 24108 34354
rect 23996 34300 24108 34302
rect 23996 34290 24052 34300
rect 24108 34224 24164 34300
rect 24220 34914 24276 34926
rect 24220 34862 24222 34914
rect 24274 34862 24276 34914
rect 24220 34020 24276 34862
rect 23996 33684 24052 33694
rect 23996 31948 24052 33628
rect 24220 33346 24276 33964
rect 24332 34468 24388 35084
rect 24556 34914 24612 34926
rect 24556 34862 24558 34914
rect 24610 34862 24612 34914
rect 24332 33460 24388 34412
rect 24444 34804 24500 34814
rect 24444 34354 24500 34748
rect 24444 34302 24446 34354
rect 24498 34302 24500 34354
rect 24444 34132 24500 34302
rect 24444 34066 24500 34076
rect 24556 33906 24612 34862
rect 24556 33854 24558 33906
rect 24610 33854 24612 33906
rect 24556 33842 24612 33854
rect 24332 33404 24612 33460
rect 24220 33294 24222 33346
rect 24274 33294 24276 33346
rect 24220 33282 24276 33294
rect 24556 33346 24612 33404
rect 24556 33294 24558 33346
rect 24610 33294 24612 33346
rect 24556 33282 24612 33294
rect 24332 33236 24388 33246
rect 24332 32564 24388 33180
rect 24108 32452 24164 32462
rect 24332 32432 24388 32508
rect 24108 32358 24164 32396
rect 24556 32340 24612 32350
rect 24556 32246 24612 32284
rect 23996 31892 24164 31948
rect 23996 31780 24052 31790
rect 23996 31220 24052 31724
rect 23996 31088 24052 31164
rect 24108 28980 24164 31892
rect 24444 31892 24500 31902
rect 24444 31798 24500 31836
rect 24444 30884 24500 30894
rect 24444 30790 24500 30828
rect 24556 30548 24612 30558
rect 24444 30436 24500 30446
rect 24220 30100 24276 30110
rect 24276 30044 24388 30100
rect 24220 30006 24276 30044
rect 23548 28702 23550 28754
rect 23602 28702 23604 28754
rect 23548 28690 23604 28702
rect 23660 28924 23940 28980
rect 23996 28924 24164 28980
rect 23660 28642 23716 28924
rect 23660 28590 23662 28642
rect 23714 28590 23716 28642
rect 23660 28578 23716 28590
rect 23772 28532 23828 28924
rect 23772 28466 23828 28476
rect 23212 28030 23214 28082
rect 23266 28030 23268 28082
rect 23212 28018 23268 28030
rect 23660 28420 23716 28430
rect 23660 28082 23716 28364
rect 23660 28030 23662 28082
rect 23714 28030 23716 28082
rect 23660 28018 23716 28030
rect 22988 27298 23156 27300
rect 22988 27246 22990 27298
rect 23042 27246 23156 27298
rect 22988 27244 23156 27246
rect 22988 27234 23044 27244
rect 23996 27186 24052 28924
rect 24220 28532 24276 28542
rect 24108 28420 24164 28430
rect 24108 28082 24164 28364
rect 24108 28030 24110 28082
rect 24162 28030 24164 28082
rect 24108 28018 24164 28030
rect 23996 27134 23998 27186
rect 24050 27134 24052 27186
rect 23996 27076 24052 27134
rect 23996 27010 24052 27020
rect 24220 27074 24276 28476
rect 24220 27022 24222 27074
rect 24274 27022 24276 27074
rect 24220 27010 24276 27022
rect 24332 26908 24388 30044
rect 24220 26852 24388 26908
rect 23884 26628 23940 26638
rect 23884 26514 23940 26572
rect 23884 26462 23886 26514
rect 23938 26462 23940 26514
rect 23884 26450 23940 26462
rect 23660 26402 23716 26414
rect 23660 26350 23662 26402
rect 23714 26350 23716 26402
rect 23548 26292 23604 26302
rect 23548 26198 23604 26236
rect 22988 25956 23044 25966
rect 22988 25618 23044 25900
rect 23660 25732 23716 26350
rect 23660 25666 23716 25676
rect 22988 25566 22990 25618
rect 23042 25566 23044 25618
rect 22988 25554 23044 25566
rect 23548 25620 23604 25630
rect 23548 25526 23604 25564
rect 24108 25508 24164 25518
rect 23772 25506 24164 25508
rect 23772 25454 24110 25506
rect 24162 25454 24164 25506
rect 23772 25452 24164 25454
rect 23100 24722 23156 24734
rect 23100 24670 23102 24722
rect 23154 24670 23156 24722
rect 22988 23716 23044 23726
rect 22988 23622 23044 23660
rect 23100 23268 23156 24670
rect 23772 24722 23828 25452
rect 24108 25442 24164 25452
rect 23772 24670 23774 24722
rect 23826 24670 23828 24722
rect 23660 24052 23716 24062
rect 23772 24052 23828 24670
rect 23660 24050 23828 24052
rect 23660 23998 23662 24050
rect 23714 23998 23828 24050
rect 23660 23996 23828 23998
rect 23660 23986 23716 23996
rect 23772 23826 23828 23838
rect 23772 23774 23774 23826
rect 23826 23774 23828 23826
rect 23548 23714 23604 23726
rect 23548 23662 23550 23714
rect 23602 23662 23604 23714
rect 23548 23492 23604 23662
rect 22988 23212 23100 23268
rect 22988 22370 23044 23212
rect 23100 23202 23156 23212
rect 23436 23436 23604 23492
rect 23660 23604 23716 23614
rect 22988 22318 22990 22370
rect 23042 22318 23044 22370
rect 22988 22306 23044 22318
rect 23100 23044 23156 23054
rect 23436 23044 23492 23436
rect 23660 23380 23716 23548
rect 23100 23042 23492 23044
rect 23100 22990 23102 23042
rect 23154 22990 23492 23042
rect 23100 22988 23492 22990
rect 23548 23324 23716 23380
rect 22876 21746 22932 21756
rect 23100 21700 23156 22988
rect 23548 22482 23604 23324
rect 23660 23044 23716 23054
rect 23660 22950 23716 22988
rect 23548 22430 23550 22482
rect 23602 22430 23604 22482
rect 23548 22418 23604 22430
rect 23436 22148 23492 22158
rect 23548 22148 23604 22158
rect 23436 22146 23548 22148
rect 23436 22094 23438 22146
rect 23490 22094 23548 22146
rect 23436 22092 23548 22094
rect 23436 22082 23492 22092
rect 22764 21420 23044 21476
rect 22652 21186 22708 21196
rect 22092 20132 22596 20188
rect 22652 20690 22708 20702
rect 22652 20638 22654 20690
rect 22706 20638 22708 20690
rect 21644 18274 21700 18284
rect 21756 18508 21924 18564
rect 21980 20130 22148 20132
rect 21980 20078 22094 20130
rect 22146 20078 22148 20130
rect 21980 20076 22148 20078
rect 21756 17780 21812 18508
rect 21644 17724 21812 17780
rect 21644 17108 21700 17724
rect 21980 17668 22036 20076
rect 22092 20066 22148 20076
rect 22652 20020 22708 20638
rect 22988 20580 23044 21420
rect 22652 19954 22708 19964
rect 22876 20524 23044 20580
rect 22204 19796 22260 19806
rect 22204 19702 22260 19740
rect 22876 19460 22932 20524
rect 23100 20468 23156 21644
rect 23324 21924 23380 21934
rect 23212 21588 23268 21598
rect 23212 20692 23268 21532
rect 23324 21026 23380 21868
rect 23324 20974 23326 21026
rect 23378 20974 23380 21026
rect 23324 20962 23380 20974
rect 23548 21474 23604 22092
rect 23660 22146 23716 22158
rect 23660 22094 23662 22146
rect 23714 22094 23716 22146
rect 23660 21924 23716 22094
rect 23772 22148 23828 23774
rect 24220 23716 24276 26852
rect 24444 24834 24500 30380
rect 24556 29538 24612 30492
rect 24556 29486 24558 29538
rect 24610 29486 24612 29538
rect 24556 29474 24612 29486
rect 24668 29540 24724 41132
rect 24892 40514 24948 42588
rect 24892 40462 24894 40514
rect 24946 40462 24948 40514
rect 24892 40450 24948 40462
rect 25004 41300 25060 43374
rect 25116 43314 25172 43708
rect 25116 43262 25118 43314
rect 25170 43262 25172 43314
rect 25116 43250 25172 43262
rect 25116 42868 25172 42878
rect 25116 42774 25172 42812
rect 24780 40292 24836 40302
rect 24780 35812 24836 40236
rect 25004 39732 25060 41244
rect 25228 41860 25284 44604
rect 25676 44548 25732 44830
rect 25676 44482 25732 44492
rect 25788 44660 25844 44670
rect 25788 44434 25844 44604
rect 25788 44382 25790 44434
rect 25842 44382 25844 44434
rect 25788 44370 25844 44382
rect 25452 43428 25508 43438
rect 25228 41300 25284 41804
rect 25228 41234 25284 41244
rect 25340 42868 25396 42878
rect 25228 41076 25284 41086
rect 25228 40982 25284 41020
rect 25340 40852 25396 42812
rect 25228 40796 25396 40852
rect 24892 39676 25060 39732
rect 25116 39732 25172 39742
rect 24892 37490 24948 39676
rect 25116 39638 25172 39676
rect 25004 38722 25060 38734
rect 25004 38670 25006 38722
rect 25058 38670 25060 38722
rect 25004 38388 25060 38670
rect 25004 38322 25060 38332
rect 24892 37438 24894 37490
rect 24946 37438 24948 37490
rect 24892 37042 24948 37438
rect 24892 36990 24894 37042
rect 24946 36990 24948 37042
rect 24892 36978 24948 36990
rect 25004 36370 25060 36382
rect 25004 36318 25006 36370
rect 25058 36318 25060 36370
rect 25004 35924 25060 36318
rect 25004 35858 25060 35868
rect 25116 36258 25172 36270
rect 25116 36206 25118 36258
rect 25170 36206 25172 36258
rect 24780 35756 24948 35812
rect 24780 35586 24836 35598
rect 24780 35534 24782 35586
rect 24834 35534 24836 35586
rect 24780 34468 24836 35534
rect 24780 34402 24836 34412
rect 24892 34244 24948 35756
rect 24780 34188 24948 34244
rect 24780 30436 24836 34188
rect 24892 34020 24948 34030
rect 24892 30996 24948 33964
rect 25116 33012 25172 36206
rect 25228 36148 25284 40796
rect 25340 40404 25396 40414
rect 25340 36482 25396 40348
rect 25340 36430 25342 36482
rect 25394 36430 25396 36482
rect 25340 36418 25396 36430
rect 25452 39396 25508 43372
rect 25564 43316 25620 43326
rect 25564 40626 25620 43260
rect 25676 43092 25732 43102
rect 25676 42308 25732 43036
rect 25900 42866 25956 46844
rect 26012 46450 26068 46462
rect 26012 46398 26014 46450
rect 26066 46398 26068 46450
rect 26012 46004 26068 46398
rect 26012 45938 26068 45948
rect 26012 44884 26068 44894
rect 26012 44790 26068 44828
rect 26012 43876 26068 43886
rect 26012 43762 26068 43820
rect 26012 43710 26014 43762
rect 26066 43710 26068 43762
rect 26012 43698 26068 43710
rect 25900 42814 25902 42866
rect 25954 42814 25956 42866
rect 25900 42802 25956 42814
rect 26124 42754 26180 47068
rect 26236 47012 26292 50428
rect 26684 50036 26740 50046
rect 26796 50036 26852 51996
rect 26908 51986 26964 51996
rect 27132 52052 27188 52062
rect 27132 51958 27188 51996
rect 27244 50820 27300 52780
rect 27468 52770 27524 52780
rect 27692 52612 27748 55132
rect 27356 52556 27748 52612
rect 27916 52834 27972 57260
rect 28700 56978 28756 57372
rect 28700 56926 28702 56978
rect 28754 56926 28756 56978
rect 28700 56914 28756 56926
rect 29484 56980 29540 57822
rect 29820 58660 29876 58670
rect 29820 57874 29876 58604
rect 29932 58546 29988 58940
rect 29932 58494 29934 58546
rect 29986 58494 29988 58546
rect 29932 58482 29988 58494
rect 30044 58772 30100 59276
rect 30156 59238 30212 59276
rect 30716 59332 30772 59342
rect 30716 59238 30772 59276
rect 32620 59332 32676 59342
rect 32620 59330 32788 59332
rect 32620 59278 32622 59330
rect 32674 59278 32788 59330
rect 32620 59276 32788 59278
rect 32620 59266 32676 59276
rect 30828 59220 30884 59230
rect 30828 59126 30884 59164
rect 32508 59218 32564 59230
rect 32508 59166 32510 59218
rect 32562 59166 32564 59218
rect 31276 59106 31332 59118
rect 31276 59054 31278 59106
rect 31330 59054 31332 59106
rect 30716 58996 30772 59006
rect 30716 58902 30772 58940
rect 29820 57822 29822 57874
rect 29874 57822 29876 57874
rect 29820 57810 29876 57822
rect 29708 57762 29764 57774
rect 29708 57710 29710 57762
rect 29762 57710 29764 57762
rect 29708 57652 29764 57710
rect 30044 57764 30100 58716
rect 31276 58772 31332 59054
rect 31276 58706 31332 58716
rect 30156 58660 30212 58670
rect 30156 58566 30212 58604
rect 30604 58660 30660 58670
rect 30492 58436 30548 58446
rect 30492 58342 30548 58380
rect 30044 57652 30100 57708
rect 29708 57596 30100 57652
rect 30604 57650 30660 58604
rect 31500 58436 31556 58446
rect 31276 58434 31556 58436
rect 31276 58382 31502 58434
rect 31554 58382 31556 58434
rect 31276 58380 31556 58382
rect 30604 57598 30606 57650
rect 30658 57598 30660 57650
rect 29596 56980 29652 56990
rect 29484 56978 29652 56980
rect 29484 56926 29598 56978
rect 29650 56926 29652 56978
rect 29484 56924 29652 56926
rect 29596 56914 29652 56924
rect 28812 56868 28868 56878
rect 28812 56774 28868 56812
rect 28028 56756 28084 56766
rect 28028 55410 28084 56700
rect 28588 56756 28644 56766
rect 28588 56662 28644 56700
rect 29260 56532 29316 56542
rect 28028 55358 28030 55410
rect 28082 55358 28084 55410
rect 28028 55346 28084 55358
rect 28252 55970 28308 55982
rect 28252 55918 28254 55970
rect 28306 55918 28308 55970
rect 28140 54516 28196 54526
rect 28140 54422 28196 54460
rect 28252 53620 28308 55918
rect 28476 55636 28532 55646
rect 28476 55186 28532 55580
rect 28476 55134 28478 55186
rect 28530 55134 28532 55186
rect 28476 55076 28532 55134
rect 28476 55010 28532 55020
rect 28588 54516 28644 54526
rect 29036 54516 29092 54526
rect 28588 54514 28756 54516
rect 28588 54462 28590 54514
rect 28642 54462 28756 54514
rect 28588 54460 28756 54462
rect 28588 54450 28644 54460
rect 28700 53954 28756 54460
rect 29036 54422 29092 54460
rect 28700 53902 28702 53954
rect 28754 53902 28756 53954
rect 28700 53732 28756 53902
rect 28700 53666 28756 53676
rect 28252 53554 28308 53564
rect 28812 53620 28868 53630
rect 28812 53618 29204 53620
rect 28812 53566 28814 53618
rect 28866 53566 29204 53618
rect 28812 53564 29204 53566
rect 28812 53554 28868 53564
rect 27916 52782 27918 52834
rect 27970 52782 27972 52834
rect 27356 52050 27412 52556
rect 27916 52164 27972 52782
rect 27916 52098 27972 52108
rect 28028 53506 28084 53518
rect 28028 53454 28030 53506
rect 28082 53454 28084 53506
rect 28028 53396 28084 53454
rect 27356 51998 27358 52050
rect 27410 51998 27412 52050
rect 27356 51986 27412 51998
rect 27468 52050 27524 52062
rect 27468 51998 27470 52050
rect 27522 51998 27524 52050
rect 27244 50754 27300 50764
rect 27468 51266 27524 51998
rect 27468 51214 27470 51266
rect 27522 51214 27524 51266
rect 27020 50706 27076 50718
rect 27020 50654 27022 50706
rect 27074 50654 27076 50706
rect 26908 50596 26964 50606
rect 26908 50502 26964 50540
rect 26684 50034 26852 50036
rect 26684 49982 26686 50034
rect 26738 49982 26852 50034
rect 26684 49980 26852 49982
rect 26684 49970 26740 49980
rect 27020 49700 27076 50654
rect 27356 50708 27412 50718
rect 27468 50708 27524 51214
rect 27356 50706 27524 50708
rect 27356 50654 27358 50706
rect 27410 50654 27524 50706
rect 27356 50652 27524 50654
rect 27804 52052 27860 52062
rect 27804 51378 27860 51996
rect 27804 51326 27806 51378
rect 27858 51326 27860 51378
rect 27356 50642 27412 50652
rect 27244 50596 27300 50606
rect 27244 49810 27300 50540
rect 27244 49758 27246 49810
rect 27298 49758 27300 49810
rect 27244 49746 27300 49758
rect 27356 49812 27412 49822
rect 26908 49698 27076 49700
rect 26908 49646 27022 49698
rect 27074 49646 27076 49698
rect 26908 49644 27076 49646
rect 26908 49476 26964 49644
rect 27020 49634 27076 49644
rect 26908 49420 27300 49476
rect 26460 49364 26516 49374
rect 26348 49140 26404 49150
rect 26348 49046 26404 49084
rect 26236 46946 26292 46956
rect 26348 48916 26404 48926
rect 26460 48916 26516 49308
rect 26404 48860 26516 48916
rect 27020 49252 27076 49262
rect 26236 46676 26292 46686
rect 26236 46582 26292 46620
rect 26348 46452 26404 48860
rect 26796 48804 26852 48814
rect 26796 48710 26852 48748
rect 26684 48580 26740 48590
rect 26572 48356 26628 48366
rect 26572 48262 26628 48300
rect 26572 47682 26628 47694
rect 26572 47630 26574 47682
rect 26626 47630 26628 47682
rect 26572 47570 26628 47630
rect 26572 47518 26574 47570
rect 26626 47518 26628 47570
rect 26572 47506 26628 47518
rect 26236 46396 26404 46452
rect 26236 43092 26292 46396
rect 26348 46116 26404 46126
rect 26348 44660 26404 46060
rect 26348 44594 26404 44604
rect 26460 44324 26516 44334
rect 26460 44230 26516 44268
rect 26348 44212 26404 44222
rect 26348 44118 26404 44156
rect 26572 44100 26628 44110
rect 26684 44100 26740 48524
rect 26796 47682 26852 47694
rect 26796 47630 26798 47682
rect 26850 47630 26852 47682
rect 26796 46676 26852 47630
rect 26796 46620 26964 46676
rect 26908 46228 26964 46620
rect 26908 46162 26964 46172
rect 26908 46004 26964 46014
rect 26908 45910 26964 45948
rect 26796 45778 26852 45790
rect 26796 45726 26798 45778
rect 26850 45726 26852 45778
rect 26796 45220 26852 45726
rect 26796 45154 26852 45164
rect 26908 45780 26964 45790
rect 26908 45106 26964 45724
rect 26908 45054 26910 45106
rect 26962 45054 26964 45106
rect 26908 44772 26964 45054
rect 27020 45108 27076 49196
rect 27132 48804 27188 48814
rect 27132 47458 27188 48748
rect 27244 47570 27300 49420
rect 27356 48804 27412 49756
rect 27580 48804 27636 48814
rect 27356 48738 27412 48748
rect 27468 48802 27636 48804
rect 27468 48750 27582 48802
rect 27634 48750 27636 48802
rect 27468 48748 27636 48750
rect 27244 47518 27246 47570
rect 27298 47518 27300 47570
rect 27244 47506 27300 47518
rect 27356 48132 27412 48142
rect 27132 47406 27134 47458
rect 27186 47406 27188 47458
rect 27132 47394 27188 47406
rect 27356 47460 27412 48076
rect 27356 47366 27412 47404
rect 27468 46228 27524 48748
rect 27580 48738 27636 48748
rect 27804 48580 27860 51326
rect 27916 51938 27972 51950
rect 27916 51886 27918 51938
rect 27970 51886 27972 51938
rect 27916 51044 27972 51886
rect 28028 51380 28084 53340
rect 29036 53060 29092 53070
rect 29036 52966 29092 53004
rect 28588 52948 28644 52958
rect 28364 52834 28420 52846
rect 28364 52782 28366 52834
rect 28418 52782 28420 52834
rect 28364 52500 28420 52782
rect 28364 52434 28420 52444
rect 28252 52164 28308 52174
rect 28252 51490 28308 52108
rect 28252 51438 28254 51490
rect 28306 51438 28308 51490
rect 28252 51426 28308 51438
rect 28476 51938 28532 51950
rect 28476 51886 28478 51938
rect 28530 51886 28532 51938
rect 28028 51314 28084 51324
rect 27916 50988 28196 51044
rect 28028 50820 28084 50830
rect 27916 50706 27972 50718
rect 27916 50654 27918 50706
rect 27970 50654 27972 50706
rect 27916 50596 27972 50654
rect 27916 50530 27972 50540
rect 28028 50482 28084 50764
rect 28028 50430 28030 50482
rect 28082 50430 28084 50482
rect 28028 50418 28084 50430
rect 28028 50148 28084 50158
rect 27916 49812 27972 49822
rect 27916 49718 27972 49756
rect 27916 49140 27972 49150
rect 28028 49140 28084 50092
rect 27972 49084 28084 49140
rect 27916 49008 27972 49084
rect 27804 48524 27972 48580
rect 27916 48018 27972 48524
rect 27916 47966 27918 48018
rect 27970 47966 27972 48018
rect 27916 47954 27972 47966
rect 27580 47348 27636 47358
rect 27580 47254 27636 47292
rect 27916 47348 27972 47358
rect 27804 46564 27860 46574
rect 27804 46470 27860 46508
rect 27468 46162 27524 46172
rect 27132 45780 27188 45790
rect 27132 45778 27300 45780
rect 27132 45726 27134 45778
rect 27186 45726 27300 45778
rect 27132 45724 27300 45726
rect 27132 45714 27188 45724
rect 27020 45042 27076 45052
rect 27244 45218 27300 45724
rect 27356 45778 27412 45790
rect 27356 45726 27358 45778
rect 27410 45726 27412 45778
rect 27356 45332 27412 45726
rect 27356 45266 27412 45276
rect 27580 45220 27636 45230
rect 27244 45166 27246 45218
rect 27298 45166 27300 45218
rect 27020 44884 27076 44894
rect 27020 44882 27188 44884
rect 27020 44830 27022 44882
rect 27074 44830 27188 44882
rect 27020 44828 27188 44830
rect 27020 44818 27076 44828
rect 26572 44098 26740 44100
rect 26572 44046 26574 44098
rect 26626 44046 26740 44098
rect 26572 44044 26740 44046
rect 26796 44716 26964 44772
rect 26236 43026 26292 43036
rect 26460 43876 26516 43886
rect 26460 43762 26516 43820
rect 26460 43710 26462 43762
rect 26514 43710 26516 43762
rect 26124 42702 26126 42754
rect 26178 42702 26180 42754
rect 25900 42642 25956 42654
rect 25900 42590 25902 42642
rect 25954 42590 25956 42642
rect 25676 42242 25732 42252
rect 25788 42532 25844 42542
rect 25564 40574 25566 40626
rect 25618 40574 25620 40626
rect 25564 40292 25620 40574
rect 25564 40226 25620 40236
rect 25228 36082 25284 36092
rect 25340 34468 25396 34478
rect 25116 32956 25284 33012
rect 25116 32452 25172 32462
rect 25004 32340 25060 32350
rect 25004 32246 25060 32284
rect 25004 31892 25060 31902
rect 25116 31892 25172 32396
rect 25004 31890 25172 31892
rect 25004 31838 25006 31890
rect 25058 31838 25172 31890
rect 25004 31836 25172 31838
rect 25004 31218 25060 31836
rect 25004 31166 25006 31218
rect 25058 31166 25060 31218
rect 25004 31154 25060 31166
rect 25116 31668 25172 31678
rect 25004 30996 25060 31006
rect 24892 30940 25004 30996
rect 24780 30370 24836 30380
rect 24668 29484 24948 29540
rect 24892 29092 24948 29484
rect 25004 29316 25060 30940
rect 25116 30884 25172 31612
rect 25116 30818 25172 30828
rect 25228 30210 25284 32956
rect 25340 30548 25396 34412
rect 25452 32004 25508 39340
rect 25676 39732 25732 39742
rect 25788 39732 25844 42476
rect 25900 42308 25956 42590
rect 26124 42644 26180 42702
rect 26124 42578 26180 42588
rect 26348 42532 26404 42542
rect 25900 42242 25956 42252
rect 26236 42530 26404 42532
rect 26236 42478 26350 42530
rect 26402 42478 26404 42530
rect 26236 42476 26404 42478
rect 25900 41858 25956 41870
rect 25900 41806 25902 41858
rect 25954 41806 25956 41858
rect 25900 40852 25956 41806
rect 25900 40786 25956 40796
rect 26236 40404 26292 42476
rect 26348 42466 26404 42476
rect 26460 42532 26516 43710
rect 26460 42466 26516 42476
rect 26572 42308 26628 44044
rect 26796 43708 26852 44716
rect 27020 44322 27076 44334
rect 27020 44270 27022 44322
rect 27074 44270 27076 44322
rect 27020 43764 27076 44270
rect 27132 43876 27188 44828
rect 27244 44772 27300 45166
rect 27468 45218 27636 45220
rect 27468 45166 27582 45218
rect 27634 45166 27636 45218
rect 27468 45164 27636 45166
rect 27468 45108 27524 45164
rect 27580 45154 27636 45164
rect 27244 44706 27300 44716
rect 27356 45052 27524 45108
rect 27692 45106 27748 45118
rect 27692 45054 27694 45106
rect 27746 45054 27748 45106
rect 27132 43810 27188 43820
rect 26796 43652 26964 43708
rect 27020 43698 27076 43708
rect 26796 43428 26852 43438
rect 26796 43334 26852 43372
rect 26684 42868 26740 42878
rect 26684 42774 26740 42812
rect 26796 42756 26852 42766
rect 26908 42756 26964 43596
rect 27356 43540 27412 45052
rect 27580 44772 27636 44782
rect 27468 44324 27524 44334
rect 27468 44230 27524 44268
rect 27580 44098 27636 44716
rect 27692 44546 27748 45054
rect 27804 45108 27860 45118
rect 27804 45014 27860 45052
rect 27916 44660 27972 47292
rect 28028 46004 28084 49084
rect 28140 48356 28196 50988
rect 28252 50484 28308 50494
rect 28252 50390 28308 50428
rect 28364 49700 28420 49710
rect 28476 49700 28532 51886
rect 28364 49698 28532 49700
rect 28364 49646 28366 49698
rect 28418 49646 28532 49698
rect 28364 49644 28532 49646
rect 28364 49634 28420 49644
rect 28364 49252 28420 49262
rect 28364 49138 28420 49196
rect 28364 49086 28366 49138
rect 28418 49086 28420 49138
rect 28364 49074 28420 49086
rect 28364 48468 28420 48478
rect 28252 48356 28308 48366
rect 28140 48300 28252 48356
rect 28252 48242 28308 48300
rect 28252 48190 28254 48242
rect 28306 48190 28308 48242
rect 28140 48130 28196 48142
rect 28140 48078 28142 48130
rect 28194 48078 28196 48130
rect 28140 46676 28196 48078
rect 28140 46452 28196 46620
rect 28252 47124 28308 48190
rect 28364 47570 28420 48412
rect 28364 47518 28366 47570
rect 28418 47518 28420 47570
rect 28364 47236 28420 47518
rect 28364 47170 28420 47180
rect 28252 46674 28308 47068
rect 28252 46622 28254 46674
rect 28306 46622 28308 46674
rect 28252 46610 28308 46622
rect 28140 46386 28196 46396
rect 28476 46452 28532 49644
rect 28028 45938 28084 45948
rect 28252 46228 28308 46238
rect 28252 45780 28308 46172
rect 28028 45666 28084 45678
rect 28028 45614 28030 45666
rect 28082 45614 28084 45666
rect 28028 45332 28084 45614
rect 28028 45266 28084 45276
rect 28140 45668 28196 45678
rect 27692 44494 27694 44546
rect 27746 44494 27748 44546
rect 27692 44482 27748 44494
rect 27804 44604 27972 44660
rect 28028 45108 28084 45118
rect 28028 44772 28084 45052
rect 27580 44046 27582 44098
rect 27634 44046 27636 44098
rect 27580 44034 27636 44046
rect 27244 43428 27300 43438
rect 27244 43334 27300 43372
rect 26852 42700 26964 42756
rect 26796 42624 26852 42700
rect 26236 40338 26292 40348
rect 26348 42252 26628 42308
rect 26124 40290 26180 40302
rect 26124 40238 26126 40290
rect 26178 40238 26180 40290
rect 26124 40180 26180 40238
rect 26124 40114 26180 40124
rect 26348 39844 26404 42252
rect 26572 42082 26628 42094
rect 26572 42030 26574 42082
rect 26626 42030 26628 42082
rect 26460 41076 26516 41086
rect 26572 41076 26628 42030
rect 26684 41970 26740 41982
rect 26684 41918 26686 41970
rect 26738 41918 26740 41970
rect 26684 41748 26740 41918
rect 26740 41692 26852 41748
rect 26684 41682 26740 41692
rect 26516 41020 26740 41076
rect 26460 40944 26516 41020
rect 26572 40628 26628 40638
rect 26572 40402 26628 40572
rect 26572 40350 26574 40402
rect 26626 40350 26628 40402
rect 26572 40338 26628 40350
rect 26684 40404 26740 41020
rect 26796 41074 26852 41692
rect 26796 41022 26798 41074
rect 26850 41022 26852 41074
rect 26796 40628 26852 41022
rect 26796 40562 26852 40572
rect 27020 41412 27076 41422
rect 26908 40516 26964 40526
rect 26796 40404 26852 40414
rect 26684 40402 26852 40404
rect 26684 40350 26798 40402
rect 26850 40350 26852 40402
rect 26684 40348 26852 40350
rect 26796 40338 26852 40348
rect 26908 40180 26964 40460
rect 26348 39778 26404 39788
rect 26684 40124 26964 40180
rect 25676 39730 25844 39732
rect 25676 39678 25678 39730
rect 25730 39678 25844 39730
rect 25676 39676 25844 39678
rect 25676 38164 25732 39676
rect 26124 39508 26180 39518
rect 26124 39394 26180 39452
rect 26124 39342 26126 39394
rect 26178 39342 26180 39394
rect 25788 38948 25844 38958
rect 25788 38834 25844 38892
rect 26012 38836 26068 38846
rect 25788 38782 25790 38834
rect 25842 38782 25844 38834
rect 25788 38770 25844 38782
rect 25900 38834 26068 38836
rect 25900 38782 26014 38834
rect 26066 38782 26068 38834
rect 25900 38780 26068 38782
rect 25900 38724 25956 38780
rect 26012 38770 26068 38780
rect 26124 38668 26180 39342
rect 26348 38948 26404 38958
rect 25900 38612 26068 38668
rect 26124 38612 26292 38668
rect 25564 37938 25620 37950
rect 25564 37886 25566 37938
rect 25618 37886 25620 37938
rect 25564 35700 25620 37886
rect 25676 37492 25732 38108
rect 25900 37492 25956 37502
rect 25676 37490 25956 37492
rect 25676 37438 25902 37490
rect 25954 37438 25956 37490
rect 25676 37436 25956 37438
rect 25900 37426 25956 37436
rect 26012 36596 26068 38612
rect 25900 36540 26068 36596
rect 26124 37940 26180 37950
rect 26124 37156 26180 37884
rect 25900 36484 25956 36540
rect 25564 34018 25620 35644
rect 25676 36482 25956 36484
rect 25676 36430 25902 36482
rect 25954 36430 25956 36482
rect 25676 36428 25956 36430
rect 25676 35252 25732 36428
rect 25900 36418 25956 36428
rect 26124 36482 26180 37100
rect 26124 36430 26126 36482
rect 26178 36430 26180 36482
rect 26124 36418 26180 36430
rect 26012 36372 26068 36382
rect 26012 36278 26068 36316
rect 25900 36260 25956 36270
rect 26236 36260 26292 38612
rect 26348 38162 26404 38892
rect 26348 38110 26350 38162
rect 26402 38110 26404 38162
rect 26348 38098 26404 38110
rect 26572 38500 26628 38510
rect 26572 38050 26628 38444
rect 26572 37998 26574 38050
rect 26626 37998 26628 38050
rect 26572 37986 26628 37998
rect 26348 37268 26404 37278
rect 26348 37174 26404 37212
rect 26572 36484 26628 36494
rect 26572 36390 26628 36428
rect 26236 36204 26628 36260
rect 25788 36036 25844 36046
rect 25788 35700 25844 35980
rect 25788 35606 25844 35644
rect 25900 35698 25956 36204
rect 26124 36148 26180 36158
rect 26012 35924 26068 35934
rect 26012 35830 26068 35868
rect 26124 35922 26180 36092
rect 26124 35870 26126 35922
rect 26178 35870 26180 35922
rect 26124 35858 26180 35870
rect 25900 35646 25902 35698
rect 25954 35646 25956 35698
rect 25676 35186 25732 35196
rect 25564 33966 25566 34018
rect 25618 33966 25620 34018
rect 25564 33908 25620 33966
rect 25564 33842 25620 33852
rect 25676 35028 25732 35038
rect 25676 34802 25732 34972
rect 25676 34750 25678 34802
rect 25730 34750 25732 34802
rect 25676 33796 25732 34750
rect 25676 33730 25732 33740
rect 25900 33460 25956 35646
rect 26348 35698 26404 35710
rect 26348 35646 26350 35698
rect 26402 35646 26404 35698
rect 26348 35588 26404 35646
rect 26348 35522 26404 35532
rect 26460 35364 26516 35374
rect 26348 34692 26404 34702
rect 26236 34636 26348 34692
rect 26012 34356 26068 34366
rect 26012 34262 26068 34300
rect 25452 31938 25508 31948
rect 25564 33404 25956 33460
rect 25564 31780 25620 33404
rect 25788 33234 25844 33246
rect 25788 33182 25790 33234
rect 25842 33182 25844 33234
rect 25452 31724 25620 31780
rect 25676 32674 25732 32686
rect 25676 32622 25678 32674
rect 25730 32622 25732 32674
rect 25452 30660 25508 31724
rect 25564 31554 25620 31566
rect 25564 31502 25566 31554
rect 25618 31502 25620 31554
rect 25564 30996 25620 31502
rect 25676 31108 25732 32622
rect 25788 32004 25844 33182
rect 26236 32900 26292 34636
rect 26348 34598 26404 34636
rect 26460 34468 26516 35308
rect 26236 32834 26292 32844
rect 26348 34412 26516 34468
rect 26348 33122 26404 34412
rect 26460 34244 26516 34254
rect 26460 33908 26516 34188
rect 26460 33842 26516 33852
rect 26348 33070 26350 33122
rect 26402 33070 26404 33122
rect 26348 32676 26404 33070
rect 26572 32788 26628 36204
rect 26684 35924 26740 40124
rect 27020 39618 27076 41356
rect 27244 41186 27300 41198
rect 27244 41134 27246 41186
rect 27298 41134 27300 41186
rect 27132 40964 27188 40974
rect 27132 40870 27188 40908
rect 27244 40516 27300 41134
rect 27244 40450 27300 40460
rect 27132 40404 27188 40414
rect 27132 40310 27188 40348
rect 27244 40068 27300 40078
rect 27244 39732 27300 40012
rect 27356 39956 27412 43484
rect 27692 42978 27748 42990
rect 27692 42926 27694 42978
rect 27746 42926 27748 42978
rect 27468 42530 27524 42542
rect 27468 42478 27470 42530
rect 27522 42478 27524 42530
rect 27468 42196 27524 42478
rect 27468 42130 27524 42140
rect 27692 41858 27748 42926
rect 27692 41806 27694 41858
rect 27746 41806 27748 41858
rect 27692 41794 27748 41806
rect 27804 41188 27860 44604
rect 27916 44436 27972 44446
rect 27916 44342 27972 44380
rect 28028 43988 28084 44716
rect 28140 44546 28196 45612
rect 28140 44494 28142 44546
rect 28194 44494 28196 44546
rect 28140 44482 28196 44494
rect 28028 43762 28084 43932
rect 28252 43988 28308 45724
rect 28364 45668 28420 45678
rect 28476 45668 28532 46396
rect 28588 46228 28644 52892
rect 28924 52162 28980 52174
rect 28924 52110 28926 52162
rect 28978 52110 28980 52162
rect 28700 52052 28756 52062
rect 28700 51266 28756 51996
rect 28700 51214 28702 51266
rect 28754 51214 28756 51266
rect 28700 50484 28756 51214
rect 28700 50418 28756 50428
rect 28812 50482 28868 50494
rect 28812 50430 28814 50482
rect 28866 50430 28868 50482
rect 28812 49924 28868 50430
rect 28924 50372 28980 52110
rect 29148 51602 29204 53564
rect 29148 51550 29150 51602
rect 29202 51550 29204 51602
rect 29148 51538 29204 51550
rect 29260 50596 29316 56476
rect 29708 56308 29764 57596
rect 30604 57586 30660 57598
rect 30716 58212 30772 58222
rect 31164 58212 31220 58222
rect 30044 56866 30100 56878
rect 30044 56814 30046 56866
rect 30098 56814 30100 56866
rect 30044 56756 30100 56814
rect 30492 56868 30548 56878
rect 30492 56774 30548 56812
rect 30044 56690 30100 56700
rect 30156 56308 30212 56318
rect 29708 56306 30212 56308
rect 29708 56254 30158 56306
rect 30210 56254 30212 56306
rect 29708 56252 30212 56254
rect 30156 56242 30212 56252
rect 30716 56306 30772 58156
rect 31052 58210 31220 58212
rect 31052 58158 31166 58210
rect 31218 58158 31220 58210
rect 31052 58156 31220 58158
rect 31052 56866 31108 58156
rect 31164 58146 31220 58156
rect 31276 57762 31332 58380
rect 31500 58370 31556 58380
rect 32060 58434 32116 58446
rect 32060 58382 32062 58434
rect 32114 58382 32116 58434
rect 32060 58212 32116 58382
rect 32508 58436 32564 59166
rect 32732 58548 32788 59276
rect 32844 59220 32900 59258
rect 32844 59154 32900 59164
rect 33628 59108 33684 59724
rect 33740 59778 33796 59790
rect 33740 59726 33742 59778
rect 33794 59726 33796 59778
rect 33740 59668 33796 59726
rect 33740 59602 33796 59612
rect 34188 59442 34244 59948
rect 50428 60002 50484 60014
rect 50428 59950 50430 60002
rect 50482 59950 50484 60002
rect 43708 59890 43764 59902
rect 43708 59838 43710 59890
rect 43762 59838 43764 59890
rect 34748 59778 34804 59790
rect 34748 59726 34750 59778
rect 34802 59726 34804 59778
rect 34748 59444 34804 59726
rect 35532 59780 35588 59790
rect 35532 59686 35588 59724
rect 36316 59780 36372 59790
rect 34188 59390 34190 59442
rect 34242 59390 34244 59442
rect 33964 59220 34020 59230
rect 33964 59126 34020 59164
rect 33852 59108 33908 59118
rect 33628 59052 33852 59108
rect 32732 58482 32788 58492
rect 32844 58996 32900 59006
rect 32508 58370 32564 58380
rect 32284 58324 32340 58334
rect 32060 58146 32116 58156
rect 32172 58268 32284 58324
rect 31276 57710 31278 57762
rect 31330 57710 31332 57762
rect 31276 57698 31332 57710
rect 31164 57652 31220 57662
rect 31164 57558 31220 57596
rect 32060 57650 32116 57662
rect 32060 57598 32062 57650
rect 32114 57598 32116 57650
rect 31724 57540 31780 57550
rect 31052 56814 31054 56866
rect 31106 56814 31108 56866
rect 31052 56644 31108 56814
rect 31500 56980 31556 56990
rect 31500 56756 31556 56924
rect 31724 56866 31780 57484
rect 31724 56814 31726 56866
rect 31778 56814 31780 56866
rect 31724 56802 31780 56814
rect 31500 56662 31556 56700
rect 31052 56578 31108 56588
rect 31388 56642 31444 56654
rect 31388 56590 31390 56642
rect 31442 56590 31444 56642
rect 31388 56532 31444 56590
rect 31388 56466 31444 56476
rect 30716 56254 30718 56306
rect 30770 56254 30772 56306
rect 30716 56242 30772 56254
rect 31276 55972 31332 55982
rect 29932 55188 29988 55198
rect 29932 55186 30212 55188
rect 29932 55134 29934 55186
rect 29986 55134 30212 55186
rect 29932 55132 30212 55134
rect 29932 55122 29988 55132
rect 29820 55074 29876 55086
rect 29820 55022 29822 55074
rect 29874 55022 29876 55074
rect 29708 53844 29764 53854
rect 29708 53750 29764 53788
rect 29596 53732 29652 53742
rect 29596 53638 29652 53676
rect 29820 53730 29876 55022
rect 30156 54516 30212 55132
rect 30156 54422 30212 54460
rect 30940 54740 30996 54750
rect 29820 53678 29822 53730
rect 29874 53678 29876 53730
rect 29820 53666 29876 53678
rect 29932 54402 29988 54414
rect 29932 54350 29934 54402
rect 29986 54350 29988 54402
rect 29932 53732 29988 54350
rect 30828 54404 30884 54414
rect 30828 54310 30884 54348
rect 29932 53666 29988 53676
rect 30156 53730 30212 53742
rect 30156 53678 30158 53730
rect 30210 53678 30212 53730
rect 29708 52946 29764 52958
rect 29708 52894 29710 52946
rect 29762 52894 29764 52946
rect 29708 52164 29764 52894
rect 29708 52070 29764 52108
rect 30044 52946 30100 52958
rect 30044 52894 30046 52946
rect 30098 52894 30100 52946
rect 30044 51716 30100 52894
rect 30156 52834 30212 53678
rect 30604 53732 30660 53742
rect 30156 52782 30158 52834
rect 30210 52782 30212 52834
rect 30156 52770 30212 52782
rect 30268 53058 30324 53070
rect 30268 53006 30270 53058
rect 30322 53006 30324 53058
rect 30044 51650 30100 51660
rect 30156 52162 30212 52174
rect 30156 52110 30158 52162
rect 30210 52110 30212 52162
rect 30156 51604 30212 52110
rect 30156 51538 30212 51548
rect 29372 51490 29428 51502
rect 29372 51438 29374 51490
rect 29426 51438 29428 51490
rect 29372 50708 29428 51438
rect 29484 51380 29540 51390
rect 30268 51380 30324 53006
rect 30604 52274 30660 53676
rect 30604 52222 30606 52274
rect 30658 52222 30660 52274
rect 30604 52210 30660 52222
rect 30716 51716 30772 51726
rect 29484 51378 30212 51380
rect 29484 51326 29486 51378
rect 29538 51326 30212 51378
rect 29484 51324 30212 51326
rect 29484 51314 29540 51324
rect 29372 50652 29988 50708
rect 29260 50540 29428 50596
rect 28924 50306 28980 50316
rect 28700 49868 28868 49924
rect 28700 46564 28756 49868
rect 28812 49700 28868 49710
rect 29148 49700 29204 49710
rect 28812 49698 28980 49700
rect 28812 49646 28814 49698
rect 28866 49646 28980 49698
rect 28812 49644 28980 49646
rect 28812 49634 28868 49644
rect 28812 49140 28868 49150
rect 28812 49046 28868 49084
rect 28812 48132 28868 48142
rect 28812 47572 28868 48076
rect 28812 47440 28868 47516
rect 28924 46676 28980 49644
rect 28924 46610 28980 46620
rect 28700 46498 28756 46508
rect 28588 46162 28644 46172
rect 28364 45666 28532 45668
rect 28364 45614 28366 45666
rect 28418 45614 28532 45666
rect 28364 45612 28532 45614
rect 28364 45602 28420 45612
rect 28476 44884 28532 45612
rect 28588 45668 28644 45678
rect 28588 45106 28644 45612
rect 28924 45666 28980 45678
rect 28924 45614 28926 45666
rect 28978 45614 28980 45666
rect 28588 45054 28590 45106
rect 28642 45054 28644 45106
rect 28588 45042 28644 45054
rect 28812 45556 28868 45566
rect 28812 45106 28868 45500
rect 28812 45054 28814 45106
rect 28866 45054 28868 45106
rect 28812 45042 28868 45054
rect 28700 44884 28756 44894
rect 28476 44828 28644 44884
rect 28588 44546 28644 44828
rect 28588 44494 28590 44546
rect 28642 44494 28644 44546
rect 28588 44482 28644 44494
rect 28028 43710 28030 43762
rect 28082 43710 28084 43762
rect 28028 43698 28084 43710
rect 28140 43764 28196 43774
rect 28140 43670 28196 43708
rect 28252 43762 28308 43932
rect 28252 43710 28254 43762
rect 28306 43710 28308 43762
rect 27916 43540 27972 43550
rect 27916 43446 27972 43484
rect 28252 42978 28308 43710
rect 28476 43652 28532 43662
rect 28476 43558 28532 43596
rect 28252 42926 28254 42978
rect 28306 42926 28308 42978
rect 28252 42914 28308 42926
rect 27916 42868 27972 42878
rect 27916 42774 27972 42812
rect 28028 42532 28084 42542
rect 28028 41972 28084 42476
rect 27916 41412 27972 41422
rect 27916 41318 27972 41356
rect 28028 41410 28084 41916
rect 28364 42530 28420 42542
rect 28364 42478 28366 42530
rect 28418 42478 28420 42530
rect 28364 41970 28420 42478
rect 28364 41918 28366 41970
rect 28418 41918 28420 41970
rect 28364 41524 28420 41918
rect 28364 41458 28420 41468
rect 28476 42084 28532 42094
rect 28028 41358 28030 41410
rect 28082 41358 28084 41410
rect 28028 41346 28084 41358
rect 28252 41412 28308 41422
rect 28252 41318 28308 41356
rect 27804 41132 28084 41188
rect 27356 39890 27412 39900
rect 27580 40740 27636 40750
rect 27244 39730 27524 39732
rect 27244 39678 27246 39730
rect 27298 39678 27524 39730
rect 27244 39676 27524 39678
rect 27244 39666 27300 39676
rect 27020 39566 27022 39618
rect 27074 39566 27076 39618
rect 27020 37268 27076 39566
rect 27020 37202 27076 37212
rect 27132 39620 27188 39630
rect 26796 35924 26852 35934
rect 26684 35922 26852 35924
rect 26684 35870 26798 35922
rect 26850 35870 26852 35922
rect 26684 35868 26852 35870
rect 26796 35476 26852 35868
rect 26796 35410 26852 35420
rect 27020 35140 27076 35150
rect 27020 35026 27076 35084
rect 27020 34974 27022 35026
rect 27074 34974 27076 35026
rect 27020 34962 27076 34974
rect 27132 34132 27188 39564
rect 27468 38668 27524 39676
rect 27356 38612 27524 38668
rect 27580 38668 27636 40684
rect 27804 40740 27860 40750
rect 27804 40626 27860 40684
rect 27804 40574 27806 40626
rect 27858 40574 27860 40626
rect 27804 40562 27860 40574
rect 28028 40628 28084 41132
rect 27692 40516 27748 40526
rect 28028 40496 28084 40572
rect 28140 41076 28196 41086
rect 27692 40422 27748 40460
rect 28028 40404 28084 40414
rect 27692 40180 27748 40190
rect 27692 39620 27748 40124
rect 27692 39554 27748 39564
rect 27804 39172 27860 39182
rect 27804 38946 27860 39116
rect 27804 38894 27806 38946
rect 27858 38894 27860 38946
rect 27804 38882 27860 38894
rect 27580 38612 27748 38668
rect 27244 38276 27300 38286
rect 27244 38162 27300 38220
rect 27244 38110 27246 38162
rect 27298 38110 27300 38162
rect 27244 38098 27300 38110
rect 27356 37940 27412 38612
rect 27580 37940 27636 37950
rect 27244 37884 27412 37940
rect 27468 37884 27580 37940
rect 27244 35700 27300 37884
rect 27356 37604 27412 37614
rect 27356 37378 27412 37548
rect 27356 37326 27358 37378
rect 27410 37326 27412 37378
rect 27356 37044 27412 37326
rect 27468 37266 27524 37884
rect 27580 37874 27636 37884
rect 27468 37214 27470 37266
rect 27522 37214 27524 37266
rect 27468 37156 27524 37214
rect 27468 37090 27524 37100
rect 27580 37154 27636 37166
rect 27580 37102 27582 37154
rect 27634 37102 27636 37154
rect 27356 36978 27412 36988
rect 27468 35700 27524 35710
rect 27244 35698 27524 35700
rect 27244 35646 27470 35698
rect 27522 35646 27524 35698
rect 27244 35644 27524 35646
rect 27020 34076 27188 34132
rect 26796 33572 26852 33582
rect 26796 33458 26852 33516
rect 26796 33406 26798 33458
rect 26850 33406 26852 33458
rect 26796 33394 26852 33406
rect 26572 32722 26628 32732
rect 26908 33236 26964 33246
rect 26236 32620 26404 32676
rect 26012 32564 26068 32574
rect 26012 32470 26068 32508
rect 25900 32450 25956 32462
rect 25900 32398 25902 32450
rect 25954 32398 25956 32450
rect 25900 32228 25956 32398
rect 26236 32340 26292 32620
rect 26908 32562 26964 33180
rect 26908 32510 26910 32562
rect 26962 32510 26964 32562
rect 26908 32452 26964 32510
rect 26908 32386 26964 32396
rect 25900 32162 25956 32172
rect 26012 32284 26292 32340
rect 27020 32340 27076 34076
rect 27244 34020 27300 34030
rect 27132 33908 27188 33918
rect 27132 33814 27188 33852
rect 27244 33906 27300 33964
rect 27244 33854 27246 33906
rect 27298 33854 27300 33906
rect 27244 33348 27300 33854
rect 27356 33572 27412 35644
rect 27468 35634 27524 35644
rect 27580 35588 27636 37102
rect 27692 35700 27748 38612
rect 27804 37940 27860 37978
rect 27804 37874 27860 37884
rect 27916 37826 27972 37838
rect 27916 37774 27918 37826
rect 27970 37774 27972 37826
rect 27916 37604 27972 37774
rect 27916 37538 27972 37548
rect 27804 37268 27860 37278
rect 27804 37174 27860 37212
rect 28028 36708 28084 40348
rect 28140 38050 28196 41020
rect 28476 39730 28532 42028
rect 28700 40740 28756 44828
rect 28812 44546 28868 44558
rect 28812 44494 28814 44546
rect 28866 44494 28868 44546
rect 28812 44098 28868 44494
rect 28924 44212 28980 45614
rect 28924 44146 28980 44156
rect 29036 44994 29092 45006
rect 29036 44942 29038 44994
rect 29090 44942 29092 44994
rect 28812 44046 28814 44098
rect 28866 44046 28868 44098
rect 28812 42756 28868 44046
rect 29036 43764 29092 44942
rect 29036 43698 29092 43708
rect 28812 42662 28868 42700
rect 29036 41972 29092 41982
rect 29036 41878 29092 41916
rect 28924 41858 28980 41870
rect 28924 41806 28926 41858
rect 28978 41806 28980 41858
rect 28924 41412 28980 41806
rect 28924 41346 28980 41356
rect 28812 41300 28868 41310
rect 29148 41300 29204 49644
rect 29372 46450 29428 50540
rect 29596 50034 29652 50652
rect 29932 50594 29988 50652
rect 29932 50542 29934 50594
rect 29986 50542 29988 50594
rect 29932 50530 29988 50542
rect 30156 50706 30212 51324
rect 30268 51378 30660 51380
rect 30268 51326 30270 51378
rect 30322 51326 30660 51378
rect 30268 51324 30660 51326
rect 30268 51314 30324 51324
rect 30156 50654 30158 50706
rect 30210 50654 30212 50706
rect 29596 49982 29598 50034
rect 29650 49982 29652 50034
rect 29596 49970 29652 49982
rect 29708 50484 29764 50494
rect 29484 49922 29540 49934
rect 29484 49870 29486 49922
rect 29538 49870 29540 49922
rect 29484 47460 29540 49870
rect 29708 49812 29764 50428
rect 30156 50428 30212 50654
rect 30604 50706 30660 51324
rect 30604 50654 30606 50706
rect 30658 50654 30660 50706
rect 30604 50484 30660 50654
rect 30156 50372 30436 50428
rect 30604 50418 30660 50428
rect 30716 51266 30772 51660
rect 30716 51214 30718 51266
rect 30770 51214 30772 51266
rect 30380 50034 30436 50372
rect 30380 49982 30382 50034
rect 30434 49982 30436 50034
rect 30380 49970 30436 49982
rect 30492 50372 30548 50382
rect 30492 50034 30548 50316
rect 30492 49982 30494 50034
rect 30546 49982 30548 50034
rect 30492 49970 30548 49982
rect 30604 50036 30660 50046
rect 29708 49718 29764 49756
rect 30268 49810 30324 49822
rect 30268 49758 30270 49810
rect 30322 49758 30324 49810
rect 30268 49700 30324 49758
rect 30268 49634 30324 49644
rect 29484 47394 29540 47404
rect 29820 49252 29876 49262
rect 29708 47236 29764 47246
rect 29708 47142 29764 47180
rect 29372 46398 29374 46450
rect 29426 46398 29428 46450
rect 29372 46386 29428 46398
rect 29596 46002 29652 46014
rect 29596 45950 29598 46002
rect 29650 45950 29652 46002
rect 29596 45556 29652 45950
rect 29708 46004 29764 46014
rect 29708 45778 29764 45948
rect 29708 45726 29710 45778
rect 29762 45726 29764 45778
rect 29708 45714 29764 45726
rect 29596 45490 29652 45500
rect 29484 45332 29540 45342
rect 29484 45238 29540 45276
rect 29372 45220 29428 45230
rect 29372 45126 29428 45164
rect 29260 45108 29316 45118
rect 29260 45014 29316 45052
rect 29484 44212 29540 44222
rect 29484 44118 29540 44156
rect 29260 43426 29316 43438
rect 29260 43374 29262 43426
rect 29314 43374 29316 43426
rect 29260 42084 29316 43374
rect 29708 43426 29764 43438
rect 29708 43374 29710 43426
rect 29762 43374 29764 43426
rect 29708 43316 29764 43374
rect 29260 42018 29316 42028
rect 29484 43260 29764 43316
rect 29484 41860 29540 43260
rect 29484 41794 29540 41804
rect 29596 42082 29652 42094
rect 29596 42030 29598 42082
rect 29650 42030 29652 42082
rect 29148 41244 29540 41300
rect 28812 41206 28868 41244
rect 29372 40852 29428 40862
rect 28700 40684 29092 40740
rect 28476 39678 28478 39730
rect 28530 39678 28532 39730
rect 28476 39508 28532 39678
rect 28476 39442 28532 39452
rect 28588 40628 28644 40638
rect 28140 37998 28142 38050
rect 28194 37998 28196 38050
rect 28140 37986 28196 37998
rect 28588 39058 28644 40572
rect 29036 40626 29092 40684
rect 29036 40574 29038 40626
rect 29090 40574 29092 40626
rect 28700 40290 28756 40302
rect 28700 40238 28702 40290
rect 28754 40238 28756 40290
rect 28700 40178 28756 40238
rect 28700 40126 28702 40178
rect 28754 40126 28756 40178
rect 28700 40114 28756 40126
rect 28588 39006 28590 39058
rect 28642 39006 28644 39058
rect 27916 36652 28084 36708
rect 28364 36708 28420 36718
rect 27804 35700 27860 35710
rect 27692 35698 27860 35700
rect 27692 35646 27806 35698
rect 27858 35646 27860 35698
rect 27692 35644 27860 35646
rect 27580 35522 27636 35532
rect 27692 35476 27748 35486
rect 27468 35364 27524 35374
rect 27468 34914 27524 35308
rect 27468 34862 27470 34914
rect 27522 34862 27524 34914
rect 27468 34850 27524 34862
rect 27692 34468 27748 35420
rect 27804 34692 27860 35644
rect 27804 34626 27860 34636
rect 27692 34412 27860 34468
rect 27468 34132 27524 34142
rect 27468 33908 27524 34076
rect 27468 33906 27748 33908
rect 27468 33854 27470 33906
rect 27522 33854 27748 33906
rect 27468 33852 27748 33854
rect 27468 33842 27524 33852
rect 27356 33506 27412 33516
rect 27692 33458 27748 33852
rect 27692 33406 27694 33458
rect 27746 33406 27748 33458
rect 27580 33348 27636 33358
rect 27244 33346 27636 33348
rect 27244 33294 27582 33346
rect 27634 33294 27636 33346
rect 27244 33292 27636 33294
rect 27580 33282 27636 33292
rect 25788 31938 25844 31948
rect 25900 31780 25956 31818
rect 25900 31714 25956 31724
rect 25676 31042 25732 31052
rect 25900 31556 25956 31566
rect 25564 30930 25620 30940
rect 25900 30994 25956 31500
rect 25900 30942 25902 30994
rect 25954 30942 25956 30994
rect 25900 30930 25956 30942
rect 25676 30884 25732 30894
rect 25676 30790 25732 30828
rect 26012 30772 26068 32284
rect 27020 32274 27076 32284
rect 27580 32340 27636 32350
rect 27580 32246 27636 32284
rect 27692 31948 27748 33406
rect 26572 31890 26628 31902
rect 26572 31838 26574 31890
rect 26626 31838 26628 31890
rect 26124 31780 26180 31790
rect 26124 31220 26180 31724
rect 26572 31780 26628 31838
rect 26796 31892 27748 31948
rect 26572 31714 26628 31724
rect 26684 31778 26740 31790
rect 26684 31726 26686 31778
rect 26738 31726 26740 31778
rect 26684 31556 26740 31726
rect 26684 31490 26740 31500
rect 26124 30994 26180 31164
rect 26124 30942 26126 30994
rect 26178 30942 26180 30994
rect 26124 30930 26180 30942
rect 26236 31332 26292 31342
rect 26012 30716 26180 30772
rect 25900 30660 25956 30670
rect 25452 30604 25732 30660
rect 25340 30492 25620 30548
rect 25228 30158 25230 30210
rect 25282 30158 25284 30210
rect 25228 30146 25284 30158
rect 25340 30212 25396 30222
rect 25340 30118 25396 30156
rect 25116 30098 25172 30110
rect 25116 30046 25118 30098
rect 25170 30046 25172 30098
rect 25116 29988 25172 30046
rect 25116 29540 25172 29932
rect 25564 29652 25620 30492
rect 25676 30324 25732 30604
rect 25676 30258 25732 30268
rect 25900 30210 25956 30604
rect 26012 30324 26068 30334
rect 26012 30230 26068 30268
rect 25900 30158 25902 30210
rect 25954 30158 25956 30210
rect 25900 30146 25956 30158
rect 25676 30100 25732 30110
rect 25676 30098 25844 30100
rect 25676 30046 25678 30098
rect 25730 30046 25844 30098
rect 25676 30044 25844 30046
rect 25676 30034 25732 30044
rect 25676 29652 25732 29662
rect 25564 29596 25676 29652
rect 25676 29520 25732 29596
rect 25788 29650 25844 30044
rect 26124 29876 26180 30716
rect 26124 29810 26180 29820
rect 25788 29598 25790 29650
rect 25842 29598 25844 29650
rect 25788 29586 25844 29598
rect 25900 29652 25956 29662
rect 26236 29652 26292 31276
rect 25900 29558 25956 29596
rect 26012 29596 26292 29652
rect 26460 31108 26516 31118
rect 26460 29652 26516 31052
rect 26572 30772 26628 30782
rect 26572 30678 26628 30716
rect 26796 30210 26852 31892
rect 27804 31780 27860 34412
rect 27916 33460 27972 36652
rect 28364 36614 28420 36652
rect 28588 36596 28644 39006
rect 29036 38724 29092 40574
rect 28812 37826 28868 37838
rect 28812 37774 28814 37826
rect 28866 37774 28868 37826
rect 28588 36530 28644 36540
rect 28700 37492 28756 37502
rect 28028 36484 28084 36494
rect 28028 35026 28084 36428
rect 28476 36484 28532 36494
rect 28476 36390 28532 36428
rect 28252 35588 28308 35598
rect 28252 35138 28308 35532
rect 28700 35308 28756 37436
rect 28812 37268 28868 37774
rect 29036 37268 29092 38668
rect 29148 40178 29204 40190
rect 29148 40126 29150 40178
rect 29202 40126 29204 40178
rect 29148 38946 29204 40126
rect 29148 38894 29150 38946
rect 29202 38894 29204 38946
rect 29148 37380 29204 38894
rect 29148 37286 29204 37324
rect 29260 38164 29316 38174
rect 29260 37378 29316 38108
rect 29260 37326 29262 37378
rect 29314 37326 29316 37378
rect 29260 37314 29316 37326
rect 28812 37266 29092 37268
rect 28812 37214 29038 37266
rect 29090 37214 29092 37266
rect 28812 37212 29092 37214
rect 28812 36370 28868 36382
rect 28812 36318 28814 36370
rect 28866 36318 28868 36370
rect 28812 35588 28868 36318
rect 28812 35522 28868 35532
rect 28924 35700 28980 35710
rect 28924 35586 28980 35644
rect 28924 35534 28926 35586
rect 28978 35534 28980 35586
rect 28924 35522 28980 35534
rect 28700 35252 28868 35308
rect 28252 35086 28254 35138
rect 28306 35086 28308 35138
rect 28252 35074 28308 35086
rect 28028 34974 28030 35026
rect 28082 34974 28084 35026
rect 28028 34962 28084 34974
rect 28588 34692 28644 34702
rect 28588 34598 28644 34636
rect 28588 34132 28644 34142
rect 28476 34130 28644 34132
rect 28476 34078 28590 34130
rect 28642 34078 28644 34130
rect 28476 34076 28644 34078
rect 28028 34020 28084 34030
rect 28028 34018 28196 34020
rect 28028 33966 28030 34018
rect 28082 33966 28196 34018
rect 28028 33964 28196 33966
rect 28028 33954 28084 33964
rect 27916 33404 28084 33460
rect 27916 33234 27972 33246
rect 27916 33182 27918 33234
rect 27970 33182 27972 33234
rect 27916 32452 27972 33182
rect 27916 32358 27972 32396
rect 27916 31892 27972 31902
rect 28028 31892 28084 33404
rect 28140 32564 28196 33964
rect 28140 32432 28196 32508
rect 28476 33908 28532 34076
rect 28588 34066 28644 34076
rect 28476 33346 28532 33852
rect 28476 33294 28478 33346
rect 28530 33294 28532 33346
rect 28252 32228 28308 32238
rect 27916 31890 28084 31892
rect 27916 31838 27918 31890
rect 27970 31838 28084 31890
rect 27916 31836 28084 31838
rect 27916 31826 27972 31836
rect 27468 31724 27860 31780
rect 27356 31666 27412 31678
rect 27356 31614 27358 31666
rect 27410 31614 27412 31666
rect 27356 30996 27412 31614
rect 27356 30930 27412 30940
rect 26796 30158 26798 30210
rect 26850 30158 26852 30210
rect 26796 30146 26852 30158
rect 27132 30212 27188 30222
rect 26796 29876 26852 29886
rect 27132 29876 27188 30156
rect 27132 29820 27300 29876
rect 26460 29596 26628 29652
rect 25116 29474 25172 29484
rect 25004 29260 25172 29316
rect 24668 29036 24948 29092
rect 24556 28868 24612 28878
rect 24556 28754 24612 28812
rect 24556 28702 24558 28754
rect 24610 28702 24612 28754
rect 24556 28690 24612 28702
rect 24556 27860 24612 27870
rect 24556 27766 24612 27804
rect 24556 27524 24612 27534
rect 24556 26514 24612 27468
rect 24556 26462 24558 26514
rect 24610 26462 24612 26514
rect 24556 26450 24612 26462
rect 24668 25844 24724 29036
rect 25004 28308 25060 28318
rect 25004 28082 25060 28252
rect 25004 28030 25006 28082
rect 25058 28030 25060 28082
rect 25004 28018 25060 28030
rect 25004 27076 25060 27086
rect 24892 26962 24948 26974
rect 24892 26910 24894 26962
rect 24946 26910 24948 26962
rect 24892 26628 24948 26910
rect 24668 25778 24724 25788
rect 24780 26572 24948 26628
rect 24668 25508 24724 25518
rect 24668 25414 24724 25452
rect 24444 24782 24446 24834
rect 24498 24782 24500 24834
rect 24444 24770 24500 24782
rect 24668 24724 24724 24734
rect 24220 23650 24276 23660
rect 24444 23940 24500 23950
rect 23772 22082 23828 22092
rect 24108 22932 24164 22942
rect 23660 21858 23716 21868
rect 23548 21422 23550 21474
rect 23602 21422 23604 21474
rect 23212 20598 23268 20636
rect 23324 20580 23380 20590
rect 23324 20468 23380 20524
rect 23548 20468 23604 21422
rect 23100 20412 23380 20468
rect 23436 20412 23604 20468
rect 23660 20692 23716 20702
rect 22988 20356 23044 20366
rect 23044 20300 23268 20356
rect 22988 20290 23044 20300
rect 23100 19908 23156 19918
rect 23100 19814 23156 19852
rect 22092 19404 22932 19460
rect 22092 19122 22148 19404
rect 22316 19236 22372 19246
rect 22316 19142 22372 19180
rect 22092 19070 22094 19122
rect 22146 19070 22148 19122
rect 22092 19058 22148 19070
rect 22876 19124 22932 19404
rect 23100 19236 23156 19246
rect 22988 19124 23044 19134
rect 22876 19122 23044 19124
rect 22876 19070 22990 19122
rect 23042 19070 23044 19122
rect 22876 19068 23044 19070
rect 22204 19010 22260 19022
rect 22764 19012 22820 19022
rect 22204 18958 22206 19010
rect 22258 18958 22260 19010
rect 21644 17042 21700 17052
rect 21756 17612 22036 17668
rect 22092 17668 22148 17678
rect 22204 17668 22260 18958
rect 22092 17666 22260 17668
rect 22092 17614 22094 17666
rect 22146 17614 22260 17666
rect 22092 17612 22260 17614
rect 22540 19010 22820 19012
rect 22540 18958 22766 19010
rect 22818 18958 22820 19010
rect 22540 18956 22820 18958
rect 22540 17666 22596 18956
rect 22764 18946 22820 18956
rect 22540 17614 22542 17666
rect 22594 17614 22596 17666
rect 21644 16212 21700 16222
rect 21756 16212 21812 17612
rect 22092 17602 22148 17612
rect 22540 17602 22596 17614
rect 22652 18564 22708 18574
rect 22876 18564 22932 19068
rect 22988 19058 23044 19068
rect 22652 18562 22932 18564
rect 22652 18510 22654 18562
rect 22706 18510 22932 18562
rect 22652 18508 22932 18510
rect 21868 17442 21924 17454
rect 21868 17390 21870 17442
rect 21922 17390 21924 17442
rect 21868 17332 21924 17390
rect 21980 17444 22036 17454
rect 21980 17350 22036 17388
rect 21868 17266 21924 17276
rect 22316 17332 22372 17342
rect 21868 16994 21924 17006
rect 21868 16942 21870 16994
rect 21922 16942 21924 16994
rect 21868 16884 21924 16942
rect 22204 16996 22260 17006
rect 22204 16902 22260 16940
rect 21868 16818 21924 16828
rect 21644 16210 21756 16212
rect 21644 16158 21646 16210
rect 21698 16158 21756 16210
rect 21644 16156 21756 16158
rect 21644 16146 21700 16156
rect 21756 16080 21812 16156
rect 22316 16210 22372 17276
rect 22652 16324 22708 18508
rect 22876 18338 22932 18350
rect 22876 18286 22878 18338
rect 22930 18286 22932 18338
rect 22764 17668 22820 17678
rect 22876 17668 22932 18286
rect 22988 17892 23044 17902
rect 23100 17892 23156 19180
rect 23212 19124 23268 20300
rect 23436 19908 23492 20412
rect 23660 20356 23716 20636
rect 23548 20244 23604 20254
rect 23548 20130 23604 20188
rect 23660 20242 23716 20300
rect 23996 20690 24052 20702
rect 23996 20638 23998 20690
rect 24050 20638 24052 20690
rect 23660 20190 23662 20242
rect 23714 20190 23716 20242
rect 23660 20178 23716 20190
rect 23884 20244 23940 20254
rect 23996 20244 24052 20638
rect 23884 20242 24052 20244
rect 23884 20190 23886 20242
rect 23938 20190 24052 20242
rect 23884 20188 24052 20190
rect 23884 20178 23940 20188
rect 24108 20132 24164 22876
rect 24220 22370 24276 22382
rect 24220 22318 24222 22370
rect 24274 22318 24276 22370
rect 24220 22148 24276 22318
rect 24220 22082 24276 22092
rect 24444 21586 24500 23884
rect 24668 23604 24724 24668
rect 24780 23604 24836 26572
rect 24892 26404 24948 26414
rect 24892 26310 24948 26348
rect 24892 23604 24948 23614
rect 24780 23548 24892 23604
rect 24556 23268 24612 23278
rect 24556 21698 24612 23212
rect 24668 23266 24724 23548
rect 24892 23538 24948 23548
rect 24668 23214 24670 23266
rect 24722 23214 24724 23266
rect 24668 23202 24724 23214
rect 24780 23268 24836 23278
rect 24780 23174 24836 23212
rect 24892 23156 24948 23166
rect 24780 22932 24836 22942
rect 24892 22932 24948 23100
rect 24780 22930 24948 22932
rect 24780 22878 24782 22930
rect 24834 22878 24948 22930
rect 24780 22876 24948 22878
rect 24780 22866 24836 22876
rect 24780 22260 24836 22270
rect 24556 21646 24558 21698
rect 24610 21646 24612 21698
rect 24556 21634 24612 21646
rect 24668 22258 24836 22260
rect 24668 22206 24782 22258
rect 24834 22206 24836 22258
rect 24668 22204 24836 22206
rect 24668 21812 24724 22204
rect 24780 22194 24836 22204
rect 24444 21534 24446 21586
rect 24498 21534 24500 21586
rect 24332 20916 24388 20926
rect 24332 20822 24388 20860
rect 24220 20580 24276 20590
rect 24220 20486 24276 20524
rect 23548 20078 23550 20130
rect 23602 20078 23604 20130
rect 23548 20066 23604 20078
rect 23996 20076 24164 20132
rect 24444 20356 24500 21534
rect 24444 20242 24500 20300
rect 24444 20190 24446 20242
rect 24498 20190 24500 20242
rect 23436 19852 23716 19908
rect 23212 19058 23268 19068
rect 23548 18564 23604 18574
rect 23548 18470 23604 18508
rect 22988 17890 23156 17892
rect 22988 17838 22990 17890
rect 23042 17838 23156 17890
rect 22988 17836 23156 17838
rect 22988 17826 23044 17836
rect 23100 17668 23156 17678
rect 22876 17612 23100 17668
rect 22764 17108 22820 17612
rect 23100 17536 23156 17612
rect 23548 17220 23604 17230
rect 23660 17220 23716 19852
rect 23772 19796 23828 19806
rect 23772 19346 23828 19740
rect 23772 19294 23774 19346
rect 23826 19294 23828 19346
rect 23772 19282 23828 19294
rect 23772 19124 23828 19134
rect 23772 18340 23828 19068
rect 23884 18564 23940 18574
rect 23884 18470 23940 18508
rect 23772 18284 23940 18340
rect 23772 17890 23828 17902
rect 23772 17838 23774 17890
rect 23826 17838 23828 17890
rect 23772 17778 23828 17838
rect 23772 17726 23774 17778
rect 23826 17726 23828 17778
rect 23772 17714 23828 17726
rect 23884 17220 23940 18284
rect 23604 17164 23716 17220
rect 23772 17164 23940 17220
rect 22988 17108 23044 17118
rect 22764 17106 23044 17108
rect 22764 17054 22990 17106
rect 23042 17054 23044 17106
rect 22764 17052 23044 17054
rect 22988 16996 23044 17052
rect 22988 16930 23044 16940
rect 23212 17108 23268 17118
rect 22652 16258 22708 16268
rect 22316 16158 22318 16210
rect 22370 16158 22372 16210
rect 22316 16146 22372 16158
rect 23212 16210 23268 17052
rect 23548 17106 23604 17164
rect 23548 17054 23550 17106
rect 23602 17054 23604 17106
rect 23548 17042 23604 17054
rect 23212 16158 23214 16210
rect 23266 16158 23268 16210
rect 23212 16146 23268 16158
rect 23324 16212 23380 16222
rect 22428 16098 22484 16110
rect 22428 16046 22430 16098
rect 22482 16046 22484 16098
rect 22204 15988 22260 15998
rect 22204 15894 22260 15932
rect 22428 15540 22484 16046
rect 22204 15484 22484 15540
rect 22540 15988 22596 15998
rect 22204 15426 22260 15484
rect 22204 15374 22206 15426
rect 22258 15374 22260 15426
rect 22204 15316 22260 15374
rect 22204 15250 22260 15260
rect 21644 15202 21700 15214
rect 21644 15150 21646 15202
rect 21698 15150 21700 15202
rect 21644 15148 21700 15150
rect 21644 15092 21812 15148
rect 21756 14532 21812 15092
rect 21868 14532 21924 14542
rect 21756 14530 21924 14532
rect 21756 14478 21870 14530
rect 21922 14478 21924 14530
rect 21756 14476 21924 14478
rect 21868 14466 21924 14476
rect 21644 14308 21700 14318
rect 21644 14214 21700 14252
rect 22540 13970 22596 15932
rect 22764 15986 22820 15998
rect 22764 15934 22766 15986
rect 22818 15934 22820 15986
rect 22764 14642 22820 15934
rect 22764 14590 22766 14642
rect 22818 14590 22820 14642
rect 22764 14578 22820 14590
rect 22876 15316 22932 15326
rect 22764 14420 22820 14430
rect 22876 14420 22932 15260
rect 22764 14418 22932 14420
rect 22764 14366 22766 14418
rect 22818 14366 22932 14418
rect 22764 14364 22932 14366
rect 22988 15202 23044 15214
rect 22988 15150 22990 15202
rect 23042 15150 23044 15202
rect 22988 14420 23044 15150
rect 22764 14354 22820 14364
rect 22988 14326 23044 14364
rect 22540 13918 22542 13970
rect 22594 13918 22596 13970
rect 22540 13906 22596 13918
rect 22428 13748 22484 13758
rect 22316 13746 22484 13748
rect 22316 13694 22430 13746
rect 22482 13694 22484 13746
rect 22316 13692 22484 13694
rect 22316 12962 22372 13692
rect 22428 13682 22484 13692
rect 22652 13748 22708 13758
rect 22652 13746 22820 13748
rect 22652 13694 22654 13746
rect 22706 13694 22820 13746
rect 22652 13692 22820 13694
rect 22652 13682 22708 13692
rect 22316 12910 22318 12962
rect 22370 12910 22372 12962
rect 21756 12738 21812 12750
rect 21756 12686 21758 12738
rect 21810 12686 21812 12738
rect 21756 12290 21812 12686
rect 21756 12238 21758 12290
rect 21810 12238 21812 12290
rect 21756 12226 21812 12238
rect 21532 12012 21812 12068
rect 19628 11506 19684 12012
rect 19628 11454 19630 11506
rect 19682 11454 19684 11506
rect 19628 11442 19684 11454
rect 21644 11508 21700 11518
rect 21644 11414 21700 11452
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19628 10724 19684 10734
rect 19628 10630 19684 10668
rect 19964 10612 20020 10622
rect 19964 10518 20020 10556
rect 20524 10612 20580 10622
rect 20524 10518 20580 10556
rect 21196 10612 21252 10622
rect 21196 10518 21252 10556
rect 21420 10500 21476 10510
rect 21420 10406 21476 10444
rect 19292 9886 19294 9938
rect 19346 9886 19348 9938
rect 18956 9716 19012 9726
rect 18956 9622 19012 9660
rect 18396 9604 18452 9614
rect 18396 9510 18452 9548
rect 18732 9604 18788 9614
rect 15484 8978 15540 8988
rect 16492 9042 16548 9054
rect 16492 8990 16494 9042
rect 16546 8990 16548 9042
rect 16492 8708 16548 8990
rect 17052 9044 17108 9054
rect 17052 8950 17108 8988
rect 17612 9044 17668 9054
rect 16492 8642 16548 8652
rect 17612 8930 17668 8988
rect 17612 8878 17614 8930
rect 17666 8878 17668 8930
rect 17612 8484 17668 8878
rect 18060 8930 18116 8942
rect 18060 8878 18062 8930
rect 18114 8878 18116 8930
rect 15148 8372 15540 8428
rect 17612 8418 17668 8428
rect 17948 8596 18004 8606
rect 15036 8206 15038 8258
rect 15090 8206 15092 8258
rect 14028 6414 14030 6466
rect 14082 6414 14084 6466
rect 13244 6132 13300 6142
rect 13244 6038 13300 6076
rect 14028 6132 14084 6414
rect 14476 6692 14532 6702
rect 14476 6466 14532 6636
rect 14476 6414 14478 6466
rect 14530 6414 14532 6466
rect 14028 6066 14084 6076
rect 14364 6132 14420 6142
rect 14364 6038 14420 6076
rect 13804 5682 13860 5694
rect 13804 5630 13806 5682
rect 13858 5630 13860 5682
rect 13804 5572 13860 5630
rect 13804 5506 13860 5516
rect 14252 5684 14308 5694
rect 13132 5394 13188 5404
rect 13580 5236 13636 5246
rect 13580 5142 13636 5180
rect 14252 5234 14308 5628
rect 14252 5182 14254 5234
rect 14306 5182 14308 5234
rect 14252 5170 14308 5182
rect 13020 5012 13076 5022
rect 13020 4338 13076 4956
rect 13020 4286 13022 4338
rect 13074 4286 13076 4338
rect 13020 4274 13076 4286
rect 11228 4050 11284 4060
rect 10108 3614 10110 3666
rect 10162 3614 10164 3666
rect 10108 3602 10164 3614
rect 7644 3490 7700 3500
rect 12908 3444 12964 3454
rect 12908 800 12964 3388
rect 13692 3444 13748 3454
rect 13692 3350 13748 3388
rect 14476 3332 14532 6414
rect 15036 6690 15092 8206
rect 15036 6638 15038 6690
rect 15090 6638 15092 6690
rect 15036 6132 15092 6638
rect 15372 8258 15428 8270
rect 15372 8206 15374 8258
rect 15426 8206 15428 8258
rect 15372 6580 15428 8206
rect 15372 6514 15428 6524
rect 15148 6132 15204 6142
rect 15036 6130 15204 6132
rect 15036 6078 15150 6130
rect 15202 6078 15204 6130
rect 15036 6076 15204 6078
rect 14924 5236 14980 5246
rect 15036 5236 15092 6076
rect 15148 6066 15204 6076
rect 15484 5236 15540 8372
rect 15708 8036 15764 8046
rect 15708 6690 15764 7980
rect 15708 6638 15710 6690
rect 15762 6638 15764 6690
rect 15708 6626 15764 6638
rect 17948 8034 18004 8540
rect 17948 7982 17950 8034
rect 18002 7982 18004 8034
rect 17948 6466 18004 7982
rect 17948 6414 17950 6466
rect 18002 6414 18004 6466
rect 15708 5908 15764 5918
rect 15708 5814 15764 5852
rect 16156 5906 16212 5918
rect 16156 5854 16158 5906
rect 16210 5854 16212 5906
rect 14924 5234 15428 5236
rect 14924 5182 14926 5234
rect 14978 5182 15428 5234
rect 14924 5180 15428 5182
rect 14924 5170 14980 5180
rect 15036 4450 15092 5180
rect 15372 5124 15428 5180
rect 15484 5170 15540 5180
rect 16044 5348 16100 5358
rect 15372 4992 15428 5068
rect 16044 5122 16100 5292
rect 16044 5070 16046 5122
rect 16098 5070 16100 5122
rect 16044 5058 16100 5070
rect 15036 4398 15038 4450
rect 15090 4398 15092 4450
rect 15036 4386 15092 4398
rect 15036 3668 15092 3678
rect 16156 3668 16212 5854
rect 16716 5908 16772 5918
rect 16716 5814 16772 5852
rect 17612 5906 17668 5918
rect 17612 5854 17614 5906
rect 17666 5854 17668 5906
rect 16604 5684 16660 5694
rect 15036 3666 16212 3668
rect 15036 3614 15038 3666
rect 15090 3614 16212 3666
rect 15036 3612 16212 3614
rect 16380 5236 16436 5246
rect 16380 3666 16436 5180
rect 16604 5236 16660 5628
rect 16604 5170 16660 5180
rect 16380 3614 16382 3666
rect 16434 3614 16436 3666
rect 15036 3602 15092 3612
rect 16380 3602 16436 3614
rect 16828 5124 16884 5134
rect 16828 3666 16884 5068
rect 17612 5124 17668 5854
rect 17612 4338 17668 5068
rect 17612 4286 17614 4338
rect 17666 4286 17668 4338
rect 17612 4274 17668 4286
rect 17948 5908 18004 6414
rect 16828 3614 16830 3666
rect 16882 3614 16884 3666
rect 16828 3602 16884 3614
rect 17724 3556 17780 3566
rect 17724 3462 17780 3500
rect 17948 3556 18004 5852
rect 18060 6132 18116 8878
rect 18620 8930 18676 8942
rect 18620 8878 18622 8930
rect 18674 8878 18676 8930
rect 18620 8708 18676 8878
rect 18620 8642 18676 8652
rect 18732 8596 18788 9548
rect 18620 8260 18676 8270
rect 18620 8166 18676 8204
rect 18732 7698 18788 8540
rect 19292 9604 19348 9886
rect 19292 8428 19348 9548
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 21308 9268 21364 9278
rect 21308 9174 21364 9212
rect 21644 9042 21700 9054
rect 21644 8990 21646 9042
rect 21698 8990 21700 9042
rect 21644 8428 21700 8990
rect 18732 7646 18734 7698
rect 18786 7646 18788 7698
rect 18732 7634 18788 7646
rect 19068 8372 19124 8382
rect 19292 8372 19572 8428
rect 19068 7700 19124 8316
rect 19516 8034 19572 8372
rect 21084 8372 21700 8428
rect 19516 7982 19518 8034
rect 19570 7982 19572 8034
rect 19180 7700 19236 7710
rect 19068 7698 19236 7700
rect 19068 7646 19182 7698
rect 19234 7646 19236 7698
rect 19068 7644 19236 7646
rect 19516 7700 19572 7982
rect 20636 8148 20692 8158
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19516 7644 20132 7700
rect 19180 7634 19236 7644
rect 19628 7476 19684 7486
rect 19628 7362 19684 7420
rect 19628 7310 19630 7362
rect 19682 7310 19684 7362
rect 18732 6916 18788 6926
rect 18732 6822 18788 6860
rect 19628 6916 19684 7310
rect 19628 6850 19684 6860
rect 19628 6690 19684 6702
rect 19628 6638 19630 6690
rect 19682 6638 19684 6690
rect 18060 4900 18116 6076
rect 18060 4834 18116 4844
rect 18172 6468 18228 6478
rect 18172 4338 18228 6412
rect 19404 6468 19460 6478
rect 19404 6374 19460 6412
rect 18284 5908 18340 5918
rect 18284 5814 18340 5852
rect 19068 5124 19124 5134
rect 19068 5030 19124 5068
rect 18172 4286 18174 4338
rect 18226 4286 18228 4338
rect 18172 4274 18228 4286
rect 18284 4900 18340 4910
rect 18172 3668 18228 3678
rect 18284 3668 18340 4844
rect 19628 4564 19684 6638
rect 20076 6692 20132 7644
rect 20076 6636 20244 6692
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 20188 6132 20244 6636
rect 20636 6690 20692 8092
rect 20860 8034 20916 8046
rect 20860 7982 20862 8034
rect 20914 7982 20916 8034
rect 20860 7588 20916 7982
rect 20860 7494 20916 7532
rect 21084 7474 21140 8372
rect 21644 8036 21700 8046
rect 21644 7942 21700 7980
rect 21084 7422 21086 7474
rect 21138 7422 21140 7474
rect 21084 7410 21140 7422
rect 20636 6638 20638 6690
rect 20690 6638 20692 6690
rect 20636 6626 20692 6638
rect 21756 6692 21812 12012
rect 22316 11506 22372 12910
rect 22316 11454 22318 11506
rect 22370 11454 22372 11506
rect 22316 11442 22372 11454
rect 22652 12628 22708 12638
rect 22652 12402 22708 12572
rect 22652 12350 22654 12402
rect 22706 12350 22708 12402
rect 22652 11508 22708 12350
rect 22764 12402 22820 13692
rect 22764 12350 22766 12402
rect 22818 12350 22820 12402
rect 22764 12338 22820 12350
rect 23100 13746 23156 13758
rect 23100 13694 23102 13746
rect 23154 13694 23156 13746
rect 23100 12404 23156 13694
rect 23212 12852 23268 12862
rect 23212 12758 23268 12796
rect 23324 12628 23380 16156
rect 23660 16212 23716 16222
rect 23772 16212 23828 17164
rect 23996 17106 24052 20076
rect 24332 19122 24388 19134
rect 24332 19070 24334 19122
rect 24386 19070 24388 19122
rect 24332 18564 24388 19070
rect 24332 18498 24388 18508
rect 24332 18340 24388 18350
rect 24332 17668 24388 18284
rect 24444 17890 24500 20190
rect 24668 21586 24724 21756
rect 25004 21588 25060 27020
rect 25116 26852 25172 29260
rect 25900 29204 25956 29214
rect 25228 28980 25284 28990
rect 25228 28754 25284 28924
rect 25228 28702 25230 28754
rect 25282 28702 25284 28754
rect 25228 28690 25284 28702
rect 25788 28980 25844 28990
rect 25788 28754 25844 28924
rect 25788 28702 25790 28754
rect 25842 28702 25844 28754
rect 25788 28690 25844 28702
rect 25900 28196 25956 29148
rect 25788 28140 25956 28196
rect 25116 26786 25172 26796
rect 25452 27972 25508 27982
rect 25452 26404 25508 27916
rect 25676 27634 25732 27646
rect 25676 27582 25678 27634
rect 25730 27582 25732 27634
rect 25676 26908 25732 27582
rect 25788 27074 25844 28140
rect 25900 27972 25956 27982
rect 25900 27878 25956 27916
rect 26012 27746 26068 29596
rect 26124 29426 26180 29438
rect 26124 29374 26126 29426
rect 26178 29374 26180 29426
rect 26124 28644 26180 29374
rect 26460 29428 26516 29438
rect 26460 29334 26516 29372
rect 26124 28578 26180 28588
rect 26236 29204 26292 29214
rect 26236 28642 26292 29148
rect 26236 28590 26238 28642
rect 26290 28590 26292 28642
rect 26012 27694 26014 27746
rect 26066 27694 26068 27746
rect 26012 27682 26068 27694
rect 25788 27022 25790 27074
rect 25842 27022 25844 27074
rect 25788 27010 25844 27022
rect 26012 27186 26068 27198
rect 26236 27188 26292 28590
rect 26460 27748 26516 27758
rect 26012 27134 26014 27186
rect 26066 27134 26068 27186
rect 26012 27076 26068 27134
rect 26012 27010 26068 27020
rect 26124 27132 26292 27188
rect 26348 27746 26516 27748
rect 26348 27694 26462 27746
rect 26514 27694 26516 27746
rect 26348 27692 26516 27694
rect 26348 27300 26404 27692
rect 26460 27682 26516 27692
rect 25676 26852 25956 26908
rect 26124 26852 26180 27132
rect 26348 26908 26404 27244
rect 26572 27188 26628 29596
rect 26572 27122 26628 27132
rect 25676 26404 25732 26414
rect 25452 26402 25732 26404
rect 25452 26350 25678 26402
rect 25730 26350 25732 26402
rect 25452 26348 25732 26350
rect 25116 25508 25172 25518
rect 25116 23826 25172 25452
rect 25116 23774 25118 23826
rect 25170 23774 25172 23826
rect 25452 23940 25508 26348
rect 25676 26338 25732 26348
rect 25900 26066 25956 26852
rect 26012 26796 26180 26852
rect 26236 26852 26404 26908
rect 26460 26962 26516 26974
rect 26460 26910 26462 26962
rect 26514 26910 26516 26962
rect 26012 26516 26068 26796
rect 26236 26740 26292 26852
rect 26012 26450 26068 26460
rect 26124 26684 26292 26740
rect 25900 26014 25902 26066
rect 25954 26014 25956 26066
rect 25452 23808 25508 23884
rect 25788 25396 25844 25406
rect 25788 24610 25844 25340
rect 25788 24558 25790 24610
rect 25842 24558 25844 24610
rect 25116 21812 25172 23774
rect 25676 23716 25732 23726
rect 25676 22260 25732 23660
rect 25788 22482 25844 24558
rect 25900 24164 25956 26014
rect 26124 25618 26180 26684
rect 26236 26516 26292 26526
rect 26236 26422 26292 26460
rect 26460 25732 26516 26910
rect 26796 26516 26852 29820
rect 27132 29540 27188 29550
rect 27132 29446 27188 29484
rect 27244 29538 27300 29820
rect 27244 29486 27246 29538
rect 27298 29486 27300 29538
rect 27244 29474 27300 29486
rect 26908 29428 26964 29438
rect 26908 29334 26964 29372
rect 27468 29204 27524 31724
rect 28028 31444 28084 31836
rect 28028 31378 28084 31388
rect 28140 32002 28196 32014
rect 28140 31950 28142 32002
rect 28194 31950 28196 32002
rect 27580 30994 27636 31006
rect 27580 30942 27582 30994
rect 27634 30942 27636 30994
rect 27580 30772 27636 30942
rect 27580 30098 27636 30716
rect 27804 30996 27860 31006
rect 27804 30210 27860 30940
rect 27804 30158 27806 30210
rect 27858 30158 27860 30210
rect 27804 30146 27860 30158
rect 27580 30046 27582 30098
rect 27634 30046 27636 30098
rect 27580 30034 27636 30046
rect 26908 29148 27524 29204
rect 27580 29876 27636 29886
rect 26908 26516 26964 29148
rect 27132 28644 27188 28654
rect 27020 28532 27076 28542
rect 27020 28438 27076 28476
rect 27020 27972 27076 27982
rect 27020 27074 27076 27916
rect 27132 27186 27188 28588
rect 27580 27972 27636 29820
rect 28140 29426 28196 31950
rect 28140 29374 28142 29426
rect 28194 29374 28196 29426
rect 28028 29316 28084 29326
rect 28028 28866 28084 29260
rect 28028 28814 28030 28866
rect 28082 28814 28084 28866
rect 28028 28756 28084 28814
rect 28028 28690 28084 28700
rect 27580 27906 27636 27916
rect 27692 28642 27748 28654
rect 27692 28590 27694 28642
rect 27746 28590 27748 28642
rect 27692 28532 27748 28590
rect 27804 28644 27860 28654
rect 27804 28550 27860 28588
rect 27692 27858 27748 28476
rect 28140 28532 28196 29374
rect 28140 28466 28196 28476
rect 27692 27806 27694 27858
rect 27746 27806 27748 27858
rect 27692 27794 27748 27806
rect 28028 27860 28084 27870
rect 28028 27412 28084 27804
rect 28028 27346 28084 27356
rect 27132 27134 27134 27186
rect 27186 27134 27188 27186
rect 27132 27122 27188 27134
rect 28028 27188 28084 27198
rect 27020 27022 27022 27074
rect 27074 27022 27076 27074
rect 27020 27010 27076 27022
rect 28028 27076 28084 27132
rect 28140 27076 28196 27086
rect 28028 27074 28196 27076
rect 28028 27022 28142 27074
rect 28194 27022 28196 27074
rect 28028 27020 28196 27022
rect 27244 26964 27300 27002
rect 27244 26898 27300 26908
rect 27468 26850 27524 26862
rect 27468 26798 27470 26850
rect 27522 26798 27524 26850
rect 26908 26460 27300 26516
rect 26796 26450 26852 26460
rect 26908 26292 26964 26302
rect 26908 25844 26964 26236
rect 27132 26290 27188 26302
rect 27132 26238 27134 26290
rect 27186 26238 27188 26290
rect 27132 26068 27188 26238
rect 27244 26068 27300 26460
rect 27356 26292 27412 26302
rect 27356 26198 27412 26236
rect 27468 26178 27524 26798
rect 28028 26628 28084 27020
rect 28140 27010 28196 27020
rect 28252 26962 28308 32172
rect 28476 32002 28532 33294
rect 28700 32564 28756 32574
rect 28700 32470 28756 32508
rect 28476 31950 28478 32002
rect 28530 31950 28532 32002
rect 28476 31938 28532 31950
rect 28812 31780 28868 35252
rect 28700 31724 28868 31780
rect 28924 34356 28980 34366
rect 28364 31556 28420 31566
rect 28364 31462 28420 31500
rect 28476 30996 28532 31006
rect 28476 30902 28532 30940
rect 28364 30322 28420 30334
rect 28364 30270 28366 30322
rect 28418 30270 28420 30322
rect 28364 28084 28420 30270
rect 28476 29426 28532 29438
rect 28476 29374 28478 29426
rect 28530 29374 28532 29426
rect 28476 28644 28532 29374
rect 28588 29316 28644 29326
rect 28588 29222 28644 29260
rect 28476 28578 28532 28588
rect 28588 28532 28644 28542
rect 28588 28438 28644 28476
rect 28364 28018 28420 28028
rect 28252 26910 28254 26962
rect 28306 26910 28308 26962
rect 28252 26908 28308 26910
rect 27916 26572 28084 26628
rect 28140 26852 28308 26908
rect 28476 27972 28532 27982
rect 28476 26908 28532 27916
rect 28700 27860 28756 31724
rect 28812 31554 28868 31566
rect 28812 31502 28814 31554
rect 28866 31502 28868 31554
rect 28812 31220 28868 31502
rect 28812 31154 28868 31164
rect 28924 29988 28980 34300
rect 29036 34018 29092 37212
rect 29036 33966 29038 34018
rect 29090 33966 29092 34018
rect 29036 33236 29092 33966
rect 29036 33170 29092 33180
rect 29260 37156 29316 37166
rect 29260 33012 29316 37100
rect 29372 34132 29428 40796
rect 29484 37156 29540 41244
rect 29596 40628 29652 42030
rect 29820 40852 29876 49196
rect 30492 49138 30548 49150
rect 30492 49086 30494 49138
rect 30546 49086 30548 49138
rect 30044 48468 30100 48478
rect 30044 48242 30100 48412
rect 30492 48468 30548 49086
rect 30492 48402 30548 48412
rect 30604 48916 30660 49980
rect 30716 49250 30772 51214
rect 30940 50428 30996 54684
rect 31276 54740 31332 55916
rect 31836 55972 31892 55982
rect 31836 55878 31892 55916
rect 31388 55860 31444 55870
rect 31388 55468 31444 55804
rect 32060 55860 32116 57598
rect 32172 57652 32228 58268
rect 32284 58230 32340 58268
rect 32172 57586 32228 57596
rect 32396 58212 32452 58222
rect 32396 57650 32452 58156
rect 32396 57598 32398 57650
rect 32450 57598 32452 57650
rect 32396 57586 32452 57598
rect 32732 57652 32788 57662
rect 32844 57652 32900 58940
rect 32956 58548 33012 58558
rect 32956 58454 33012 58492
rect 33180 58436 33236 58446
rect 33180 58342 33236 58380
rect 33516 58436 33572 58446
rect 33516 58342 33572 58380
rect 33740 58436 33796 58446
rect 33628 58324 33684 58334
rect 33628 57762 33684 58268
rect 33740 57874 33796 58380
rect 33740 57822 33742 57874
rect 33794 57822 33796 57874
rect 33740 57810 33796 57822
rect 33852 57876 33908 59052
rect 34076 58996 34132 59006
rect 34076 58902 34132 58940
rect 33964 57876 34020 57886
rect 33852 57874 34020 57876
rect 33852 57822 33966 57874
rect 34018 57822 34020 57874
rect 33852 57820 34020 57822
rect 33964 57810 34020 57820
rect 33628 57710 33630 57762
rect 33682 57710 33684 57762
rect 33628 57698 33684 57710
rect 32732 57650 32900 57652
rect 32732 57598 32734 57650
rect 32786 57598 32900 57650
rect 32732 57596 32900 57598
rect 32732 57586 32788 57596
rect 32508 57540 32564 57550
rect 32508 57446 32564 57484
rect 34188 57092 34244 59390
rect 34412 59388 34804 59444
rect 34412 59332 34468 59388
rect 34300 59330 34468 59332
rect 34300 59278 34414 59330
rect 34466 59278 34468 59330
rect 34300 59276 34468 59278
rect 34300 57652 34356 59276
rect 34412 59266 34468 59276
rect 34524 59220 34580 59230
rect 35196 59220 35252 59230
rect 34412 58436 34468 58446
rect 34412 58342 34468 58380
rect 34524 57762 34580 59164
rect 34972 59218 35252 59220
rect 34972 59166 35198 59218
rect 35250 59166 35252 59218
rect 34972 59164 35252 59166
rect 34748 58996 34804 59006
rect 34748 58434 34804 58940
rect 34748 58382 34750 58434
rect 34802 58382 34804 58434
rect 34748 58370 34804 58382
rect 34972 58660 35028 59164
rect 35196 59154 35252 59164
rect 36316 59218 36372 59724
rect 36988 59780 37044 59790
rect 36988 59442 37044 59724
rect 36988 59390 36990 59442
rect 37042 59390 37044 59442
rect 36988 59378 37044 59390
rect 39676 59780 39732 59790
rect 36428 59332 36484 59342
rect 38220 59332 38276 59342
rect 36428 59330 36596 59332
rect 36428 59278 36430 59330
rect 36482 59278 36596 59330
rect 36428 59276 36596 59278
rect 36428 59266 36484 59276
rect 36316 59166 36318 59218
rect 36370 59166 36372 59218
rect 34972 58434 35028 58604
rect 34972 58382 34974 58434
rect 35026 58382 35028 58434
rect 34860 58212 34916 58222
rect 34860 58118 34916 58156
rect 34972 57764 35028 58382
rect 35084 58994 35140 59006
rect 35084 58942 35086 58994
rect 35138 58942 35140 58994
rect 35084 58436 35140 58942
rect 35420 58996 35476 59034
rect 35420 58930 35476 58940
rect 35532 58994 35588 59006
rect 35532 58942 35534 58994
rect 35586 58942 35588 58994
rect 35196 58828 35460 58838
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35196 58762 35460 58772
rect 35084 58370 35140 58380
rect 34524 57710 34526 57762
rect 34578 57710 34580 57762
rect 34524 57698 34580 57710
rect 34860 57708 35028 57764
rect 34300 57586 34356 57596
rect 34748 57652 34804 57662
rect 34748 57558 34804 57596
rect 34636 57092 34692 57102
rect 34188 57090 34692 57092
rect 34188 57038 34638 57090
rect 34690 57038 34692 57090
rect 34188 57036 34692 57038
rect 32284 56868 32340 56878
rect 32172 56756 32228 56766
rect 32172 56662 32228 56700
rect 32060 55794 32116 55804
rect 31388 55412 31556 55468
rect 31276 54674 31332 54684
rect 31164 52162 31220 52174
rect 31164 52110 31166 52162
rect 31218 52110 31220 52162
rect 31052 51268 31108 51278
rect 31052 51174 31108 51212
rect 30716 49198 30718 49250
rect 30770 49198 30772 49250
rect 30716 49186 30772 49198
rect 30828 50372 30996 50428
rect 30828 49140 30884 50372
rect 30940 49810 30996 49822
rect 30940 49758 30942 49810
rect 30994 49758 30996 49810
rect 30940 49700 30996 49758
rect 31164 49700 31220 52110
rect 31388 51716 31444 51726
rect 31276 51604 31332 51614
rect 31276 50818 31332 51548
rect 31276 50766 31278 50818
rect 31330 50766 31332 50818
rect 31276 50754 31332 50766
rect 31388 50594 31444 51660
rect 31388 50542 31390 50594
rect 31442 50542 31444 50594
rect 31388 50530 31444 50542
rect 31276 50484 31332 50494
rect 31276 50390 31332 50428
rect 30940 49644 31444 49700
rect 30828 49074 30884 49084
rect 30044 48190 30046 48242
rect 30098 48190 30100 48242
rect 30044 48178 30100 48190
rect 29932 48132 29988 48142
rect 29932 48038 29988 48076
rect 30156 48132 30212 48142
rect 29932 46676 29988 46686
rect 29932 46116 29988 46620
rect 30156 46674 30212 48076
rect 30156 46622 30158 46674
rect 30210 46622 30212 46674
rect 30156 46610 30212 46622
rect 30604 46674 30660 48860
rect 30716 49026 30772 49038
rect 30716 48974 30718 49026
rect 30770 48974 30772 49026
rect 30716 47236 30772 48974
rect 31052 48468 31108 48478
rect 30716 47170 30772 47180
rect 30828 48356 30884 48366
rect 30828 48242 30884 48300
rect 30828 48190 30830 48242
rect 30882 48190 30884 48242
rect 30604 46622 30606 46674
rect 30658 46622 30660 46674
rect 30604 46610 30660 46622
rect 30828 46674 30884 48190
rect 30828 46622 30830 46674
rect 30882 46622 30884 46674
rect 30828 46452 30884 46622
rect 30828 46386 30884 46396
rect 30940 46116 30996 46126
rect 29932 46050 29988 46060
rect 30716 46114 30996 46116
rect 30716 46062 30942 46114
rect 30994 46062 30996 46114
rect 30716 46060 30996 46062
rect 30268 46004 30324 46014
rect 29932 45780 29988 45790
rect 29932 45686 29988 45724
rect 30268 45330 30324 45948
rect 30716 45890 30772 46060
rect 30940 46050 30996 46060
rect 30716 45838 30718 45890
rect 30770 45838 30772 45890
rect 30716 45826 30772 45838
rect 30604 45780 30660 45790
rect 30492 45778 30660 45780
rect 30492 45726 30606 45778
rect 30658 45726 30660 45778
rect 30492 45724 30660 45726
rect 30380 45668 30436 45678
rect 30380 45574 30436 45612
rect 30268 45278 30270 45330
rect 30322 45278 30324 45330
rect 29932 45220 29988 45230
rect 29932 42978 29988 45164
rect 30044 45108 30100 45118
rect 30044 44546 30100 45052
rect 30044 44494 30046 44546
rect 30098 44494 30100 44546
rect 30044 44482 30100 44494
rect 30156 44996 30212 45006
rect 30156 44210 30212 44940
rect 30156 44158 30158 44210
rect 30210 44158 30212 44210
rect 30156 44146 30212 44158
rect 29932 42926 29934 42978
rect 29986 42926 29988 42978
rect 29932 42914 29988 42926
rect 30268 43762 30324 45278
rect 30492 45332 30548 45724
rect 30604 45714 30660 45724
rect 31052 45556 31108 48412
rect 30492 45200 30548 45276
rect 30604 45500 31108 45556
rect 31164 48242 31220 48254
rect 31164 48190 31166 48242
rect 31218 48190 31220 48242
rect 31164 48020 31220 48190
rect 31164 46002 31220 47964
rect 31276 47570 31332 47582
rect 31276 47518 31278 47570
rect 31330 47518 31332 47570
rect 31276 47012 31332 47518
rect 31276 46946 31332 46956
rect 31388 46788 31444 49644
rect 31164 45950 31166 46002
rect 31218 45950 31220 46002
rect 30604 45330 30660 45500
rect 30604 45278 30606 45330
rect 30658 45278 30660 45330
rect 30380 45106 30436 45118
rect 30380 45054 30382 45106
rect 30434 45054 30436 45106
rect 30380 44660 30436 45054
rect 30604 44884 30660 45278
rect 30940 45332 30996 45342
rect 30828 45220 30884 45230
rect 30940 45220 30996 45276
rect 30828 45218 30996 45220
rect 30828 45166 30830 45218
rect 30882 45166 30996 45218
rect 30828 45164 30996 45166
rect 30828 45154 30884 45164
rect 30604 44828 30772 44884
rect 30380 44604 30548 44660
rect 30268 43710 30270 43762
rect 30322 43710 30324 43762
rect 30044 42644 30100 42654
rect 30044 42642 30212 42644
rect 30044 42590 30046 42642
rect 30098 42590 30212 42642
rect 30044 42588 30212 42590
rect 30044 42578 30100 42588
rect 29820 40786 29876 40796
rect 29932 42530 29988 42542
rect 29932 42478 29934 42530
rect 29986 42478 29988 42530
rect 29932 41186 29988 42478
rect 29932 41134 29934 41186
rect 29986 41134 29988 41186
rect 29932 40628 29988 41134
rect 29596 40572 29988 40628
rect 30156 41300 30212 42588
rect 30156 41074 30212 41244
rect 30156 41022 30158 41074
rect 30210 41022 30212 41074
rect 29596 40514 29652 40572
rect 29596 40462 29598 40514
rect 29650 40462 29652 40514
rect 29596 40450 29652 40462
rect 29820 40404 29876 40414
rect 30156 40404 30212 41022
rect 29820 40402 30212 40404
rect 29820 40350 29822 40402
rect 29874 40350 30212 40402
rect 29820 40348 30212 40350
rect 30268 42196 30324 43710
rect 29820 40338 29876 40348
rect 30156 40180 30212 40190
rect 30268 40180 30324 42140
rect 30156 40178 30324 40180
rect 30156 40126 30158 40178
rect 30210 40126 30324 40178
rect 30156 40124 30324 40126
rect 30380 44436 30436 44446
rect 30156 40114 30212 40124
rect 29820 39956 29876 39966
rect 29820 39618 29876 39900
rect 29820 39566 29822 39618
rect 29874 39566 29876 39618
rect 29820 39554 29876 39566
rect 29708 38834 29764 38846
rect 29708 38782 29710 38834
rect 29762 38782 29764 38834
rect 29708 38164 29764 38782
rect 30044 38836 30100 38846
rect 29820 38724 29876 38762
rect 30044 38742 30100 38780
rect 29820 38658 29876 38668
rect 29708 38098 29764 38108
rect 29484 37090 29540 37100
rect 29596 37826 29652 37838
rect 30044 37828 30100 37838
rect 29596 37774 29598 37826
rect 29650 37774 29652 37826
rect 29484 36596 29540 36606
rect 29484 36482 29540 36540
rect 29484 36430 29486 36482
rect 29538 36430 29540 36482
rect 29484 36418 29540 36430
rect 29596 36372 29652 37774
rect 29932 37826 30100 37828
rect 29932 37774 30046 37826
rect 30098 37774 30100 37826
rect 29932 37772 30100 37774
rect 29708 37492 29764 37502
rect 29708 37398 29764 37436
rect 29484 35698 29540 35710
rect 29484 35646 29486 35698
rect 29538 35646 29540 35698
rect 29484 35476 29540 35646
rect 29484 35410 29540 35420
rect 29596 35364 29652 36316
rect 29596 35298 29652 35308
rect 29932 36482 29988 37772
rect 30044 37762 30100 37772
rect 30044 37380 30100 37390
rect 30044 36594 30100 37324
rect 30156 37156 30212 37166
rect 30156 37062 30212 37100
rect 30380 36708 30436 44380
rect 30492 43092 30548 44604
rect 30716 44436 30772 44828
rect 30716 44370 30772 44380
rect 30828 44098 30884 44110
rect 30828 44046 30830 44098
rect 30882 44046 30884 44098
rect 30828 43988 30884 44046
rect 30828 43922 30884 43932
rect 31052 43652 31108 43662
rect 31164 43652 31220 45950
rect 31276 46732 31444 46788
rect 31276 44884 31332 46732
rect 31500 45892 31556 55412
rect 32284 55410 32340 56812
rect 34636 56756 34692 57036
rect 34748 56980 34804 56990
rect 34860 56980 34916 57708
rect 35084 57650 35140 57662
rect 35084 57598 35086 57650
rect 35138 57598 35140 57650
rect 34972 57538 35028 57550
rect 34972 57486 34974 57538
rect 35026 57486 35028 57538
rect 34972 57092 35028 57486
rect 34972 57026 35028 57036
rect 34748 56978 34916 56980
rect 34748 56926 34750 56978
rect 34802 56926 34916 56978
rect 34748 56924 34916 56926
rect 34748 56914 34804 56924
rect 35084 56756 35140 57598
rect 35196 57260 35460 57270
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35196 57194 35460 57204
rect 35532 57092 35588 58942
rect 35644 58772 35700 58782
rect 35644 57874 35700 58716
rect 36092 58436 36148 58446
rect 36316 58436 36372 59166
rect 36092 58434 36372 58436
rect 36092 58382 36094 58434
rect 36146 58382 36372 58434
rect 36092 58380 36372 58382
rect 36428 58546 36484 58558
rect 36428 58494 36430 58546
rect 36482 58494 36484 58546
rect 36092 58100 36148 58380
rect 36092 58034 36148 58044
rect 35644 57822 35646 57874
rect 35698 57822 35700 57874
rect 35644 57652 35700 57822
rect 36428 57874 36484 58494
rect 36428 57822 36430 57874
rect 36482 57822 36484 57874
rect 36428 57810 36484 57822
rect 35644 57586 35700 57596
rect 35756 57764 35812 57774
rect 35644 57092 35700 57102
rect 35532 57090 35700 57092
rect 35532 57038 35646 57090
rect 35698 57038 35700 57090
rect 35532 57036 35700 57038
rect 35644 57026 35700 57036
rect 34636 56700 35140 56756
rect 32620 56642 32676 56654
rect 32620 56590 32622 56642
rect 32674 56590 32676 56642
rect 32620 55860 32676 56590
rect 35532 56308 35588 56318
rect 35532 56214 35588 56252
rect 35084 55972 35140 55982
rect 35084 55878 35140 55916
rect 32620 55794 32676 55804
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 35756 55468 35812 57708
rect 36316 57764 36372 57774
rect 36316 57670 36372 57708
rect 36540 57428 36596 59276
rect 38220 59238 38276 59276
rect 39340 59332 39396 59342
rect 36652 59218 36708 59230
rect 36652 59166 36654 59218
rect 36706 59166 36708 59218
rect 36652 58436 36708 59166
rect 38108 59218 38164 59230
rect 38108 59166 38110 59218
rect 38162 59166 38164 59218
rect 36764 59108 36820 59118
rect 36764 58546 36820 59052
rect 38108 59108 38164 59166
rect 38444 59220 38500 59230
rect 38444 59218 38612 59220
rect 38444 59166 38446 59218
rect 38498 59166 38612 59218
rect 38444 59164 38612 59166
rect 38444 59154 38500 59164
rect 38108 59042 38164 59052
rect 37660 58660 37716 58670
rect 37660 58566 37716 58604
rect 36764 58494 36766 58546
rect 36818 58494 36820 58546
rect 36764 58482 36820 58494
rect 36652 58370 36708 58380
rect 37548 58436 37604 58446
rect 38556 58436 38612 59164
rect 39340 59108 39396 59276
rect 39452 59108 39508 59118
rect 39340 59106 39508 59108
rect 39340 59054 39454 59106
rect 39506 59054 39508 59106
rect 39340 59052 39508 59054
rect 38892 58994 38948 59006
rect 38892 58942 38894 58994
rect 38946 58942 38948 58994
rect 38668 58436 38724 58446
rect 38556 58434 38724 58436
rect 38556 58382 38670 58434
rect 38722 58382 38724 58434
rect 38556 58380 38724 58382
rect 37548 58342 37604 58380
rect 38668 58370 38724 58380
rect 38892 58436 38948 58942
rect 39228 58996 39284 59006
rect 39228 58902 39284 58940
rect 38892 58370 38948 58380
rect 39116 58660 39172 58670
rect 39116 58434 39172 58604
rect 39116 58382 39118 58434
rect 39170 58382 39172 58434
rect 39116 58370 39172 58382
rect 37660 58324 37716 58334
rect 37660 58230 37716 58268
rect 38108 58212 38164 58222
rect 38108 57874 38164 58156
rect 38780 58212 38836 58222
rect 38780 58118 38836 58156
rect 38892 58210 38948 58222
rect 39340 58212 39396 59052
rect 39452 59042 39508 59052
rect 39452 58436 39508 58446
rect 39452 58342 39508 58380
rect 38892 58158 38894 58210
rect 38946 58158 38948 58210
rect 38108 57822 38110 57874
rect 38162 57822 38164 57874
rect 36988 57764 37044 57774
rect 36988 57670 37044 57708
rect 36540 57334 36596 57372
rect 37436 57538 37492 57550
rect 37436 57486 37438 57538
rect 37490 57486 37492 57538
rect 36540 57204 36596 57214
rect 35868 57092 35924 57102
rect 35868 56998 35924 57036
rect 36316 57092 36372 57102
rect 36092 56866 36148 56878
rect 36092 56814 36094 56866
rect 36146 56814 36148 56866
rect 32284 55358 32286 55410
rect 32338 55358 32340 55410
rect 32284 55346 32340 55358
rect 35532 55412 35812 55468
rect 35868 56308 35924 56318
rect 32172 55300 32228 55310
rect 32172 55206 32228 55244
rect 32844 55300 32900 55310
rect 32508 55188 32564 55198
rect 32508 55186 32676 55188
rect 32508 55134 32510 55186
rect 32562 55134 32676 55186
rect 32508 55132 32676 55134
rect 32508 55122 32564 55132
rect 32396 54514 32452 54526
rect 32396 54462 32398 54514
rect 32450 54462 32452 54514
rect 32284 54068 32340 54078
rect 32172 51938 32228 51950
rect 32172 51886 32174 51938
rect 32226 51886 32228 51938
rect 32060 51044 32116 51054
rect 31948 50988 32060 51044
rect 31948 50034 32004 50988
rect 32060 50978 32116 50988
rect 31948 49982 31950 50034
rect 32002 49982 32004 50034
rect 31948 49970 32004 49982
rect 32060 50818 32116 50830
rect 32060 50766 32062 50818
rect 32114 50766 32116 50818
rect 32060 50482 32116 50766
rect 32060 50430 32062 50482
rect 32114 50430 32116 50482
rect 31724 49924 31780 49934
rect 31724 49830 31780 49868
rect 31612 49810 31668 49822
rect 31612 49758 31614 49810
rect 31666 49758 31668 49810
rect 31612 48692 31668 49758
rect 31612 48626 31668 48636
rect 31724 47458 31780 47470
rect 31724 47406 31726 47458
rect 31778 47406 31780 47458
rect 31724 47236 31780 47406
rect 31724 47124 31780 47180
rect 31724 47068 32004 47124
rect 31612 47012 31668 47022
rect 31612 46004 31668 46956
rect 31612 45872 31668 45948
rect 31724 46114 31780 46126
rect 31724 46062 31726 46114
rect 31778 46062 31780 46114
rect 31500 45220 31556 45836
rect 31724 45330 31780 46062
rect 31724 45278 31726 45330
rect 31778 45278 31780 45330
rect 31724 45266 31780 45278
rect 31836 46004 31892 46014
rect 31612 45220 31668 45230
rect 31500 45218 31668 45220
rect 31500 45166 31614 45218
rect 31666 45166 31668 45218
rect 31500 45164 31668 45166
rect 31612 45154 31668 45164
rect 31388 45108 31444 45118
rect 31388 45014 31444 45052
rect 31276 44828 31668 44884
rect 31500 44322 31556 44334
rect 31500 44270 31502 44322
rect 31554 44270 31556 44322
rect 31052 43650 31220 43652
rect 31052 43598 31054 43650
rect 31106 43598 31220 43650
rect 31052 43596 31220 43598
rect 31052 43586 31108 43596
rect 31164 43540 31220 43596
rect 31164 43474 31220 43484
rect 31388 44100 31444 44110
rect 30492 43026 30548 43036
rect 31276 43316 31332 43326
rect 30492 42756 30548 42766
rect 30492 39618 30548 42700
rect 30828 42532 30884 42542
rect 31276 42532 31332 43260
rect 30716 42530 31332 42532
rect 30716 42478 30830 42530
rect 30882 42478 31332 42530
rect 30716 42476 31332 42478
rect 30716 41970 30772 42476
rect 30828 42466 30884 42476
rect 30828 42196 30884 42206
rect 30828 42082 30884 42140
rect 30828 42030 30830 42082
rect 30882 42030 30884 42082
rect 30828 42018 30884 42030
rect 31164 42084 31220 42094
rect 31164 41990 31220 42028
rect 30716 41918 30718 41970
rect 30770 41918 30772 41970
rect 30716 40628 30772 41918
rect 31052 41858 31108 41870
rect 31052 41806 31054 41858
rect 31106 41806 31108 41858
rect 30940 41636 30996 41646
rect 30940 41298 30996 41580
rect 30940 41246 30942 41298
rect 30994 41246 30996 41298
rect 30828 40628 30884 40638
rect 30716 40572 30828 40628
rect 30828 40534 30884 40572
rect 30492 39566 30494 39618
rect 30546 39566 30548 39618
rect 30492 36932 30548 39566
rect 30716 38836 30772 38846
rect 30716 38742 30772 38780
rect 30604 38724 30660 38734
rect 30604 38162 30660 38668
rect 30604 38110 30606 38162
rect 30658 38110 30660 38162
rect 30604 38098 30660 38110
rect 30716 38050 30772 38062
rect 30716 37998 30718 38050
rect 30770 37998 30772 38050
rect 30716 37492 30772 37998
rect 30716 37426 30772 37436
rect 30716 37156 30772 37166
rect 30940 37156 30996 41246
rect 31052 38668 31108 41806
rect 31388 40290 31444 44044
rect 31500 42756 31556 44270
rect 31500 42690 31556 42700
rect 31612 43314 31668 44828
rect 31836 44322 31892 45948
rect 31836 44270 31838 44322
rect 31890 44270 31892 44322
rect 31836 44258 31892 44270
rect 31948 43652 32004 47068
rect 32060 46116 32116 50430
rect 32172 50372 32228 51886
rect 32172 50306 32228 50316
rect 32060 46050 32116 46060
rect 32172 46564 32228 46574
rect 32172 45668 32228 46508
rect 32284 46452 32340 54012
rect 32396 53620 32452 54462
rect 32508 54404 32564 54414
rect 32508 53954 32564 54348
rect 32620 54292 32676 55132
rect 32620 54226 32676 54236
rect 32732 55186 32788 55198
rect 32732 55134 32734 55186
rect 32786 55134 32788 55186
rect 32508 53902 32510 53954
rect 32562 53902 32564 53954
rect 32508 53890 32564 53902
rect 32732 53842 32788 55134
rect 32844 54626 32900 55244
rect 33404 55300 33460 55310
rect 33404 55206 33460 55244
rect 33740 55298 33796 55310
rect 33740 55246 33742 55298
rect 33794 55246 33796 55298
rect 32844 54574 32846 54626
rect 32898 54574 32900 54626
rect 32844 54562 32900 54574
rect 33180 55076 33236 55086
rect 32732 53790 32734 53842
rect 32786 53790 32788 53842
rect 32732 53778 32788 53790
rect 32732 53620 32788 53630
rect 32396 53564 32732 53620
rect 32732 53488 32788 53564
rect 33068 52948 33124 52958
rect 33068 52274 33124 52892
rect 33068 52222 33070 52274
rect 33122 52222 33124 52274
rect 32396 51378 32452 51390
rect 32396 51326 32398 51378
rect 32450 51326 32452 51378
rect 32396 51044 32452 51326
rect 32620 51380 32676 51390
rect 32620 51286 32676 51324
rect 32732 51268 32788 51278
rect 32732 51174 32788 51212
rect 32396 50978 32452 50988
rect 32508 50818 32564 50830
rect 32508 50766 32510 50818
rect 32562 50766 32564 50818
rect 32508 50706 32564 50766
rect 32508 50654 32510 50706
rect 32562 50654 32564 50706
rect 32508 50642 32564 50654
rect 33068 50484 33124 52222
rect 33068 50390 33124 50428
rect 33180 50428 33236 55020
rect 33740 54404 33796 55246
rect 34300 55300 34356 55310
rect 34300 55206 34356 55244
rect 35420 55300 35476 55310
rect 35420 54738 35476 55244
rect 35420 54686 35422 54738
rect 35474 54686 35476 54738
rect 35420 54674 35476 54686
rect 35532 54738 35588 55412
rect 35644 55300 35700 55310
rect 35644 55206 35700 55244
rect 35532 54686 35534 54738
rect 35586 54686 35588 54738
rect 35532 54674 35588 54686
rect 35756 54516 35812 54526
rect 35644 54514 35812 54516
rect 35644 54462 35758 54514
rect 35810 54462 35812 54514
rect 35644 54460 35812 54462
rect 33740 54402 33908 54404
rect 33740 54350 33742 54402
rect 33794 54350 33908 54402
rect 33740 54348 33908 54350
rect 33740 54338 33796 54348
rect 33628 54292 33684 54302
rect 33628 54198 33684 54236
rect 33404 53620 33460 53630
rect 33404 53526 33460 53564
rect 33516 53618 33572 53630
rect 33516 53566 33518 53618
rect 33570 53566 33572 53618
rect 33516 52388 33572 53566
rect 33852 53172 33908 54348
rect 35644 54402 35700 54460
rect 35756 54450 35812 54460
rect 35644 54350 35646 54402
rect 35698 54350 35700 54402
rect 35644 54338 35700 54350
rect 34076 54292 34132 54302
rect 33964 53172 34020 53182
rect 33852 53170 34020 53172
rect 33852 53118 33966 53170
rect 34018 53118 34020 53170
rect 33852 53116 34020 53118
rect 33964 53106 34020 53116
rect 33740 53058 33796 53070
rect 33740 53006 33742 53058
rect 33794 53006 33796 53058
rect 33628 52948 33684 52958
rect 33628 52854 33684 52892
rect 33516 52332 33684 52388
rect 33292 52052 33348 52062
rect 33292 50596 33348 51996
rect 33628 51604 33684 52332
rect 33740 52052 33796 53006
rect 33740 51986 33796 51996
rect 33852 51604 33908 51614
rect 33628 51602 33908 51604
rect 33628 51550 33854 51602
rect 33906 51550 33908 51602
rect 33628 51548 33908 51550
rect 33852 51538 33908 51548
rect 33740 51378 33796 51390
rect 33740 51326 33742 51378
rect 33794 51326 33796 51378
rect 33740 51044 33796 51326
rect 33964 51380 34020 51390
rect 33964 51286 34020 51324
rect 34076 51378 34132 54236
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 35420 53732 35476 53742
rect 35756 53732 35812 53742
rect 35420 53730 35812 53732
rect 35420 53678 35422 53730
rect 35474 53678 35758 53730
rect 35810 53678 35812 53730
rect 35420 53676 35812 53678
rect 35420 53666 35476 53676
rect 35756 53666 35812 53676
rect 35084 53620 35140 53630
rect 35084 52274 35140 53564
rect 35196 53508 35252 53518
rect 35196 53414 35252 53452
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 35084 52222 35086 52274
rect 35138 52222 35140 52274
rect 35084 52210 35140 52222
rect 34076 51326 34078 51378
rect 34130 51326 34132 51378
rect 34076 51314 34132 51326
rect 34636 52162 34692 52174
rect 34636 52110 34638 52162
rect 34690 52110 34692 52162
rect 34636 51268 34692 52110
rect 34636 51174 34692 51212
rect 33740 50978 33796 50988
rect 34412 51154 34468 51166
rect 34412 51102 34414 51154
rect 34466 51102 34468 51154
rect 33404 50820 33460 50830
rect 33404 50726 33460 50764
rect 34412 50820 34468 51102
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 34412 50754 34468 50764
rect 34076 50708 34132 50718
rect 33404 50596 33460 50606
rect 33292 50594 33460 50596
rect 33292 50542 33406 50594
rect 33458 50542 33460 50594
rect 33292 50540 33460 50542
rect 33404 50484 33460 50540
rect 33404 50428 33684 50484
rect 32620 50372 32676 50382
rect 33180 50372 33348 50428
rect 32620 50034 32676 50316
rect 32620 49982 32622 50034
rect 32674 49982 32676 50034
rect 32620 49970 32676 49982
rect 32396 49812 32452 49822
rect 32396 49718 32452 49756
rect 32284 46386 32340 46396
rect 32508 49700 32564 49710
rect 32508 46116 32564 49644
rect 32732 49586 32788 49598
rect 32732 49534 32734 49586
rect 32786 49534 32788 49586
rect 32620 49140 32676 49150
rect 32620 49026 32676 49084
rect 32620 48974 32622 49026
rect 32674 48974 32676 49026
rect 32620 47012 32676 48974
rect 32732 48244 32788 49534
rect 32732 48178 32788 48188
rect 32956 49026 33012 49038
rect 32956 48974 32958 49026
rect 33010 48974 33012 49026
rect 32956 48132 33012 48974
rect 32956 47570 33012 48076
rect 32956 47518 32958 47570
rect 33010 47518 33012 47570
rect 32956 47506 33012 47518
rect 32620 46898 32676 46956
rect 32620 46846 32622 46898
rect 32674 46846 32676 46898
rect 32620 46834 32676 46846
rect 33180 47458 33236 47470
rect 33180 47406 33182 47458
rect 33234 47406 33236 47458
rect 32508 46050 32564 46060
rect 33068 45780 33124 45790
rect 32172 45574 32228 45612
rect 32844 45668 32900 45678
rect 32060 45332 32116 45342
rect 32060 45106 32116 45276
rect 32060 45054 32062 45106
rect 32114 45054 32116 45106
rect 32060 45042 32116 45054
rect 32508 44996 32564 45006
rect 32172 43652 32228 43662
rect 31948 43596 32172 43652
rect 31948 43428 32004 43596
rect 32172 43586 32228 43596
rect 31948 43362 32004 43372
rect 31612 43262 31614 43314
rect 31666 43262 31668 43314
rect 31388 40238 31390 40290
rect 31442 40238 31444 40290
rect 31388 40226 31444 40238
rect 31500 40514 31556 40526
rect 31500 40462 31502 40514
rect 31554 40462 31556 40514
rect 31500 38948 31556 40462
rect 31500 38882 31556 38892
rect 31276 38836 31332 38846
rect 31052 38612 31220 38668
rect 30716 37154 31108 37156
rect 30716 37102 30718 37154
rect 30770 37102 31108 37154
rect 30716 37100 31108 37102
rect 30716 37090 30772 37100
rect 30492 36876 30996 36932
rect 30436 36652 30660 36708
rect 30380 36642 30436 36652
rect 30044 36542 30046 36594
rect 30098 36542 30100 36594
rect 30044 36530 30100 36542
rect 29932 36430 29934 36482
rect 29986 36430 29988 36482
rect 29932 35140 29988 36430
rect 30268 36484 30324 36494
rect 30156 36372 30212 36382
rect 30156 36278 30212 36316
rect 30268 35698 30324 36428
rect 30268 35646 30270 35698
rect 30322 35646 30324 35698
rect 30268 35634 30324 35646
rect 30380 35588 30436 35598
rect 30380 35494 30436 35532
rect 30492 35476 30548 35486
rect 29932 35084 30212 35140
rect 30044 34916 30100 34926
rect 30044 34822 30100 34860
rect 29708 34804 29764 34814
rect 29708 34356 29764 34748
rect 29932 34690 29988 34702
rect 29932 34638 29934 34690
rect 29986 34638 29988 34690
rect 29820 34356 29876 34366
rect 29708 34354 29876 34356
rect 29708 34302 29822 34354
rect 29874 34302 29876 34354
rect 29708 34300 29876 34302
rect 29820 34290 29876 34300
rect 29932 34132 29988 34638
rect 29372 34076 29540 34132
rect 28924 29922 28980 29932
rect 29036 32956 29316 33012
rect 28700 27794 28756 27804
rect 28588 27746 28644 27758
rect 28588 27694 28590 27746
rect 28642 27694 28644 27746
rect 28588 27524 28644 27694
rect 28588 27458 28644 27468
rect 28700 27186 28756 27198
rect 28700 27134 28702 27186
rect 28754 27134 28756 27186
rect 28700 27076 28756 27134
rect 28700 27010 28756 27020
rect 28812 26964 28868 26974
rect 28476 26852 28644 26908
rect 27468 26126 27470 26178
rect 27522 26126 27524 26178
rect 27468 26114 27524 26126
rect 27580 26290 27636 26302
rect 27580 26238 27582 26290
rect 27634 26238 27636 26290
rect 27580 26180 27636 26238
rect 27580 26114 27636 26124
rect 27244 26012 27412 26068
rect 27132 26002 27188 26012
rect 26460 25666 26516 25676
rect 26796 25788 26964 25844
rect 26124 25566 26126 25618
rect 26178 25566 26180 25618
rect 26124 25554 26180 25566
rect 26796 25396 26852 25788
rect 26908 25620 26964 25630
rect 26908 25618 27300 25620
rect 26908 25566 26910 25618
rect 26962 25566 27300 25618
rect 26908 25564 27300 25566
rect 26908 25554 26964 25564
rect 27244 25508 27300 25564
rect 27244 25442 27300 25452
rect 27356 25506 27412 26012
rect 27356 25454 27358 25506
rect 27410 25454 27412 25506
rect 26796 25340 26908 25396
rect 26460 25284 26516 25294
rect 26852 25284 26908 25340
rect 26852 25228 26964 25284
rect 26348 24834 26404 24846
rect 26348 24782 26350 24834
rect 26402 24782 26404 24834
rect 26236 24724 26292 24734
rect 26236 24630 26292 24668
rect 25900 24098 25956 24108
rect 26236 24500 26292 24510
rect 26012 23940 26068 23950
rect 25788 22430 25790 22482
rect 25842 22430 25844 22482
rect 25788 22418 25844 22430
rect 25900 23938 26068 23940
rect 25900 23886 26014 23938
rect 26066 23886 26068 23938
rect 25900 23884 26068 23886
rect 25900 22932 25956 23884
rect 26012 23874 26068 23884
rect 26124 23268 26180 23278
rect 26124 23174 26180 23212
rect 25900 22370 25956 22876
rect 25900 22318 25902 22370
rect 25954 22318 25956 22370
rect 25900 22306 25956 22318
rect 26012 23154 26068 23166
rect 26012 23102 26014 23154
rect 26066 23102 26068 23154
rect 26012 22260 26068 23102
rect 26236 22708 26292 24444
rect 26348 23268 26404 24782
rect 26348 23202 26404 23212
rect 26236 22652 26404 22708
rect 25676 22204 25844 22260
rect 25116 21746 25172 21756
rect 25676 21812 25732 21822
rect 25676 21718 25732 21756
rect 24668 21534 24670 21586
rect 24722 21534 24724 21586
rect 24668 20244 24724 21534
rect 24668 20178 24724 20188
rect 24892 21532 25060 21588
rect 24892 20132 24948 21532
rect 25788 20916 25844 22204
rect 26012 22194 26068 22204
rect 26236 22260 26292 22270
rect 26012 21028 26068 21038
rect 25900 20916 25956 20926
rect 25788 20914 25956 20916
rect 25788 20862 25902 20914
rect 25954 20862 25956 20914
rect 25788 20860 25956 20862
rect 25900 20850 25956 20860
rect 25004 20692 25060 20702
rect 25004 20598 25060 20636
rect 25452 20580 25508 20590
rect 25452 20486 25508 20524
rect 26012 20580 26068 20972
rect 25116 20468 25172 20478
rect 25004 20132 25060 20142
rect 24892 20130 25060 20132
rect 24892 20078 25006 20130
rect 25058 20078 25060 20130
rect 24892 20076 25060 20078
rect 25004 20066 25060 20076
rect 24892 19236 24948 19246
rect 24444 17838 24446 17890
rect 24498 17838 24500 17890
rect 24444 17826 24500 17838
rect 24556 19124 24612 19134
rect 24556 18450 24612 19068
rect 24556 18398 24558 18450
rect 24610 18398 24612 18450
rect 24444 17668 24500 17678
rect 24332 17666 24500 17668
rect 24332 17614 24446 17666
rect 24498 17614 24500 17666
rect 24332 17612 24500 17614
rect 24444 17602 24500 17612
rect 23996 17054 23998 17106
rect 24050 17054 24052 17106
rect 23996 17042 24052 17054
rect 24108 16996 24164 17006
rect 24108 16548 24164 16940
rect 24444 16996 24500 17006
rect 24556 16996 24612 18398
rect 24780 18564 24836 18574
rect 24780 18450 24836 18508
rect 24780 18398 24782 18450
rect 24834 18398 24836 18450
rect 24780 18386 24836 18398
rect 24892 18450 24948 19180
rect 25004 19234 25060 19246
rect 25004 19182 25006 19234
rect 25058 19182 25060 19234
rect 25004 18676 25060 19182
rect 25004 18610 25060 18620
rect 24892 18398 24894 18450
rect 24946 18398 24948 18450
rect 24892 18386 24948 18398
rect 24892 17780 24948 17790
rect 25116 17780 25172 20412
rect 25676 19906 25732 19918
rect 25676 19854 25678 19906
rect 25730 19854 25732 19906
rect 25676 19572 25732 19854
rect 25676 19124 25732 19516
rect 26012 19906 26068 20524
rect 26012 19854 26014 19906
rect 26066 19854 26068 19906
rect 26012 19124 26068 19854
rect 26124 19124 26180 19134
rect 26012 19122 26180 19124
rect 26012 19070 26126 19122
rect 26178 19070 26180 19122
rect 26012 19068 26180 19070
rect 25676 19058 25732 19068
rect 25676 18676 25732 18686
rect 25676 18582 25732 18620
rect 25900 18564 25956 18574
rect 25900 18470 25956 18508
rect 25788 18338 25844 18350
rect 25788 18286 25790 18338
rect 25842 18286 25844 18338
rect 24892 17778 25172 17780
rect 24892 17726 24894 17778
rect 24946 17726 25172 17778
rect 24892 17724 25172 17726
rect 25340 17778 25396 17790
rect 25340 17726 25342 17778
rect 25394 17726 25396 17778
rect 24892 17714 24948 17724
rect 25340 17668 25396 17726
rect 25340 17602 25396 17612
rect 25676 17668 25732 17678
rect 25676 17574 25732 17612
rect 25004 17108 25060 17118
rect 25004 17014 25060 17052
rect 25788 16996 25844 18286
rect 24500 16940 24612 16996
rect 25564 16940 25844 16996
rect 25900 17554 25956 17566
rect 25900 17502 25902 17554
rect 25954 17502 25956 17554
rect 24444 16902 24500 16940
rect 23660 16210 23828 16212
rect 23660 16158 23662 16210
rect 23714 16158 23828 16210
rect 23660 16156 23828 16158
rect 23996 16492 24164 16548
rect 23660 16146 23716 16156
rect 23884 16100 23940 16110
rect 23884 15426 23940 16044
rect 23884 15374 23886 15426
rect 23938 15374 23940 15426
rect 23772 15316 23828 15326
rect 23772 15222 23828 15260
rect 23884 15148 23940 15374
rect 23548 15092 23940 15148
rect 23436 13972 23492 13982
rect 23548 13972 23604 15092
rect 23884 14644 23940 14654
rect 23996 14644 24052 16492
rect 24892 16212 24948 16222
rect 24892 16118 24948 16156
rect 25340 15986 25396 15998
rect 25340 15934 25342 15986
rect 25394 15934 25396 15986
rect 24444 15874 24500 15886
rect 24444 15822 24446 15874
rect 24498 15822 24500 15874
rect 24444 15428 24500 15822
rect 24556 15540 24612 15550
rect 24556 15446 24612 15484
rect 24444 15362 24500 15372
rect 24892 15428 24948 15438
rect 24892 15334 24948 15372
rect 23884 14642 24052 14644
rect 23884 14590 23886 14642
rect 23938 14590 24052 14642
rect 23884 14588 24052 14590
rect 24108 15316 24164 15326
rect 23884 14578 23940 14588
rect 23436 13970 23604 13972
rect 23436 13918 23438 13970
rect 23490 13918 23604 13970
rect 23436 13916 23604 13918
rect 23436 13188 23492 13916
rect 23436 13122 23492 13132
rect 23660 13074 23716 13086
rect 23660 13022 23662 13074
rect 23714 13022 23716 13074
rect 23380 12572 23604 12628
rect 23324 12562 23380 12572
rect 23324 12404 23380 12414
rect 23100 12402 23380 12404
rect 23100 12350 23326 12402
rect 23378 12350 23380 12402
rect 23100 12348 23380 12350
rect 23324 12338 23380 12348
rect 23548 12402 23604 12572
rect 23548 12350 23550 12402
rect 23602 12350 23604 12402
rect 23548 12338 23604 12350
rect 22876 12292 22932 12302
rect 22876 12198 22932 12236
rect 23660 12292 23716 13022
rect 23660 12160 23716 12236
rect 22652 11442 22708 11452
rect 23212 11508 23268 11518
rect 23212 11414 23268 11452
rect 22092 11396 22148 11406
rect 21980 11394 22148 11396
rect 21980 11342 22094 11394
rect 22146 11342 22148 11394
rect 21980 11340 22148 11342
rect 21980 10500 22036 11340
rect 22092 11330 22148 11340
rect 22428 11394 22484 11406
rect 22428 11342 22430 11394
rect 22482 11342 22484 11394
rect 22428 10836 22484 11342
rect 22092 10780 22484 10836
rect 22764 11282 22820 11294
rect 22764 11230 22766 11282
rect 22818 11230 22820 11282
rect 22092 10722 22148 10780
rect 22092 10670 22094 10722
rect 22146 10670 22148 10722
rect 22092 10612 22148 10670
rect 22092 10546 22148 10556
rect 22652 10612 22708 10622
rect 21980 10434 22036 10444
rect 22540 10500 22596 10510
rect 21868 9268 21924 9278
rect 22540 9268 22596 10444
rect 22652 9826 22708 10556
rect 22764 9938 22820 11230
rect 23548 10724 23604 10734
rect 22988 10500 23044 10510
rect 22988 10050 23044 10444
rect 22988 9998 22990 10050
rect 23042 9998 23044 10050
rect 22988 9986 23044 9998
rect 22764 9886 22766 9938
rect 22818 9886 22820 9938
rect 22764 9874 22820 9886
rect 23548 9938 23604 10668
rect 23772 10724 23828 10734
rect 23772 10630 23828 10668
rect 23660 10612 23716 10622
rect 23660 10518 23716 10556
rect 23548 9886 23550 9938
rect 23602 9886 23604 9938
rect 22652 9774 22654 9826
rect 22706 9774 22708 9826
rect 22652 9762 22708 9774
rect 23548 9716 23604 9886
rect 23548 9650 23604 9660
rect 22652 9268 22708 9278
rect 22540 9266 22708 9268
rect 22540 9214 22654 9266
rect 22706 9214 22708 9266
rect 22540 9212 22708 9214
rect 21868 9174 21924 9212
rect 22652 9202 22708 9212
rect 23100 9268 23156 9278
rect 22988 9154 23044 9166
rect 22988 9102 22990 9154
rect 23042 9102 23044 9154
rect 21980 9042 22036 9054
rect 21980 8990 21982 9042
rect 22034 8990 22036 9042
rect 21980 8820 22036 8990
rect 21980 8754 22036 8764
rect 22540 9042 22596 9054
rect 22540 8990 22542 9042
rect 22594 8990 22596 9042
rect 21980 8146 22036 8158
rect 21980 8094 21982 8146
rect 22034 8094 22036 8146
rect 21980 7700 22036 8094
rect 22092 7700 22148 7710
rect 21980 7698 22148 7700
rect 21980 7646 22094 7698
rect 22146 7646 22148 7698
rect 21980 7644 22148 7646
rect 22092 7634 22148 7644
rect 22204 7586 22260 7598
rect 22204 7534 22206 7586
rect 22258 7534 22260 7586
rect 22204 7476 22260 7534
rect 22204 7410 22260 7420
rect 22540 7476 22596 8990
rect 22764 9042 22820 9054
rect 22764 8990 22766 9042
rect 22818 8990 22820 9042
rect 22652 8820 22708 8830
rect 22652 8258 22708 8764
rect 22764 8428 22820 8990
rect 22764 8372 22932 8428
rect 22876 8370 22932 8372
rect 22876 8318 22878 8370
rect 22930 8318 22932 8370
rect 22876 8306 22932 8318
rect 22652 8206 22654 8258
rect 22706 8206 22708 8258
rect 22652 8194 22708 8206
rect 22988 7812 23044 9102
rect 22876 7756 23044 7812
rect 23100 8146 23156 9212
rect 23548 9268 23604 9278
rect 23548 9174 23604 9212
rect 23996 8930 24052 8942
rect 23996 8878 23998 8930
rect 24050 8878 24052 8930
rect 23436 8820 23492 8830
rect 23100 8094 23102 8146
rect 23154 8094 23156 8146
rect 22876 7698 22932 7756
rect 22876 7646 22878 7698
rect 22930 7646 22932 7698
rect 22876 7634 22932 7646
rect 22988 7588 23044 7598
rect 22988 7494 23044 7532
rect 23100 7476 23156 8094
rect 23324 8260 23380 8270
rect 23324 7700 23380 8204
rect 23324 7634 23380 7644
rect 23436 7586 23492 8764
rect 23996 8428 24052 8878
rect 23884 8372 24052 8428
rect 23884 8260 23940 8372
rect 23884 8194 23940 8204
rect 23996 8148 24052 8158
rect 23996 8054 24052 8092
rect 23436 7534 23438 7586
rect 23490 7534 23492 7586
rect 23436 7522 23492 7534
rect 23212 7476 23268 7486
rect 23100 7474 23380 7476
rect 23100 7422 23214 7474
rect 23266 7422 23380 7474
rect 23100 7420 23380 7422
rect 22540 7410 22596 7420
rect 23212 7410 23268 7420
rect 21756 6626 21812 6636
rect 22540 6692 22596 6702
rect 20300 6580 20356 6590
rect 20300 6486 20356 6524
rect 21980 6580 22036 6590
rect 21980 6486 22036 6524
rect 21644 6466 21700 6478
rect 21644 6414 21646 6466
rect 21698 6414 21700 6466
rect 20524 6132 20580 6142
rect 20188 6130 20580 6132
rect 20188 6078 20526 6130
rect 20578 6078 20580 6130
rect 20188 6076 20580 6078
rect 20524 6066 20580 6076
rect 20188 5796 20244 5806
rect 19852 5684 19908 5694
rect 19852 5234 19908 5628
rect 20188 5460 20244 5740
rect 20188 5394 20244 5404
rect 20300 5684 20356 5694
rect 21308 5684 21364 5694
rect 19852 5182 19854 5234
rect 19906 5182 19908 5234
rect 19852 5170 19908 5182
rect 20300 5124 20356 5628
rect 20300 5030 20356 5068
rect 20860 5682 21364 5684
rect 20860 5630 21310 5682
rect 21362 5630 21364 5682
rect 20860 5628 21364 5630
rect 20860 5122 20916 5628
rect 21308 5618 21364 5628
rect 21644 5348 21700 6414
rect 22540 6356 22596 6636
rect 23100 6692 23156 6702
rect 22988 6468 23044 6478
rect 22988 6374 23044 6412
rect 22540 6290 22596 6300
rect 21980 6018 22036 6030
rect 21980 5966 21982 6018
rect 22034 5966 22036 6018
rect 21980 5908 22036 5966
rect 23100 6018 23156 6636
rect 23100 5966 23102 6018
rect 23154 5966 23156 6018
rect 22204 5908 22260 5918
rect 21980 5842 22036 5852
rect 22092 5906 22260 5908
rect 22092 5854 22206 5906
rect 22258 5854 22260 5906
rect 22092 5852 22260 5854
rect 22092 5348 22148 5852
rect 22204 5842 22260 5852
rect 23100 5908 23156 5966
rect 23100 5842 23156 5852
rect 23212 6356 23268 6366
rect 21644 5282 21700 5292
rect 21980 5292 22148 5348
rect 20860 5070 20862 5122
rect 20914 5070 20916 5122
rect 20860 5058 20916 5070
rect 21868 5012 21924 5022
rect 21868 4918 21924 4956
rect 21980 4898 22036 5292
rect 21980 4846 21982 4898
rect 22034 4846 22036 4898
rect 21980 4834 22036 4846
rect 22876 5124 22932 5134
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19628 4498 19684 4508
rect 20748 4562 20804 4574
rect 20748 4510 20750 4562
rect 20802 4510 20804 4562
rect 18228 3612 18340 3668
rect 19628 3668 19684 3678
rect 18172 3574 18228 3612
rect 19628 3574 19684 3612
rect 20748 3668 20804 4510
rect 21756 4564 21812 4574
rect 21756 4450 21812 4508
rect 21756 4398 21758 4450
rect 21810 4398 21812 4450
rect 21756 4386 21812 4398
rect 21308 4340 21364 4350
rect 21308 4246 21364 4284
rect 21532 4340 21588 4350
rect 20748 3602 20804 3612
rect 17948 3490 18004 3500
rect 18620 3556 18676 3566
rect 18620 3462 18676 3500
rect 21308 3556 21364 3566
rect 21308 3462 21364 3500
rect 21532 3442 21588 4284
rect 22204 4340 22260 4350
rect 22204 4246 22260 4284
rect 21644 4228 21700 4238
rect 21644 3554 21700 4172
rect 22652 4228 22708 4238
rect 22652 4134 22708 4172
rect 22092 3668 22148 3678
rect 22092 3574 22148 3612
rect 22876 3666 22932 5068
rect 23100 5122 23156 5134
rect 23100 5070 23102 5122
rect 23154 5070 23156 5122
rect 23100 4564 23156 5070
rect 23212 5124 23268 6300
rect 23324 6132 23380 7420
rect 23996 6578 24052 6590
rect 23996 6526 23998 6578
rect 24050 6526 24052 6578
rect 23436 6468 23492 6478
rect 23436 6132 23492 6412
rect 23324 6130 23492 6132
rect 23324 6078 23326 6130
rect 23378 6078 23492 6130
rect 23324 6076 23492 6078
rect 23324 6066 23380 6076
rect 23212 5010 23268 5068
rect 23212 4958 23214 5010
rect 23266 4958 23268 5010
rect 23212 4946 23268 4958
rect 23212 4564 23268 4574
rect 23100 4562 23268 4564
rect 23100 4510 23214 4562
rect 23266 4510 23268 4562
rect 23100 4508 23268 4510
rect 23212 4498 23268 4508
rect 23436 4562 23492 6076
rect 23548 6356 23604 6366
rect 23548 6130 23604 6300
rect 23996 6356 24052 6526
rect 23996 6290 24052 6300
rect 23548 6078 23550 6130
rect 23602 6078 23604 6130
rect 23548 6066 23604 6078
rect 23436 4510 23438 4562
rect 23490 4510 23492 4562
rect 22876 3614 22878 3666
rect 22930 3614 22932 3666
rect 22876 3602 22932 3614
rect 23324 3668 23380 3678
rect 23436 3668 23492 4510
rect 23548 5908 23604 5918
rect 23548 4450 23604 5852
rect 23660 5908 23716 5918
rect 23996 5908 24052 5918
rect 23660 5906 24052 5908
rect 23660 5854 23662 5906
rect 23714 5854 23998 5906
rect 24050 5854 24052 5906
rect 23660 5852 24052 5854
rect 23660 5842 23716 5852
rect 23996 5842 24052 5852
rect 24108 4900 24164 15260
rect 25340 15148 25396 15934
rect 25564 15148 25620 16940
rect 25676 16772 25732 16782
rect 25676 16212 25732 16716
rect 25676 16146 25732 16156
rect 25900 15540 25956 17502
rect 26012 16884 26068 16894
rect 26012 16098 26068 16828
rect 26124 16772 26180 19068
rect 26236 17106 26292 22204
rect 26348 21588 26404 22652
rect 26348 21494 26404 21532
rect 26460 20916 26516 25228
rect 26796 24052 26852 24062
rect 26796 23958 26852 23996
rect 26796 23828 26852 23838
rect 26572 23380 26628 23390
rect 26572 23286 26628 23324
rect 26684 21586 26740 21598
rect 26684 21534 26686 21586
rect 26738 21534 26740 21586
rect 26684 21476 26740 21534
rect 26684 21410 26740 21420
rect 26572 20916 26628 20926
rect 26460 20914 26628 20916
rect 26460 20862 26574 20914
rect 26626 20862 26628 20914
rect 26460 20860 26628 20862
rect 26572 20850 26628 20860
rect 26684 20916 26740 20926
rect 26796 20916 26852 23772
rect 26908 23716 26964 25228
rect 26908 23660 27188 23716
rect 26908 23492 26964 23502
rect 26908 23044 26964 23436
rect 26908 21476 26964 22988
rect 26908 21420 27076 21476
rect 26684 20914 26852 20916
rect 26684 20862 26686 20914
rect 26738 20862 26852 20914
rect 26684 20860 26852 20862
rect 26684 20850 26740 20860
rect 26460 20692 26516 20702
rect 26348 20690 26516 20692
rect 26348 20638 26462 20690
rect 26514 20638 26516 20690
rect 26348 20636 26516 20638
rect 26348 19572 26404 20636
rect 26460 20626 26516 20636
rect 26796 20468 26852 20860
rect 26908 20802 26964 20814
rect 26908 20750 26910 20802
rect 26962 20750 26964 20802
rect 26908 20580 26964 20750
rect 26908 20514 26964 20524
rect 27020 20468 27076 21420
rect 27132 21028 27188 23660
rect 27356 23492 27412 25454
rect 27468 25956 27524 25966
rect 27468 24612 27524 25900
rect 27580 24836 27636 24846
rect 27580 24742 27636 24780
rect 27468 24556 27636 24612
rect 27356 23426 27412 23436
rect 27468 23938 27524 23950
rect 27468 23886 27470 23938
rect 27522 23886 27524 23938
rect 27356 23268 27412 23278
rect 27356 22482 27412 23212
rect 27468 23156 27524 23886
rect 27468 23024 27524 23100
rect 27580 22932 27636 24556
rect 27916 24500 27972 26572
rect 28140 24724 28196 26852
rect 28588 26514 28644 26852
rect 28588 26462 28590 26514
rect 28642 26462 28644 26514
rect 28588 26450 28644 26462
rect 28700 26852 28868 26908
rect 29036 26908 29092 32956
rect 29372 31220 29428 31230
rect 29372 31106 29428 31164
rect 29372 31054 29374 31106
rect 29426 31054 29428 31106
rect 29372 31042 29428 31054
rect 29260 30212 29316 30222
rect 29148 29540 29204 29550
rect 29148 29446 29204 29484
rect 29036 26852 29204 26908
rect 28252 26290 28308 26302
rect 28252 26238 28254 26290
rect 28306 26238 28308 26290
rect 28252 25620 28308 26238
rect 28364 26290 28420 26302
rect 28364 26238 28366 26290
rect 28418 26238 28420 26290
rect 28364 25956 28420 26238
rect 28700 26290 28756 26852
rect 28700 26238 28702 26290
rect 28754 26238 28756 26290
rect 28476 26180 28532 26190
rect 28476 26086 28532 26124
rect 28364 25890 28420 25900
rect 28252 25564 28532 25620
rect 28476 25508 28532 25564
rect 28252 25394 28308 25406
rect 28252 25342 28254 25394
rect 28306 25342 28308 25394
rect 28252 25060 28308 25342
rect 28252 24994 28308 25004
rect 28364 24724 28420 24734
rect 28140 24722 28420 24724
rect 28140 24670 28366 24722
rect 28418 24670 28420 24722
rect 28140 24668 28420 24670
rect 28028 24500 28084 24510
rect 27916 24444 28028 24500
rect 27356 22430 27358 22482
rect 27410 22430 27412 22482
rect 27356 22418 27412 22430
rect 27468 22876 27636 22932
rect 28028 23938 28084 24444
rect 28028 23886 28030 23938
rect 28082 23886 28084 23938
rect 27468 21700 27524 22876
rect 27580 22370 27636 22382
rect 27580 22318 27582 22370
rect 27634 22318 27636 22370
rect 27580 22260 27636 22318
rect 27580 22194 27636 22204
rect 27916 22260 27972 22270
rect 27916 22166 27972 22204
rect 28028 22036 28084 23886
rect 27468 21634 27524 21644
rect 27580 21980 28084 22036
rect 28364 23826 28420 24668
rect 28476 24276 28532 25452
rect 28588 24500 28644 24510
rect 28588 24406 28644 24444
rect 28476 24220 28644 24276
rect 28476 24050 28532 24062
rect 28476 23998 28478 24050
rect 28530 23998 28532 24050
rect 28476 23940 28532 23998
rect 28476 23874 28532 23884
rect 28364 23774 28366 23826
rect 28418 23774 28420 23826
rect 27132 20962 27188 20972
rect 27356 20804 27412 20814
rect 27132 20692 27188 20702
rect 27188 20636 27300 20692
rect 27132 20598 27188 20636
rect 27020 20412 27188 20468
rect 26796 20402 26852 20412
rect 26908 20356 26964 20366
rect 26460 19906 26516 19918
rect 26460 19854 26462 19906
rect 26514 19854 26516 19906
rect 26460 19796 26516 19854
rect 26516 19740 26628 19796
rect 26460 19730 26516 19740
rect 26348 19506 26404 19516
rect 26460 19346 26516 19358
rect 26460 19294 26462 19346
rect 26514 19294 26516 19346
rect 26460 19236 26516 19294
rect 26460 19170 26516 19180
rect 26572 19012 26628 19740
rect 26572 18946 26628 18956
rect 26908 18788 26964 20300
rect 27132 19346 27188 20412
rect 27244 20356 27300 20636
rect 27244 20290 27300 20300
rect 27132 19294 27134 19346
rect 27186 19294 27188 19346
rect 27132 19282 27188 19294
rect 27244 20132 27300 20142
rect 26796 18732 26964 18788
rect 27020 19236 27076 19246
rect 26572 18676 26628 18686
rect 26348 18452 26404 18462
rect 26348 18358 26404 18396
rect 26572 17778 26628 18620
rect 26796 18340 26852 18732
rect 27020 18676 27076 19180
rect 27244 19012 27300 20076
rect 27244 18946 27300 18956
rect 26908 18564 26964 18574
rect 27020 18544 27076 18620
rect 26908 18470 26964 18508
rect 27356 18452 27412 20748
rect 27580 19346 27636 21980
rect 27804 21476 27860 21486
rect 27580 19294 27582 19346
rect 27634 19294 27636 19346
rect 27580 19282 27636 19294
rect 27692 21474 27860 21476
rect 27692 21422 27806 21474
rect 27858 21422 27860 21474
rect 27692 21420 27860 21422
rect 27244 18396 27412 18452
rect 27468 18564 27524 18574
rect 26796 18284 26964 18340
rect 26572 17726 26574 17778
rect 26626 17726 26628 17778
rect 26572 17714 26628 17726
rect 26236 17054 26238 17106
rect 26290 17054 26292 17106
rect 26236 17042 26292 17054
rect 26348 17666 26404 17678
rect 26348 17614 26350 17666
rect 26402 17614 26404 17666
rect 26124 16706 26180 16716
rect 26236 16212 26292 16222
rect 26348 16212 26404 17614
rect 26684 17666 26740 17678
rect 26684 17614 26686 17666
rect 26738 17614 26740 17666
rect 26236 16210 26404 16212
rect 26236 16158 26238 16210
rect 26290 16158 26404 16210
rect 26236 16156 26404 16158
rect 26236 16146 26292 16156
rect 26012 16046 26014 16098
rect 26066 16046 26068 16098
rect 26012 16034 26068 16046
rect 25676 15316 25732 15326
rect 25676 15222 25732 15260
rect 24220 15092 24276 15102
rect 24220 14306 24276 15036
rect 25116 15092 25396 15148
rect 25452 15092 25620 15148
rect 25900 15148 25956 15484
rect 26236 15540 26292 15550
rect 26236 15446 26292 15484
rect 25900 15092 26292 15148
rect 25116 14530 25172 15092
rect 25116 14478 25118 14530
rect 25170 14478 25172 14530
rect 25116 14466 25172 14478
rect 24220 14254 24222 14306
rect 24274 14254 24276 14306
rect 24220 13524 24276 14254
rect 24780 14306 24836 14318
rect 24780 14254 24782 14306
rect 24834 14254 24836 14306
rect 24220 13458 24276 13468
rect 24332 13746 24388 13758
rect 24332 13694 24334 13746
rect 24386 13694 24388 13746
rect 24332 12740 24388 13694
rect 24780 13748 24836 14254
rect 25452 13748 25508 15092
rect 24780 13682 24836 13692
rect 25228 13692 25508 13748
rect 25564 14420 25620 14430
rect 24892 13634 24948 13646
rect 24892 13582 24894 13634
rect 24946 13582 24948 13634
rect 24892 13524 24948 13582
rect 24892 13458 24948 13468
rect 24780 12852 24836 12862
rect 24780 12758 24836 12796
rect 24220 12738 24388 12740
rect 24220 12686 24334 12738
rect 24386 12686 24388 12738
rect 24220 12684 24388 12686
rect 24220 12404 24276 12684
rect 24332 12674 24388 12684
rect 24220 12338 24276 12348
rect 24332 12292 24388 12302
rect 24332 12198 24388 12236
rect 24444 12066 24500 12078
rect 24444 12014 24446 12066
rect 24498 12014 24500 12066
rect 24444 11620 24500 12014
rect 24668 11620 24724 11630
rect 24444 11618 24724 11620
rect 24444 11566 24670 11618
rect 24722 11566 24724 11618
rect 24444 11564 24724 11566
rect 24668 11554 24724 11564
rect 24220 11172 24276 11182
rect 24780 11172 24836 11182
rect 24220 11170 24724 11172
rect 24220 11118 24222 11170
rect 24274 11118 24724 11170
rect 24220 11116 24724 11118
rect 24220 11106 24276 11116
rect 24444 10948 24500 10958
rect 24444 10834 24500 10892
rect 24444 10782 24446 10834
rect 24498 10782 24500 10834
rect 24444 10770 24500 10782
rect 24668 10948 24724 11116
rect 24780 11078 24836 11116
rect 25004 11170 25060 11182
rect 25004 11118 25006 11170
rect 25058 11118 25060 11170
rect 25004 10948 25060 11118
rect 24668 10892 25060 10948
rect 24668 10610 24724 10892
rect 24668 10558 24670 10610
rect 24722 10558 24724 10610
rect 24332 10500 24388 10510
rect 24332 10406 24388 10444
rect 24668 9268 24724 10558
rect 25004 10610 25060 10622
rect 25004 10558 25006 10610
rect 25058 10558 25060 10610
rect 25004 9940 25060 10558
rect 25004 9874 25060 9884
rect 24668 9202 24724 9212
rect 25116 9602 25172 9614
rect 25116 9550 25118 9602
rect 25170 9550 25172 9602
rect 25116 9268 25172 9550
rect 25116 9202 25172 9212
rect 24220 8258 24276 8270
rect 24220 8206 24222 8258
rect 24274 8206 24276 8258
rect 24220 7476 24276 8206
rect 24668 8258 24724 8270
rect 24668 8206 24670 8258
rect 24722 8206 24724 8258
rect 24668 7588 24724 8206
rect 24668 7494 24724 7532
rect 24892 8036 24948 8046
rect 24892 7586 24948 7980
rect 24892 7534 24894 7586
rect 24946 7534 24948 7586
rect 24892 7522 24948 7534
rect 24444 7476 24500 7486
rect 24220 7474 24388 7476
rect 24220 7422 24222 7474
rect 24274 7422 24388 7474
rect 24220 7420 24388 7422
rect 24220 7410 24276 7420
rect 24220 6578 24276 6590
rect 24220 6526 24222 6578
rect 24274 6526 24276 6578
rect 24220 6468 24276 6526
rect 24220 6020 24276 6412
rect 24220 5954 24276 5964
rect 24332 5908 24388 7420
rect 24444 7382 24500 7420
rect 24668 6692 24724 6702
rect 24668 6598 24724 6636
rect 24780 6580 24836 6590
rect 24444 6466 24500 6478
rect 24444 6414 24446 6466
rect 24498 6414 24500 6466
rect 24444 6130 24500 6414
rect 24444 6078 24446 6130
rect 24498 6078 24500 6130
rect 24444 6066 24500 6078
rect 24556 5908 24612 5918
rect 24332 5906 24612 5908
rect 24332 5854 24558 5906
rect 24610 5854 24612 5906
rect 24332 5852 24612 5854
rect 24556 5842 24612 5852
rect 24668 5906 24724 5918
rect 24668 5854 24670 5906
rect 24722 5854 24724 5906
rect 24108 4562 24164 4844
rect 24108 4510 24110 4562
rect 24162 4510 24164 4562
rect 24108 4498 24164 4510
rect 24556 5348 24612 5358
rect 24556 4562 24612 5292
rect 24556 4510 24558 4562
rect 24610 4510 24612 4562
rect 24556 4498 24612 4510
rect 24668 5012 24724 5854
rect 24780 5234 24836 6524
rect 24780 5182 24782 5234
rect 24834 5182 24836 5234
rect 24780 5170 24836 5182
rect 25228 5236 25284 13692
rect 25452 13524 25508 13534
rect 25452 13074 25508 13468
rect 25452 13022 25454 13074
rect 25506 13022 25508 13074
rect 25452 13010 25508 13022
rect 25340 11396 25396 11406
rect 25340 11302 25396 11340
rect 25564 10834 25620 14364
rect 26124 14420 26180 14430
rect 25900 14308 25956 14318
rect 25900 14214 25956 14252
rect 26124 13746 26180 14364
rect 26124 13694 26126 13746
rect 26178 13694 26180 13746
rect 26124 13524 26180 13694
rect 26012 12404 26068 12414
rect 26124 12404 26180 13468
rect 26236 12516 26292 15092
rect 26348 14644 26404 16156
rect 26572 17556 26628 17566
rect 26572 15538 26628 17500
rect 26684 16884 26740 17614
rect 26684 16790 26740 16828
rect 26572 15486 26574 15538
rect 26626 15486 26628 15538
rect 26572 15148 26628 15486
rect 26908 15540 26964 18284
rect 27132 18226 27188 18238
rect 27132 18174 27134 18226
rect 27186 18174 27188 18226
rect 27132 17668 27188 18174
rect 27132 17602 27188 17612
rect 27020 17554 27076 17566
rect 27020 17502 27022 17554
rect 27074 17502 27076 17554
rect 27020 17108 27076 17502
rect 27244 17108 27300 18396
rect 27020 17042 27076 17052
rect 27132 17052 27300 17108
rect 26908 15474 26964 15484
rect 27020 15652 27076 15662
rect 27020 15538 27076 15596
rect 27020 15486 27022 15538
rect 27074 15486 27076 15538
rect 27020 15428 27076 15486
rect 27020 15362 27076 15372
rect 27132 15316 27188 17052
rect 27468 16996 27524 18508
rect 27580 18452 27636 18462
rect 27580 18358 27636 18396
rect 27692 18228 27748 21420
rect 27804 21410 27860 21420
rect 28364 21474 28420 23774
rect 28588 23716 28644 24220
rect 28476 23660 28644 23716
rect 28476 22482 28532 23660
rect 28476 22430 28478 22482
rect 28530 22430 28532 22482
rect 28476 22418 28532 22430
rect 28700 21700 28756 26238
rect 29148 26180 29204 26852
rect 29148 25620 29204 26124
rect 29148 25554 29204 25564
rect 28924 24500 28980 24510
rect 28924 24498 29092 24500
rect 28924 24446 28926 24498
rect 28978 24446 29092 24498
rect 28924 24444 29092 24446
rect 28924 24434 28980 24444
rect 28812 22148 28868 22158
rect 28812 22054 28868 22092
rect 28924 21700 28980 21710
rect 28364 21422 28366 21474
rect 28418 21422 28420 21474
rect 28364 21364 28420 21422
rect 27916 21308 28420 21364
rect 28588 21698 28980 21700
rect 28588 21646 28926 21698
rect 28978 21646 28980 21698
rect 28588 21644 28980 21646
rect 27804 21028 27860 21038
rect 27804 20802 27860 20972
rect 27804 20750 27806 20802
rect 27858 20750 27860 20802
rect 27804 20738 27860 20750
rect 27804 20132 27860 20142
rect 27804 20038 27860 20076
rect 27804 19572 27860 19582
rect 27804 18674 27860 19516
rect 27916 19012 27972 21308
rect 28588 21028 28644 21644
rect 28924 21634 28980 21644
rect 28476 20972 28644 21028
rect 28700 21028 28756 21038
rect 28364 20804 28420 20814
rect 28252 20802 28420 20804
rect 28252 20750 28366 20802
rect 28418 20750 28420 20802
rect 28252 20748 28420 20750
rect 28140 20690 28196 20702
rect 28140 20638 28142 20690
rect 28194 20638 28196 20690
rect 28140 20356 28196 20638
rect 28140 20290 28196 20300
rect 28028 20132 28084 20170
rect 28028 20066 28084 20076
rect 28028 19908 28084 19918
rect 28028 19124 28084 19852
rect 28140 19908 28196 19918
rect 28252 19908 28308 20748
rect 28364 20738 28420 20748
rect 28364 20580 28420 20590
rect 28364 20486 28420 20524
rect 28140 19906 28308 19908
rect 28140 19854 28142 19906
rect 28194 19854 28308 19906
rect 28140 19852 28308 19854
rect 28364 20356 28420 20366
rect 28140 19842 28196 19852
rect 28364 19348 28420 20300
rect 28476 20132 28532 20972
rect 28588 20804 28644 20814
rect 28588 20710 28644 20748
rect 28700 20244 28756 20972
rect 29036 20916 29092 24444
rect 29260 23042 29316 30156
rect 29484 28420 29540 34076
rect 29932 34066 29988 34076
rect 29820 33908 29876 33918
rect 29820 33458 29876 33852
rect 29820 33406 29822 33458
rect 29874 33406 29876 33458
rect 29820 33394 29876 33406
rect 29596 32564 29652 32574
rect 29596 31666 29652 32508
rect 29932 32562 29988 32574
rect 29932 32510 29934 32562
rect 29986 32510 29988 32562
rect 29932 32452 29988 32510
rect 29932 31778 29988 32396
rect 30156 31948 30212 35084
rect 30380 35026 30436 35038
rect 30380 34974 30382 35026
rect 30434 34974 30436 35026
rect 30268 34916 30324 34926
rect 30380 34916 30436 34974
rect 30268 34914 30436 34916
rect 30268 34862 30270 34914
rect 30322 34862 30436 34914
rect 30268 34860 30436 34862
rect 30268 34850 30324 34860
rect 30380 33906 30436 33918
rect 30380 33854 30382 33906
rect 30434 33854 30436 33906
rect 30380 33796 30436 33854
rect 30380 33730 30436 33740
rect 30380 33236 30436 33246
rect 30156 31892 30324 31948
rect 29932 31726 29934 31778
rect 29986 31726 29988 31778
rect 29932 31714 29988 31726
rect 29596 31614 29598 31666
rect 29650 31614 29652 31666
rect 29596 31602 29652 31614
rect 30156 31554 30212 31566
rect 30156 31502 30158 31554
rect 30210 31502 30212 31554
rect 30156 31108 30212 31502
rect 30156 31042 30212 31052
rect 29820 30770 29876 30782
rect 29820 30718 29822 30770
rect 29874 30718 29876 30770
rect 29596 29988 29652 29998
rect 29596 29894 29652 29932
rect 29820 29652 29876 30718
rect 29820 29586 29876 29596
rect 29932 30772 29988 30782
rect 29820 29316 29876 29326
rect 29820 29222 29876 29260
rect 29932 28868 29988 30716
rect 30156 29540 30212 29550
rect 29820 28812 29988 28868
rect 30044 29316 30100 29326
rect 30044 29092 30100 29260
rect 29484 28364 29652 28420
rect 29372 28084 29428 28094
rect 29372 27990 29428 28028
rect 29484 27300 29540 27310
rect 29484 27186 29540 27244
rect 29484 27134 29486 27186
rect 29538 27134 29540 27186
rect 29484 27122 29540 27134
rect 29484 26404 29540 26414
rect 29484 26310 29540 26348
rect 29372 26292 29428 26302
rect 29372 26178 29428 26236
rect 29372 26126 29374 26178
rect 29426 26126 29428 26178
rect 29372 26114 29428 26126
rect 29260 22990 29262 23042
rect 29314 22990 29316 23042
rect 29148 21812 29204 21822
rect 29148 21718 29204 21756
rect 29260 21700 29316 22990
rect 29260 21634 29316 21644
rect 29372 25956 29428 25966
rect 29372 22148 29428 25900
rect 29596 25956 29652 28364
rect 29708 26292 29764 26302
rect 29708 26198 29764 26236
rect 29596 25890 29652 25900
rect 29820 25844 29876 28812
rect 29932 28532 29988 28542
rect 29932 27858 29988 28476
rect 29932 27806 29934 27858
rect 29986 27806 29988 27858
rect 29932 27794 29988 27806
rect 29932 27188 29988 27198
rect 30044 27188 30100 29036
rect 30156 28644 30212 29484
rect 30268 29204 30324 31892
rect 30380 30548 30436 33180
rect 30492 32562 30548 35420
rect 30604 34354 30660 36652
rect 30828 35812 30884 35822
rect 30828 35718 30884 35756
rect 30828 34916 30884 34926
rect 30604 34302 30606 34354
rect 30658 34302 30660 34354
rect 30604 33908 30660 34302
rect 30604 33842 30660 33852
rect 30716 34914 30884 34916
rect 30716 34862 30830 34914
rect 30882 34862 30884 34914
rect 30716 34860 30884 34862
rect 30716 34802 30772 34860
rect 30828 34850 30884 34860
rect 30716 34750 30718 34802
rect 30770 34750 30772 34802
rect 30716 33906 30772 34750
rect 30716 33854 30718 33906
rect 30770 33854 30772 33906
rect 30716 33234 30772 33854
rect 30716 33182 30718 33234
rect 30770 33182 30772 33234
rect 30716 33170 30772 33182
rect 30492 32510 30494 32562
rect 30546 32510 30548 32562
rect 30492 31556 30548 32510
rect 30828 32674 30884 32686
rect 30828 32622 30830 32674
rect 30882 32622 30884 32674
rect 30828 32564 30884 32622
rect 30828 32498 30884 32508
rect 30828 31668 30884 31678
rect 30940 31668 30996 36876
rect 31052 36706 31108 37100
rect 31052 36654 31054 36706
rect 31106 36654 31108 36706
rect 31052 36642 31108 36654
rect 31052 36258 31108 36270
rect 31052 36206 31054 36258
rect 31106 36206 31108 36258
rect 31052 35700 31108 36206
rect 31052 35634 31108 35644
rect 31052 34916 31108 34926
rect 31052 34822 31108 34860
rect 31164 34914 31220 38612
rect 31276 37380 31332 38780
rect 31500 38724 31556 38800
rect 31388 38610 31444 38622
rect 31388 38558 31390 38610
rect 31442 38558 31444 38610
rect 31388 37604 31444 38558
rect 31388 37538 31444 37548
rect 31276 37324 31444 37380
rect 31276 37156 31332 37166
rect 31276 35028 31332 37100
rect 31276 34962 31332 34972
rect 31164 34862 31166 34914
rect 31218 34862 31220 34914
rect 31164 34804 31220 34862
rect 31164 34738 31220 34748
rect 31388 33572 31444 37324
rect 31500 37266 31556 38668
rect 31500 37214 31502 37266
rect 31554 37214 31556 37266
rect 31500 37202 31556 37214
rect 31612 37828 31668 43262
rect 32508 43316 32564 44940
rect 32844 43540 32900 45612
rect 32956 44996 33012 45006
rect 32956 44902 33012 44940
rect 32844 43538 33012 43540
rect 32844 43486 32846 43538
rect 32898 43486 33012 43538
rect 32844 43484 33012 43486
rect 32844 43474 32900 43484
rect 32956 43428 33012 43484
rect 32956 43362 33012 43372
rect 32508 43222 32564 43260
rect 32844 43316 32900 43326
rect 32844 43222 32900 43260
rect 33068 43092 33124 45724
rect 32844 43036 33124 43092
rect 33180 43988 33236 47406
rect 33292 47124 33348 50372
rect 33628 49252 33684 50428
rect 33852 50370 33908 50382
rect 33852 50318 33854 50370
rect 33906 50318 33908 50370
rect 33852 50036 33908 50318
rect 34076 50148 34132 50652
rect 35868 50708 35924 56252
rect 36092 55972 36148 56814
rect 36316 56866 36372 57036
rect 36316 56814 36318 56866
rect 36370 56814 36372 56866
rect 36316 56308 36372 56814
rect 36540 56866 36596 57148
rect 37436 57092 37492 57486
rect 37436 57026 37492 57036
rect 37548 57428 37604 57438
rect 36540 56814 36542 56866
rect 36594 56814 36596 56866
rect 36540 56802 36596 56814
rect 36428 56756 36484 56766
rect 36428 56662 36484 56700
rect 36316 56242 36372 56252
rect 37212 56644 37268 56654
rect 36092 55906 36148 55916
rect 35980 55410 36036 55422
rect 35980 55358 35982 55410
rect 36034 55358 36036 55410
rect 35980 54514 36036 55358
rect 36316 55188 36372 55198
rect 36316 55094 36372 55132
rect 35980 54462 35982 54514
rect 36034 54462 36036 54514
rect 35980 53842 36036 54462
rect 36540 54516 36596 54526
rect 36540 54514 36708 54516
rect 36540 54462 36542 54514
rect 36594 54462 36708 54514
rect 36540 54460 36708 54462
rect 36540 54450 36596 54460
rect 36428 54402 36484 54414
rect 36428 54350 36430 54402
rect 36482 54350 36484 54402
rect 36204 54292 36260 54302
rect 35980 53790 35982 53842
rect 36034 53790 36036 53842
rect 35980 53778 36036 53790
rect 36092 54290 36260 54292
rect 36092 54238 36206 54290
rect 36258 54238 36260 54290
rect 36092 54236 36260 54238
rect 36092 53620 36148 54236
rect 36204 54226 36260 54236
rect 36428 53730 36484 54350
rect 36428 53678 36430 53730
rect 36482 53678 36484 53730
rect 36428 53666 36484 53678
rect 36092 53554 36148 53564
rect 36204 53618 36260 53630
rect 36204 53566 36206 53618
rect 36258 53566 36260 53618
rect 36204 52948 36260 53566
rect 36652 53508 36708 54460
rect 36540 52948 36596 52958
rect 36204 52946 36596 52948
rect 36204 52894 36542 52946
rect 36594 52894 36596 52946
rect 36204 52892 36596 52894
rect 36540 51604 36596 52892
rect 36540 51538 36596 51548
rect 36652 52834 36708 53452
rect 36652 52782 36654 52834
rect 36706 52782 36708 52834
rect 36652 51602 36708 52782
rect 36652 51550 36654 51602
rect 36706 51550 36708 51602
rect 36652 51538 36708 51550
rect 35868 50642 35924 50652
rect 36204 51378 36260 51390
rect 36204 51326 36206 51378
rect 36258 51326 36260 51378
rect 34076 50082 34132 50092
rect 34188 50484 34244 50494
rect 33852 49970 33908 49980
rect 33964 49924 34020 49934
rect 33964 49812 34020 49868
rect 33852 49810 34020 49812
rect 33852 49758 33966 49810
rect 34018 49758 34020 49810
rect 33852 49756 34020 49758
rect 33628 49196 33796 49252
rect 33628 48804 33684 48814
rect 33628 48354 33684 48748
rect 33628 48302 33630 48354
rect 33682 48302 33684 48354
rect 33628 48290 33684 48302
rect 33740 47908 33796 49196
rect 33852 48804 33908 49756
rect 33964 49746 34020 49756
rect 34188 49476 34244 50428
rect 35196 50484 35252 50494
rect 35196 50482 35364 50484
rect 35196 50430 35198 50482
rect 35250 50430 35364 50482
rect 35196 50428 35364 50430
rect 35196 50418 35252 50428
rect 33852 48738 33908 48748
rect 33964 49420 34244 49476
rect 34300 50370 34356 50382
rect 34748 50372 34804 50382
rect 34300 50318 34302 50370
rect 34354 50318 34356 50370
rect 33292 47058 33348 47068
rect 33628 47852 33796 47908
rect 33852 48242 33908 48254
rect 33852 48190 33854 48242
rect 33906 48190 33908 48242
rect 33628 46898 33684 47852
rect 33628 46846 33630 46898
rect 33682 46846 33684 46898
rect 33628 46834 33684 46846
rect 33852 46452 33908 48190
rect 33964 46676 34020 49420
rect 34300 48468 34356 50318
rect 34300 48402 34356 48412
rect 34412 50370 34804 50372
rect 34412 50318 34750 50370
rect 34802 50318 34804 50370
rect 34412 50316 34804 50318
rect 34412 49026 34468 50316
rect 34748 50306 34804 50316
rect 34412 48974 34414 49026
rect 34466 48974 34468 49026
rect 34412 48356 34468 48974
rect 34076 48244 34132 48254
rect 34132 48188 34244 48244
rect 34076 48150 34132 48188
rect 34076 47460 34132 47470
rect 34076 47366 34132 47404
rect 33964 46620 34132 46676
rect 33964 46452 34020 46462
rect 33404 46450 34020 46452
rect 33404 46398 33966 46450
rect 34018 46398 34020 46450
rect 33404 46396 34020 46398
rect 33404 46002 33460 46396
rect 33964 46386 34020 46396
rect 33964 46228 34020 46238
rect 33404 45950 33406 46002
rect 33458 45950 33460 46002
rect 33404 45938 33460 45950
rect 33516 46116 33572 46126
rect 33516 45890 33572 46060
rect 33516 45838 33518 45890
rect 33570 45838 33572 45890
rect 33516 45826 33572 45838
rect 33740 46004 33796 46014
rect 31948 42756 32004 42766
rect 31948 42662 32004 42700
rect 32844 42194 32900 43036
rect 32844 42142 32846 42194
rect 32898 42142 32900 42194
rect 32844 42130 32900 42142
rect 33068 42756 33124 42766
rect 33180 42756 33236 43932
rect 33292 45668 33348 45678
rect 33292 42980 33348 45612
rect 33628 44996 33684 45006
rect 33628 44902 33684 44940
rect 33292 42914 33348 42924
rect 33404 44322 33460 44334
rect 33404 44270 33406 44322
rect 33458 44270 33460 44322
rect 33068 42754 33236 42756
rect 33068 42702 33070 42754
rect 33122 42702 33236 42754
rect 33068 42700 33236 42702
rect 33292 42756 33348 42766
rect 33404 42756 33460 44270
rect 33292 42754 33460 42756
rect 33292 42702 33294 42754
rect 33346 42702 33460 42754
rect 33292 42700 33460 42702
rect 33516 43428 33572 43438
rect 31724 41860 31780 41870
rect 31724 41766 31780 41804
rect 32284 41858 32340 41870
rect 32284 41806 32286 41858
rect 32338 41806 32340 41858
rect 32284 41748 32340 41806
rect 32284 41682 32340 41692
rect 32508 41860 32564 41870
rect 32508 41746 32564 41804
rect 32508 41694 32510 41746
rect 32562 41694 32564 41746
rect 32284 41188 32340 41198
rect 32508 41188 32564 41694
rect 32284 41186 32564 41188
rect 32284 41134 32286 41186
rect 32338 41134 32564 41186
rect 32284 41132 32564 41134
rect 32284 40852 32340 41132
rect 32284 40786 32340 40796
rect 32844 40962 32900 40974
rect 32844 40910 32846 40962
rect 32898 40910 32900 40962
rect 32284 40628 32340 40638
rect 32340 40572 32676 40628
rect 32284 40496 32340 40572
rect 32396 40404 32452 40414
rect 31724 40292 31780 40302
rect 31724 40198 31780 40236
rect 31836 39956 31892 39966
rect 31724 39618 31780 39630
rect 31724 39566 31726 39618
rect 31778 39566 31780 39618
rect 31724 39396 31780 39566
rect 31724 39330 31780 39340
rect 31500 36594 31556 36606
rect 31500 36542 31502 36594
rect 31554 36542 31556 36594
rect 31500 35700 31556 36542
rect 31612 36370 31668 37772
rect 31724 38834 31780 38846
rect 31724 38782 31726 38834
rect 31778 38782 31780 38834
rect 31724 37492 31780 38782
rect 31836 38724 31892 39900
rect 32172 39620 32228 39630
rect 32172 39526 32228 39564
rect 31836 38162 31892 38668
rect 31836 38110 31838 38162
rect 31890 38110 31892 38162
rect 31836 38098 31892 38110
rect 31724 37266 31780 37436
rect 32060 37940 32116 37950
rect 32060 37490 32116 37884
rect 32060 37438 32062 37490
rect 32114 37438 32116 37490
rect 32060 37426 32116 37438
rect 32396 37492 32452 40348
rect 32620 38724 32676 40572
rect 32844 40402 32900 40910
rect 32844 40350 32846 40402
rect 32898 40350 32900 40402
rect 32844 40292 32900 40350
rect 33068 40404 33124 42700
rect 33068 40338 33124 40348
rect 32844 40226 32900 40236
rect 33292 39396 33348 42700
rect 33516 41748 33572 43372
rect 33516 41074 33572 41692
rect 33516 41022 33518 41074
rect 33570 41022 33572 41074
rect 33292 39330 33348 39340
rect 33404 40852 33460 40862
rect 32620 38722 32788 38724
rect 32620 38670 32622 38722
rect 32674 38670 32788 38722
rect 32620 38668 32788 38670
rect 32620 38658 32676 38668
rect 32620 37828 32676 37838
rect 32620 37734 32676 37772
rect 32396 37426 32452 37436
rect 31724 37214 31726 37266
rect 31778 37214 31780 37266
rect 31724 37202 31780 37214
rect 32172 37154 32228 37166
rect 32172 37102 32174 37154
rect 32226 37102 32228 37154
rect 31836 37044 31892 37054
rect 31836 36484 31892 36988
rect 32172 37044 32228 37102
rect 32172 36978 32228 36988
rect 32732 37044 32788 38668
rect 33404 38668 33460 40796
rect 33516 40628 33572 41022
rect 33628 41186 33684 41198
rect 33628 41134 33630 41186
rect 33682 41134 33684 41186
rect 33628 40964 33684 41134
rect 33628 40898 33684 40908
rect 33516 40562 33572 40572
rect 33516 40402 33572 40414
rect 33516 40350 33518 40402
rect 33570 40350 33572 40402
rect 33516 40292 33572 40350
rect 33516 38948 33572 40236
rect 33740 39172 33796 45948
rect 33964 45780 34020 46172
rect 34076 46004 34132 46620
rect 34188 46674 34244 48188
rect 34412 47460 34468 48300
rect 34524 49810 34580 49822
rect 34524 49758 34526 49810
rect 34578 49758 34580 49810
rect 34524 48692 34580 49758
rect 35308 49812 35364 50428
rect 35308 49746 35364 49756
rect 35980 50260 36036 50270
rect 34636 49700 34692 49710
rect 34636 49606 34692 49644
rect 35532 49698 35588 49710
rect 35532 49646 35534 49698
rect 35586 49646 35588 49698
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 34524 47682 34580 48636
rect 34524 47630 34526 47682
rect 34578 47630 34580 47682
rect 34524 47618 34580 47630
rect 34860 49026 34916 49038
rect 34860 48974 34862 49026
rect 34914 48974 34916 49026
rect 34412 47394 34468 47404
rect 34524 47458 34580 47470
rect 34524 47406 34526 47458
rect 34578 47406 34580 47458
rect 34412 47236 34468 47246
rect 34188 46622 34190 46674
rect 34242 46622 34244 46674
rect 34188 46610 34244 46622
rect 34300 47124 34356 47134
rect 34300 46900 34356 47068
rect 34188 46004 34244 46014
rect 34076 46002 34244 46004
rect 34076 45950 34190 46002
rect 34242 45950 34244 46002
rect 34076 45948 34244 45950
rect 34188 45938 34244 45948
rect 34300 45890 34356 46844
rect 34300 45838 34302 45890
rect 34354 45838 34356 45890
rect 34300 45826 34356 45838
rect 34076 45780 34132 45790
rect 33964 45778 34132 45780
rect 33964 45726 34078 45778
rect 34130 45726 34132 45778
rect 33964 45724 34132 45726
rect 34076 45714 34132 45724
rect 34412 44772 34468 47180
rect 34524 46004 34580 47406
rect 34524 45938 34580 45948
rect 34748 47124 34804 47134
rect 34748 45890 34804 47068
rect 34748 45838 34750 45890
rect 34802 45838 34804 45890
rect 34748 45826 34804 45838
rect 34860 45556 34916 48974
rect 35532 49028 35588 49646
rect 35756 49700 35812 49710
rect 35756 49138 35812 49644
rect 35756 49086 35758 49138
rect 35810 49086 35812 49138
rect 35756 49074 35812 49086
rect 35532 48962 35588 48972
rect 35980 48804 36036 50204
rect 36092 50036 36148 50046
rect 36204 50036 36260 51326
rect 36316 51380 36372 51390
rect 36316 50594 36372 51324
rect 36540 51378 36596 51390
rect 36540 51326 36542 51378
rect 36594 51326 36596 51378
rect 36428 51044 36484 51054
rect 36540 51044 36596 51326
rect 36876 51378 36932 51390
rect 36876 51326 36878 51378
rect 36930 51326 36932 51378
rect 36540 50988 36820 51044
rect 36428 50706 36484 50988
rect 36428 50654 36430 50706
rect 36482 50654 36484 50706
rect 36428 50642 36484 50654
rect 36316 50542 36318 50594
rect 36370 50542 36372 50594
rect 36316 50428 36372 50542
rect 36764 50596 36820 50988
rect 36764 50502 36820 50540
rect 36876 50708 36932 51326
rect 36876 50428 36932 50652
rect 36316 50372 36484 50428
rect 36092 50034 36260 50036
rect 36092 49982 36094 50034
rect 36146 49982 36260 50034
rect 36092 49980 36260 49982
rect 36092 49970 36148 49980
rect 36092 49028 36148 49038
rect 36148 48972 36260 49028
rect 36092 48896 36148 48972
rect 35868 48748 36036 48804
rect 35644 48692 35700 48702
rect 35644 48130 35700 48636
rect 35644 48078 35646 48130
rect 35698 48078 35700 48130
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 35644 47012 35700 48078
rect 35868 48020 35924 48748
rect 35980 48244 36036 48254
rect 35980 48242 36148 48244
rect 35980 48190 35982 48242
rect 36034 48190 36148 48242
rect 35980 48188 36148 48190
rect 35980 48178 36036 48188
rect 35868 47964 36036 48020
rect 35644 46946 35700 46956
rect 35756 46676 35812 46686
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 35644 46004 35700 46014
rect 35756 46004 35812 46620
rect 35644 46002 35812 46004
rect 35644 45950 35646 46002
rect 35698 45950 35812 46002
rect 35644 45948 35812 45950
rect 35868 46564 35924 46574
rect 35980 46564 36036 47964
rect 36092 47460 36148 48188
rect 36204 47682 36260 48972
rect 36428 48468 36484 50372
rect 36652 50372 36932 50428
rect 36540 49700 36596 49710
rect 36540 49606 36596 49644
rect 36540 49140 36596 49150
rect 36652 49140 36708 50372
rect 36540 49138 36708 49140
rect 36540 49086 36542 49138
rect 36594 49086 36708 49138
rect 36540 49084 36708 49086
rect 36764 49700 36820 49710
rect 36540 49074 36596 49084
rect 36428 48412 36708 48468
rect 36428 48244 36484 48254
rect 36428 48150 36484 48188
rect 36204 47630 36206 47682
rect 36258 47630 36260 47682
rect 36204 47618 36260 47630
rect 36204 47460 36260 47470
rect 36092 47458 36260 47460
rect 36092 47406 36206 47458
rect 36258 47406 36260 47458
rect 36092 47404 36260 47406
rect 36204 46786 36260 47404
rect 36540 47346 36596 47358
rect 36540 47294 36542 47346
rect 36594 47294 36596 47346
rect 36540 47012 36596 47294
rect 36540 46946 36596 46956
rect 36652 46898 36708 48412
rect 36652 46846 36654 46898
rect 36706 46846 36708 46898
rect 36652 46834 36708 46846
rect 36204 46734 36206 46786
rect 36258 46734 36260 46786
rect 36204 46722 36260 46734
rect 35980 46508 36372 46564
rect 35644 45938 35700 45948
rect 35756 45778 35812 45790
rect 35756 45726 35758 45778
rect 35810 45726 35812 45778
rect 35532 45668 35588 45678
rect 35532 45574 35588 45612
rect 35756 45668 35812 45726
rect 35756 45602 35812 45612
rect 34860 45490 34916 45500
rect 34748 45444 34804 45454
rect 34636 45332 34692 45342
rect 34412 44706 34468 44716
rect 34524 45106 34580 45118
rect 34524 45054 34526 45106
rect 34578 45054 34580 45106
rect 34524 43650 34580 45054
rect 34636 43708 34692 45276
rect 34748 45330 34804 45388
rect 34748 45278 34750 45330
rect 34802 45278 34804 45330
rect 34748 45266 34804 45278
rect 34860 45106 34916 45118
rect 34860 45054 34862 45106
rect 34914 45054 34916 45106
rect 34860 44996 34916 45054
rect 35084 45108 35140 45118
rect 35084 45014 35140 45052
rect 35532 45108 35588 45118
rect 34748 44322 34804 44334
rect 34748 44270 34750 44322
rect 34802 44270 34804 44322
rect 34748 44212 34804 44270
rect 34748 44146 34804 44156
rect 34860 44100 34916 44940
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 34860 44034 34916 44044
rect 35308 44322 35364 44334
rect 35308 44270 35310 44322
rect 35362 44270 35364 44322
rect 34636 43652 34916 43708
rect 34524 43598 34526 43650
rect 34578 43598 34580 43650
rect 34076 43540 34132 43550
rect 33852 43204 33908 43214
rect 33852 41970 33908 43148
rect 33852 41918 33854 41970
rect 33906 41918 33908 41970
rect 33852 41906 33908 41918
rect 34076 41970 34132 43484
rect 34300 43538 34356 43550
rect 34300 43486 34302 43538
rect 34354 43486 34356 43538
rect 34076 41918 34078 41970
rect 34130 41918 34132 41970
rect 34076 41906 34132 41918
rect 34188 43316 34244 43326
rect 34188 42308 34244 43260
rect 34188 41412 34244 42252
rect 34300 41636 34356 43486
rect 34300 41570 34356 41580
rect 34412 42754 34468 42766
rect 34412 42702 34414 42754
rect 34466 42702 34468 42754
rect 34412 42084 34468 42702
rect 34188 41410 34356 41412
rect 34188 41358 34190 41410
rect 34242 41358 34356 41410
rect 34188 41356 34356 41358
rect 34188 41346 34244 41356
rect 34300 40402 34356 41356
rect 34300 40350 34302 40402
rect 34354 40350 34356 40402
rect 34188 40292 34244 40302
rect 33852 39172 33908 39182
rect 33740 39116 33852 39172
rect 33628 38948 33684 38958
rect 33516 38892 33628 38948
rect 33628 38854 33684 38892
rect 33852 38946 33908 39116
rect 34076 39060 34132 39070
rect 34076 38966 34132 39004
rect 33852 38894 33854 38946
rect 33906 38894 33908 38946
rect 33852 38882 33908 38894
rect 34188 38834 34244 40236
rect 34300 40180 34356 40350
rect 34300 40114 34356 40124
rect 34412 39730 34468 42028
rect 34524 41972 34580 43598
rect 34524 41746 34580 41916
rect 34524 41694 34526 41746
rect 34578 41694 34580 41746
rect 34524 41682 34580 41694
rect 34524 41412 34580 41422
rect 34524 41318 34580 41356
rect 34412 39678 34414 39730
rect 34466 39678 34468 39730
rect 34412 39666 34468 39678
rect 34524 40402 34580 40414
rect 34524 40350 34526 40402
rect 34578 40350 34580 40402
rect 34524 39620 34580 40350
rect 34524 39554 34580 39564
rect 34636 40402 34692 40414
rect 34636 40350 34638 40402
rect 34690 40350 34692 40402
rect 34636 39508 34692 40350
rect 34748 40404 34804 40414
rect 34748 39842 34804 40348
rect 34748 39790 34750 39842
rect 34802 39790 34804 39842
rect 34748 39778 34804 39790
rect 34860 39620 34916 43652
rect 35308 43652 35364 44270
rect 35420 43764 35476 43774
rect 35532 43764 35588 45052
rect 35756 45108 35812 45118
rect 35756 45014 35812 45052
rect 35420 43762 35588 43764
rect 35420 43710 35422 43762
rect 35474 43710 35588 43762
rect 35420 43708 35588 43710
rect 35756 44212 35812 44222
rect 35420 43698 35476 43708
rect 35084 43540 35140 43550
rect 35084 43446 35140 43484
rect 35308 43316 35364 43596
rect 35084 43260 35364 43316
rect 35084 42756 35140 43260
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 35756 42866 35812 44156
rect 35756 42814 35758 42866
rect 35810 42814 35812 42866
rect 35756 42802 35812 42814
rect 35308 42756 35364 42766
rect 34972 42754 35364 42756
rect 34972 42702 35310 42754
rect 35362 42702 35364 42754
rect 34972 42700 35364 42702
rect 34972 39956 35028 42700
rect 35308 42690 35364 42700
rect 35868 42644 35924 46508
rect 36092 46004 36148 46014
rect 35980 45106 36036 45118
rect 35980 45054 35982 45106
rect 36034 45054 36036 45106
rect 35980 44996 36036 45054
rect 35980 44930 36036 44940
rect 36092 44546 36148 45948
rect 36204 45892 36260 45902
rect 36204 45798 36260 45836
rect 36092 44494 36094 44546
rect 36146 44494 36148 44546
rect 36092 44482 36148 44494
rect 35980 44434 36036 44446
rect 35980 44382 35982 44434
rect 36034 44382 36036 44434
rect 35980 43708 36036 44382
rect 36316 44100 36372 46508
rect 36764 46452 36820 49644
rect 37100 49698 37156 49710
rect 37100 49646 37102 49698
rect 37154 49646 37156 49698
rect 37100 48692 37156 49646
rect 37100 48626 37156 48636
rect 36988 48132 37044 48142
rect 36988 48130 37156 48132
rect 36988 48078 36990 48130
rect 37042 48078 37156 48130
rect 36988 48076 37156 48078
rect 36988 48066 37044 48076
rect 36988 47348 37044 47358
rect 36876 46786 36932 46798
rect 36876 46734 36878 46786
rect 36930 46734 36932 46786
rect 36876 46676 36932 46734
rect 36876 46610 36932 46620
rect 36988 46674 37044 47292
rect 36988 46622 36990 46674
rect 37042 46622 37044 46674
rect 36988 46564 37044 46622
rect 36988 46498 37044 46508
rect 36764 46396 36932 46452
rect 36540 46116 36596 46126
rect 36540 45668 36596 46060
rect 36764 45892 36820 45902
rect 36652 45668 36708 45678
rect 36540 45666 36708 45668
rect 36540 45614 36654 45666
rect 36706 45614 36708 45666
rect 36540 45612 36708 45614
rect 36540 44996 36596 45612
rect 36652 45602 36708 45612
rect 36652 45220 36708 45230
rect 36652 45126 36708 45164
rect 36540 44940 36708 44996
rect 36316 44034 36372 44044
rect 35980 43652 36148 43708
rect 35980 43540 36036 43550
rect 35980 43446 36036 43484
rect 35756 42588 35924 42644
rect 35532 42420 35588 42430
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35196 40964 35252 40974
rect 35196 40870 35252 40908
rect 35532 40516 35588 42364
rect 35644 41858 35700 41870
rect 35644 41806 35646 41858
rect 35698 41806 35700 41858
rect 35644 41412 35700 41806
rect 35644 41346 35700 41356
rect 35532 40450 35588 40460
rect 35644 40290 35700 40302
rect 35644 40238 35646 40290
rect 35698 40238 35700 40290
rect 35084 40180 35140 40190
rect 35084 40178 35588 40180
rect 35084 40126 35086 40178
rect 35138 40126 35588 40178
rect 35084 40124 35588 40126
rect 35084 40114 35140 40124
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 34972 39900 35140 39956
rect 35196 39946 35460 39956
rect 34188 38782 34190 38834
rect 34242 38782 34244 38834
rect 34188 38724 34244 38782
rect 33404 38612 33572 38668
rect 34188 38658 34244 38668
rect 34524 39172 34580 39182
rect 34524 38668 34580 39116
rect 34636 39060 34692 39452
rect 34636 38994 34692 39004
rect 34748 39564 34916 39620
rect 34972 39620 35028 39630
rect 34524 38612 34692 38668
rect 33404 38276 33460 38286
rect 33068 37940 33124 37950
rect 32172 36708 32228 36718
rect 31948 36596 32004 36606
rect 31948 36502 32004 36540
rect 31612 36318 31614 36370
rect 31666 36318 31668 36370
rect 31612 36306 31668 36318
rect 31724 36482 31892 36484
rect 31724 36430 31838 36482
rect 31890 36430 31892 36482
rect 31724 36428 31892 36430
rect 31612 35700 31668 35710
rect 31500 35698 31668 35700
rect 31500 35646 31614 35698
rect 31666 35646 31668 35698
rect 31500 35644 31668 35646
rect 31612 35252 31668 35644
rect 31612 35186 31668 35196
rect 31500 34916 31556 34926
rect 31500 33908 31556 34860
rect 31724 34804 31780 36428
rect 31836 36418 31892 36428
rect 32060 36372 32116 36382
rect 32060 36278 32116 36316
rect 31836 35700 31892 35710
rect 31836 35606 31892 35644
rect 32172 35698 32228 36652
rect 32172 35646 32174 35698
rect 32226 35646 32228 35698
rect 32172 35634 32228 35646
rect 32396 36260 32452 36270
rect 32396 35812 32452 36204
rect 32620 36260 32676 36270
rect 32620 36166 32676 36204
rect 31948 35586 32004 35598
rect 31948 35534 31950 35586
rect 32002 35534 32004 35586
rect 31948 34916 32004 35534
rect 32396 35028 32452 35756
rect 32620 35924 32676 35934
rect 32172 34916 32228 34926
rect 31948 34914 32228 34916
rect 31948 34862 32174 34914
rect 32226 34862 32228 34914
rect 31948 34860 32228 34862
rect 32172 34850 32228 34860
rect 32396 34914 32452 34972
rect 32396 34862 32398 34914
rect 32450 34862 32452 34914
rect 32396 34850 32452 34862
rect 32508 35586 32564 35598
rect 32508 35534 32510 35586
rect 32562 35534 32564 35586
rect 32508 34804 32564 35534
rect 31724 34748 32116 34804
rect 31612 34692 31668 34702
rect 31612 34690 32004 34692
rect 31612 34638 31614 34690
rect 31666 34638 32004 34690
rect 31612 34636 32004 34638
rect 31612 34626 31668 34636
rect 31724 34132 31780 34142
rect 31724 34038 31780 34076
rect 31948 34130 32004 34636
rect 32060 34580 32116 34748
rect 32060 34514 32116 34524
rect 32284 34690 32340 34702
rect 32284 34638 32286 34690
rect 32338 34638 32340 34690
rect 31948 34078 31950 34130
rect 32002 34078 32004 34130
rect 31948 34066 32004 34078
rect 32060 34018 32116 34030
rect 32060 33966 32062 34018
rect 32114 33966 32116 34018
rect 31500 33852 31780 33908
rect 31388 33516 31668 33572
rect 31164 33348 31220 33358
rect 31164 33346 31556 33348
rect 31164 33294 31166 33346
rect 31218 33294 31556 33346
rect 31164 33292 31556 33294
rect 31164 33282 31220 33292
rect 30884 31612 30996 31668
rect 31276 33124 31332 33134
rect 30492 31490 30548 31500
rect 30716 31556 30772 31566
rect 30828 31556 30884 31612
rect 30716 31554 30884 31556
rect 30716 31502 30718 31554
rect 30770 31502 30884 31554
rect 30716 31500 30884 31502
rect 30716 31490 30772 31500
rect 30380 30482 30436 30492
rect 30492 30882 30548 30894
rect 30492 30830 30494 30882
rect 30546 30830 30548 30882
rect 30268 29138 30324 29148
rect 30380 30210 30436 30222
rect 30380 30158 30382 30210
rect 30434 30158 30436 30210
rect 30380 29538 30436 30158
rect 30380 29486 30382 29538
rect 30434 29486 30436 29538
rect 30156 28642 30324 28644
rect 30156 28590 30158 28642
rect 30210 28590 30324 28642
rect 30156 28588 30324 28590
rect 30156 28578 30212 28588
rect 30156 28420 30212 28430
rect 30156 28326 30212 28364
rect 30268 27970 30324 28588
rect 30268 27918 30270 27970
rect 30322 27918 30324 27970
rect 30268 27906 30324 27918
rect 29932 27186 30100 27188
rect 29932 27134 29934 27186
rect 29986 27134 30100 27186
rect 29932 27132 30100 27134
rect 30268 27748 30324 27758
rect 29932 27122 29988 27132
rect 29708 25788 29876 25844
rect 30044 26402 30100 26414
rect 30044 26350 30046 26402
rect 30098 26350 30100 26402
rect 29708 25060 29764 25788
rect 29820 25282 29876 25294
rect 29820 25230 29822 25282
rect 29874 25230 29876 25282
rect 29820 25172 29876 25230
rect 29820 25106 29876 25116
rect 29596 25004 29764 25060
rect 29484 24836 29540 24846
rect 29484 24742 29540 24780
rect 29596 24164 29652 25004
rect 29932 24836 29988 24846
rect 29372 21586 29428 22092
rect 29372 21534 29374 21586
rect 29426 21534 29428 21586
rect 29036 20850 29092 20860
rect 29260 21474 29316 21486
rect 29260 21422 29262 21474
rect 29314 21422 29316 21474
rect 29260 20804 29316 21422
rect 29260 20738 29316 20748
rect 28812 20692 28868 20702
rect 28812 20690 29204 20692
rect 28812 20638 28814 20690
rect 28866 20638 29204 20690
rect 28812 20636 29204 20638
rect 28812 20626 28868 20636
rect 28924 20244 28980 20254
rect 28700 20188 28924 20244
rect 28532 20076 28644 20132
rect 28476 20066 28532 20076
rect 28252 19346 28420 19348
rect 28252 19294 28366 19346
rect 28418 19294 28420 19346
rect 28252 19292 28420 19294
rect 28028 19068 28196 19124
rect 27916 19010 28084 19012
rect 27916 18958 27918 19010
rect 27970 18958 28084 19010
rect 27916 18956 28084 18958
rect 27916 18946 27972 18956
rect 27804 18622 27806 18674
rect 27858 18622 27860 18674
rect 27804 18610 27860 18622
rect 27916 18676 27972 18686
rect 27916 18562 27972 18620
rect 27916 18510 27918 18562
rect 27970 18510 27972 18562
rect 27916 18498 27972 18510
rect 27692 18172 27972 18228
rect 27580 17890 27636 17902
rect 27580 17838 27582 17890
rect 27634 17838 27636 17890
rect 27580 17778 27636 17838
rect 27580 17726 27582 17778
rect 27634 17726 27636 17778
rect 27580 17714 27636 17726
rect 27356 16940 27524 16996
rect 27132 15250 27188 15260
rect 27244 16882 27300 16894
rect 27244 16830 27246 16882
rect 27298 16830 27300 16882
rect 27244 15148 27300 16830
rect 27356 16660 27412 16940
rect 27356 15986 27412 16604
rect 27468 16770 27524 16782
rect 27468 16718 27470 16770
rect 27522 16718 27524 16770
rect 27468 16210 27524 16718
rect 27468 16158 27470 16210
rect 27522 16158 27524 16210
rect 27468 16146 27524 16158
rect 27580 16324 27636 16334
rect 27804 16324 27860 16334
rect 27580 16322 27860 16324
rect 27580 16270 27582 16322
rect 27634 16270 27806 16322
rect 27858 16270 27860 16322
rect 27580 16268 27860 16270
rect 27356 15934 27358 15986
rect 27410 15934 27412 15986
rect 27356 15652 27412 15934
rect 27356 15586 27412 15596
rect 27468 15314 27524 15326
rect 27468 15262 27470 15314
rect 27522 15262 27524 15314
rect 27468 15148 27524 15262
rect 26572 15092 26852 15148
rect 27244 15092 27524 15148
rect 27580 15148 27636 16268
rect 27804 16258 27860 16268
rect 27580 15092 27860 15148
rect 26572 14644 26628 14654
rect 26348 14642 26628 14644
rect 26348 14590 26574 14642
rect 26626 14590 26628 14642
rect 26348 14588 26628 14590
rect 26572 14578 26628 14588
rect 26460 14308 26516 14318
rect 26348 14306 26516 14308
rect 26348 14254 26462 14306
rect 26514 14254 26516 14306
rect 26348 14252 26516 14254
rect 26348 13748 26404 14252
rect 26460 14242 26516 14252
rect 26684 14306 26740 14318
rect 26684 14254 26686 14306
rect 26738 14254 26740 14306
rect 26348 13682 26404 13692
rect 26460 13860 26516 13870
rect 26460 13636 26516 13804
rect 26460 13634 26628 13636
rect 26460 13582 26462 13634
rect 26514 13582 26628 13634
rect 26460 13580 26628 13582
rect 26460 13570 26516 13580
rect 26348 13524 26404 13534
rect 26348 12850 26404 13468
rect 26572 13186 26628 13580
rect 26572 13134 26574 13186
rect 26626 13134 26628 13186
rect 26460 13076 26516 13086
rect 26460 12982 26516 13020
rect 26348 12798 26350 12850
rect 26402 12798 26404 12850
rect 26348 12786 26404 12798
rect 26236 12460 26404 12516
rect 26012 12402 26180 12404
rect 26012 12350 26014 12402
rect 26066 12350 26180 12402
rect 26012 12348 26180 12350
rect 26012 12338 26068 12348
rect 26124 11396 26180 11406
rect 25900 11282 25956 11294
rect 25900 11230 25902 11282
rect 25954 11230 25956 11282
rect 25900 11172 25956 11230
rect 25564 10782 25566 10834
rect 25618 10782 25620 10834
rect 25564 10770 25620 10782
rect 25676 11116 25900 11172
rect 25676 10834 25732 11116
rect 25900 11106 25956 11116
rect 26012 11282 26068 11294
rect 26012 11230 26014 11282
rect 26066 11230 26068 11282
rect 26012 11060 26068 11230
rect 26124 11284 26180 11340
rect 26124 11282 26292 11284
rect 26124 11230 26126 11282
rect 26178 11230 26292 11282
rect 26124 11228 26292 11230
rect 26124 11218 26180 11228
rect 26012 10994 26068 11004
rect 25676 10782 25678 10834
rect 25730 10782 25732 10834
rect 25676 10770 25732 10782
rect 25900 10836 25956 10846
rect 25788 9828 25844 9838
rect 25788 9734 25844 9772
rect 25676 9268 25732 9278
rect 25676 9174 25732 9212
rect 25900 8428 25956 10780
rect 26124 10724 26180 10734
rect 26124 10388 26180 10668
rect 26236 10500 26292 11228
rect 26348 11060 26404 12460
rect 26348 10994 26404 11004
rect 26460 12066 26516 12078
rect 26460 12014 26462 12066
rect 26514 12014 26516 12066
rect 26460 10836 26516 12014
rect 26572 11618 26628 13134
rect 26684 13188 26740 14254
rect 26796 14308 26852 15092
rect 27468 15026 27524 15036
rect 27692 14756 27748 14766
rect 27132 14754 27748 14756
rect 27132 14702 27694 14754
rect 27746 14702 27748 14754
rect 27132 14700 27748 14702
rect 27132 14530 27188 14700
rect 27692 14690 27748 14700
rect 27132 14478 27134 14530
rect 27186 14478 27188 14530
rect 27132 14466 27188 14478
rect 26796 14242 26852 14252
rect 27244 14420 27300 14430
rect 26684 13122 26740 13132
rect 27244 14196 27300 14364
rect 27580 14418 27636 14430
rect 27580 14366 27582 14418
rect 27634 14366 27636 14418
rect 27132 12738 27188 12750
rect 27132 12686 27134 12738
rect 27186 12686 27188 12738
rect 27132 11844 27188 12686
rect 27244 12402 27300 14140
rect 27244 12350 27246 12402
rect 27298 12350 27300 12402
rect 27244 12338 27300 12350
rect 27356 14308 27412 14318
rect 27132 11778 27188 11788
rect 26572 11566 26574 11618
rect 26626 11566 26628 11618
rect 26572 11554 26628 11566
rect 26460 10770 26516 10780
rect 27132 11282 27188 11294
rect 27132 11230 27134 11282
rect 27186 11230 27188 11282
rect 26796 10722 26852 10734
rect 26796 10670 26798 10722
rect 26850 10670 26852 10722
rect 26684 10500 26740 10510
rect 26236 10498 26740 10500
rect 26236 10446 26686 10498
rect 26738 10446 26740 10498
rect 26236 10444 26740 10446
rect 26684 10434 26740 10444
rect 26124 10332 26404 10388
rect 26348 10050 26404 10332
rect 26348 9998 26350 10050
rect 26402 9998 26404 10050
rect 26348 9986 26404 9998
rect 26684 10052 26740 10062
rect 26236 9268 26292 9278
rect 26684 9268 26740 9996
rect 26796 9828 26852 10670
rect 27132 10724 27188 11230
rect 27244 11172 27300 11182
rect 27244 11078 27300 11116
rect 27132 10658 27188 10668
rect 27020 10386 27076 10398
rect 27020 10334 27022 10386
rect 27074 10334 27076 10386
rect 27020 10052 27076 10334
rect 27020 9986 27076 9996
rect 27356 10050 27412 14252
rect 27580 13860 27636 14366
rect 27692 14306 27748 14318
rect 27692 14254 27694 14306
rect 27746 14254 27748 14306
rect 27692 14196 27748 14254
rect 27692 14130 27748 14140
rect 27580 13794 27636 13804
rect 27692 13748 27748 13758
rect 27692 13654 27748 13692
rect 27580 13522 27636 13534
rect 27580 13470 27582 13522
rect 27634 13470 27636 13522
rect 27468 12964 27524 12974
rect 27580 12964 27636 13470
rect 27468 12962 27636 12964
rect 27468 12910 27470 12962
rect 27522 12910 27636 12962
rect 27468 12908 27636 12910
rect 27468 12898 27524 12908
rect 27580 12068 27636 12078
rect 27580 11974 27636 12012
rect 27804 11844 27860 15092
rect 27916 14756 27972 18172
rect 28028 17890 28084 18956
rect 28028 17838 28030 17890
rect 28082 17838 28084 17890
rect 28028 17826 28084 17838
rect 28140 17668 28196 19068
rect 28028 17612 28196 17668
rect 28028 15538 28084 17612
rect 28140 17444 28196 17454
rect 28140 17350 28196 17388
rect 28252 16210 28308 19292
rect 28364 19282 28420 19292
rect 28476 18788 28532 18798
rect 28364 18452 28420 18462
rect 28364 18358 28420 18396
rect 28476 17444 28532 18732
rect 28476 17378 28532 17388
rect 28588 17778 28644 20076
rect 28700 20020 28756 20030
rect 28700 19926 28756 19964
rect 28924 20018 28980 20188
rect 28924 19966 28926 20018
rect 28978 19966 28980 20018
rect 28812 19348 28868 19358
rect 28812 19254 28868 19292
rect 28812 18338 28868 18350
rect 28812 18286 28814 18338
rect 28866 18286 28868 18338
rect 28812 18228 28868 18286
rect 28812 18162 28868 18172
rect 28588 17726 28590 17778
rect 28642 17726 28644 17778
rect 28364 17108 28420 17118
rect 28364 17014 28420 17052
rect 28364 16658 28420 16670
rect 28364 16606 28366 16658
rect 28418 16606 28420 16658
rect 28364 16322 28420 16606
rect 28476 16660 28532 16670
rect 28588 16660 28644 17726
rect 28700 17442 28756 17454
rect 28700 17390 28702 17442
rect 28754 17390 28756 17442
rect 28700 17332 28756 17390
rect 28700 16882 28756 17276
rect 28700 16830 28702 16882
rect 28754 16830 28756 16882
rect 28700 16818 28756 16830
rect 28588 16604 28756 16660
rect 28476 16566 28532 16604
rect 28364 16270 28366 16322
rect 28418 16270 28420 16322
rect 28364 16258 28420 16270
rect 28252 16158 28254 16210
rect 28306 16158 28308 16210
rect 28252 16146 28308 16158
rect 28028 15486 28030 15538
rect 28082 15486 28084 15538
rect 28028 15474 28084 15486
rect 28476 15876 28532 15886
rect 28476 15538 28532 15820
rect 28588 15874 28644 15886
rect 28588 15822 28590 15874
rect 28642 15822 28644 15874
rect 28588 15764 28644 15822
rect 28588 15698 28644 15708
rect 28476 15486 28478 15538
rect 28530 15486 28532 15538
rect 28476 15474 28532 15486
rect 28588 15316 28644 15326
rect 28476 15260 28588 15316
rect 28476 15148 28532 15260
rect 28588 15250 28644 15260
rect 28700 15148 28756 16604
rect 27916 12404 27972 14700
rect 28364 15092 28532 15148
rect 28588 15092 28756 15148
rect 28812 16436 28868 16446
rect 28812 15764 28868 16380
rect 28364 14306 28420 15092
rect 28364 14254 28366 14306
rect 28418 14254 28420 14306
rect 28028 13524 28084 13534
rect 28028 13074 28084 13468
rect 28028 13022 28030 13074
rect 28082 13022 28084 13074
rect 28028 13010 28084 13022
rect 28364 12740 28420 14254
rect 28588 13970 28644 15036
rect 28812 14306 28868 15708
rect 28924 15876 28980 19966
rect 29036 18452 29092 18462
rect 29036 16884 29092 18396
rect 29148 18340 29204 20636
rect 29260 19796 29316 19806
rect 29260 19702 29316 19740
rect 29372 19012 29428 21534
rect 29484 24108 29652 24164
rect 29708 24780 29932 24836
rect 29484 21810 29540 24108
rect 29596 23940 29652 23950
rect 29596 23846 29652 23884
rect 29708 22482 29764 24780
rect 29932 24742 29988 24780
rect 29708 22430 29710 22482
rect 29762 22430 29764 22482
rect 29708 22418 29764 22430
rect 29484 21758 29486 21810
rect 29538 21758 29540 21810
rect 29484 19348 29540 21758
rect 30044 21364 30100 26350
rect 30156 26292 30212 26302
rect 30156 23716 30212 26236
rect 30268 26066 30324 27692
rect 30380 27188 30436 29486
rect 30492 28532 30548 30830
rect 30716 30772 30772 30782
rect 30604 30770 30772 30772
rect 30604 30718 30718 30770
rect 30770 30718 30772 30770
rect 30604 30716 30772 30718
rect 30604 29540 30660 30716
rect 30716 30706 30772 30716
rect 30828 30212 30884 31500
rect 31164 31556 31220 31566
rect 31164 31462 31220 31500
rect 30828 30146 30884 30156
rect 30940 30996 30996 31006
rect 30604 29474 30660 29484
rect 30716 30098 30772 30110
rect 30716 30046 30718 30098
rect 30770 30046 30772 30098
rect 30492 28466 30548 28476
rect 30604 29204 30660 29214
rect 30380 27122 30436 27132
rect 30492 28308 30548 28318
rect 30268 26014 30270 26066
rect 30322 26014 30324 26066
rect 30268 25508 30324 26014
rect 30380 26066 30436 26078
rect 30380 26014 30382 26066
rect 30434 26014 30436 26066
rect 30380 25956 30436 26014
rect 30380 25890 30436 25900
rect 30268 25442 30324 25452
rect 30380 25396 30436 25406
rect 30380 25302 30436 25340
rect 30380 24948 30436 24958
rect 30492 24948 30548 28252
rect 30604 27748 30660 29148
rect 30604 27682 30660 27692
rect 30716 27300 30772 30046
rect 30828 29426 30884 29438
rect 30828 29374 30830 29426
rect 30882 29374 30884 29426
rect 30828 29316 30884 29374
rect 30828 28644 30884 29260
rect 30828 28578 30884 28588
rect 30940 28530 30996 30940
rect 31052 30772 31108 30782
rect 31052 30678 31108 30716
rect 31164 29428 31220 29438
rect 31276 29428 31332 33068
rect 31500 32786 31556 33292
rect 31500 32734 31502 32786
rect 31554 32734 31556 32786
rect 31500 32722 31556 32734
rect 31388 32676 31444 32686
rect 31388 31892 31444 32620
rect 31388 31826 31444 31836
rect 31612 29652 31668 33516
rect 31724 32786 31780 33852
rect 31724 32734 31726 32786
rect 31778 32734 31780 32786
rect 31724 32722 31780 32734
rect 31836 33684 31892 33694
rect 31836 32674 31892 33628
rect 31836 32622 31838 32674
rect 31890 32622 31892 32674
rect 31836 32610 31892 32622
rect 32060 33346 32116 33966
rect 32284 34020 32340 34638
rect 32508 34468 32564 34748
rect 32284 33954 32340 33964
rect 32396 34412 32564 34468
rect 32060 33294 32062 33346
rect 32114 33294 32116 33346
rect 31836 31780 31892 31790
rect 31836 31686 31892 31724
rect 31724 31668 31780 31678
rect 31724 31574 31780 31612
rect 31948 31556 32004 31566
rect 31948 31462 32004 31500
rect 32060 31332 32116 33294
rect 31724 31276 32116 31332
rect 32172 33796 32228 33806
rect 31724 30322 31780 31276
rect 31836 30996 31892 31006
rect 31836 30902 31892 30940
rect 31724 30270 31726 30322
rect 31778 30270 31780 30322
rect 31724 30258 31780 30270
rect 32060 29652 32116 29662
rect 31612 29650 32116 29652
rect 31612 29598 32062 29650
rect 32114 29598 32116 29650
rect 31612 29596 32116 29598
rect 32060 29586 32116 29596
rect 30940 28478 30942 28530
rect 30994 28478 30996 28530
rect 30940 28420 30996 28478
rect 30940 28354 30996 28364
rect 31052 29426 31332 29428
rect 31052 29374 31166 29426
rect 31218 29374 31332 29426
rect 31052 29372 31332 29374
rect 31388 29428 31444 29438
rect 30716 27234 30772 27244
rect 30380 24946 30548 24948
rect 30380 24894 30382 24946
rect 30434 24894 30548 24946
rect 30380 24892 30548 24894
rect 30828 27188 30884 27198
rect 30828 26514 30884 27132
rect 30940 27076 30996 27086
rect 30940 26982 30996 27020
rect 30828 26462 30830 26514
rect 30882 26462 30884 26514
rect 30828 24948 30884 26462
rect 31052 25172 31108 29372
rect 31164 29362 31220 29372
rect 31388 28980 31444 29372
rect 31948 29428 32004 29438
rect 31948 29334 32004 29372
rect 31388 28642 31444 28924
rect 31388 28590 31390 28642
rect 31442 28590 31444 28642
rect 31388 28578 31444 28590
rect 31612 28642 31668 28654
rect 31612 28590 31614 28642
rect 31666 28590 31668 28642
rect 31388 28084 31444 28094
rect 31164 27300 31220 27310
rect 31164 26964 31220 27244
rect 31276 26964 31332 26974
rect 31164 26962 31332 26964
rect 31164 26910 31278 26962
rect 31330 26910 31332 26962
rect 31164 26908 31332 26910
rect 31164 26066 31220 26908
rect 31276 26898 31332 26908
rect 31276 26180 31332 26190
rect 31388 26180 31444 28028
rect 31612 27076 31668 28590
rect 31612 27010 31668 27020
rect 31836 27970 31892 27982
rect 31836 27918 31838 27970
rect 31890 27918 31892 27970
rect 31836 26908 31892 27918
rect 32172 27860 32228 33740
rect 32396 33684 32452 34412
rect 32508 33908 32564 33918
rect 32508 33814 32564 33852
rect 32396 32786 32452 33628
rect 32620 33348 32676 35868
rect 32732 33796 32788 36988
rect 32844 37154 32900 37166
rect 32844 37102 32846 37154
rect 32898 37102 32900 37154
rect 32844 36372 32900 37102
rect 32956 36708 33012 36718
rect 32956 36594 33012 36652
rect 32956 36542 32958 36594
rect 33010 36542 33012 36594
rect 32956 36530 33012 36542
rect 32844 36306 32900 36316
rect 32844 34916 32900 34926
rect 32844 34822 32900 34860
rect 32732 33460 32788 33740
rect 32956 33460 33012 33470
rect 32732 33458 33012 33460
rect 32732 33406 32958 33458
rect 33010 33406 33012 33458
rect 32732 33404 33012 33406
rect 32956 33394 33012 33404
rect 32620 33282 32676 33292
rect 32508 33234 32564 33246
rect 32508 33182 32510 33234
rect 32562 33182 32564 33234
rect 32508 33012 32564 33182
rect 32508 32946 32564 32956
rect 32396 32734 32398 32786
rect 32450 32734 32452 32786
rect 32396 32722 32452 32734
rect 32620 32452 32676 32462
rect 32620 31780 32676 32396
rect 32732 32450 32788 32462
rect 32732 32398 32734 32450
rect 32786 32398 32788 32450
rect 32732 31948 32788 32398
rect 32732 31892 33012 31948
rect 32508 31778 32676 31780
rect 32508 31726 32622 31778
rect 32674 31726 32676 31778
rect 32508 31724 32676 31726
rect 32284 31220 32340 31230
rect 32284 28980 32340 31164
rect 32284 28914 32340 28924
rect 32396 30210 32452 30222
rect 32396 30158 32398 30210
rect 32450 30158 32452 30210
rect 32060 27858 32228 27860
rect 32060 27806 32174 27858
rect 32226 27806 32228 27858
rect 32060 27804 32228 27806
rect 31836 26852 32004 26908
rect 31948 26292 32004 26852
rect 31276 26178 31444 26180
rect 31276 26126 31278 26178
rect 31330 26126 31444 26178
rect 31276 26124 31444 26126
rect 31276 26114 31332 26124
rect 31164 26014 31166 26066
rect 31218 26014 31220 26066
rect 31164 26002 31220 26014
rect 31164 25284 31220 25294
rect 31164 25190 31220 25228
rect 31052 25106 31108 25116
rect 30828 24946 31108 24948
rect 30828 24894 30830 24946
rect 30882 24894 31108 24946
rect 30828 24892 31108 24894
rect 30380 24882 30436 24892
rect 30828 24882 30884 24892
rect 30940 23940 30996 23950
rect 30940 23846 30996 23884
rect 30156 23650 30212 23660
rect 30940 23604 30996 23614
rect 30380 23492 30436 23502
rect 30156 23044 30212 23054
rect 30156 22594 30212 22988
rect 30156 22542 30158 22594
rect 30210 22542 30212 22594
rect 30156 22530 30212 22542
rect 30380 22484 30436 23436
rect 30604 23378 30660 23390
rect 30604 23326 30606 23378
rect 30658 23326 30660 23378
rect 30604 23268 30660 23326
rect 30604 23202 30660 23212
rect 30716 23156 30772 23166
rect 30716 23062 30772 23100
rect 30940 23154 30996 23548
rect 30940 23102 30942 23154
rect 30994 23102 30996 23154
rect 30044 21298 30100 21308
rect 30268 22482 30436 22484
rect 30268 22430 30382 22482
rect 30434 22430 30436 22482
rect 30268 22428 30436 22430
rect 30268 21028 30324 22428
rect 30380 22418 30436 22428
rect 30604 22708 30660 22718
rect 30604 22370 30660 22652
rect 30604 22318 30606 22370
rect 30658 22318 30660 22370
rect 30604 22306 30660 22318
rect 30828 22372 30884 22382
rect 30828 22278 30884 22316
rect 30716 22148 30772 22158
rect 30380 22146 30772 22148
rect 30380 22094 30718 22146
rect 30770 22094 30772 22146
rect 30380 22092 30772 22094
rect 30380 21810 30436 22092
rect 30716 22082 30772 22092
rect 30380 21758 30382 21810
rect 30434 21758 30436 21810
rect 30380 21746 30436 21758
rect 30828 21812 30884 21822
rect 30828 21718 30884 21756
rect 30604 21700 30660 21710
rect 30604 21606 30660 21644
rect 30492 21474 30548 21486
rect 30940 21476 30996 23102
rect 30492 21422 30494 21474
rect 30546 21422 30548 21474
rect 30492 21364 30548 21422
rect 30492 21298 30548 21308
rect 30716 21420 30996 21476
rect 30268 20972 30660 21028
rect 29484 19282 29540 19292
rect 29708 20916 29764 20926
rect 29596 19124 29652 19134
rect 29372 18946 29428 18956
rect 29484 19010 29540 19022
rect 29484 18958 29486 19010
rect 29538 18958 29540 19010
rect 29484 18676 29540 18958
rect 29484 18610 29540 18620
rect 29596 18564 29652 19068
rect 29596 18432 29652 18508
rect 29484 18340 29540 18350
rect 29148 18338 29540 18340
rect 29148 18286 29486 18338
rect 29538 18286 29540 18338
rect 29148 18284 29540 18286
rect 29484 18274 29540 18284
rect 29036 16818 29092 16828
rect 29148 17332 29204 17342
rect 28924 15538 28980 15820
rect 28924 15486 28926 15538
rect 28978 15486 28980 15538
rect 28924 15474 28980 15486
rect 29036 16660 29092 16670
rect 28812 14254 28814 14306
rect 28866 14254 28868 14306
rect 28812 14196 28868 14254
rect 28812 14130 28868 14140
rect 28588 13918 28590 13970
rect 28642 13918 28644 13970
rect 28588 13906 28644 13918
rect 29036 12964 29092 16604
rect 29148 13970 29204 17276
rect 29372 17108 29428 17118
rect 29372 17014 29428 17052
rect 29708 16660 29764 20860
rect 30268 20802 30324 20814
rect 30268 20750 30270 20802
rect 30322 20750 30324 20802
rect 29820 20690 29876 20702
rect 29820 20638 29822 20690
rect 29874 20638 29876 20690
rect 29820 20244 29876 20638
rect 29820 20018 29876 20188
rect 29820 19966 29822 20018
rect 29874 19966 29876 20018
rect 29820 19954 29876 19966
rect 30156 20132 30212 20142
rect 30268 20132 30324 20750
rect 30156 20130 30324 20132
rect 30156 20078 30158 20130
rect 30210 20078 30324 20130
rect 30156 20076 30324 20078
rect 30156 20020 30212 20076
rect 30156 19954 30212 19964
rect 29820 19796 29876 19806
rect 29820 18564 29876 19740
rect 30380 19458 30436 19470
rect 30380 19406 30382 19458
rect 30434 19406 30436 19458
rect 30268 19348 30324 19358
rect 30268 18788 30324 19292
rect 30380 19346 30436 19406
rect 30380 19294 30382 19346
rect 30434 19294 30436 19346
rect 30380 19282 30436 19294
rect 29820 18562 30100 18564
rect 29820 18510 29822 18562
rect 29874 18510 30100 18562
rect 29820 18508 30100 18510
rect 29820 18498 29876 18508
rect 29932 18340 29988 18350
rect 29932 17106 29988 18284
rect 30044 17554 30100 18508
rect 30044 17502 30046 17554
rect 30098 17502 30100 17554
rect 30044 17490 30100 17502
rect 30156 18562 30212 18574
rect 30156 18510 30158 18562
rect 30210 18510 30212 18562
rect 29932 17054 29934 17106
rect 29986 17054 29988 17106
rect 29932 17042 29988 17054
rect 30044 17108 30100 17118
rect 30156 17108 30212 18510
rect 30268 18340 30324 18732
rect 30492 19012 30548 19022
rect 30380 18340 30436 18350
rect 30268 18338 30436 18340
rect 30268 18286 30382 18338
rect 30434 18286 30436 18338
rect 30268 18284 30436 18286
rect 30380 18274 30436 18284
rect 30492 18226 30548 18956
rect 30604 18788 30660 20972
rect 30716 19458 30772 21420
rect 30940 21028 30996 21038
rect 31052 21028 31108 24892
rect 31276 24724 31332 24734
rect 31276 24630 31332 24668
rect 31388 24612 31444 26124
rect 31724 26178 31780 26190
rect 31724 26126 31726 26178
rect 31778 26126 31780 26178
rect 31724 26066 31780 26126
rect 31724 26014 31726 26066
rect 31778 26014 31780 26066
rect 31724 24724 31780 26014
rect 31948 25620 32004 26236
rect 32060 25732 32116 27804
rect 32172 27794 32228 27804
rect 32284 28644 32340 28654
rect 32284 26964 32340 28588
rect 32396 28084 32452 30158
rect 32508 29540 32564 31724
rect 32620 31714 32676 31724
rect 32620 31220 32676 31230
rect 32620 31106 32676 31164
rect 32620 31054 32622 31106
rect 32674 31054 32676 31106
rect 32620 31042 32676 31054
rect 32732 31108 32788 31118
rect 32732 31014 32788 31052
rect 32844 30996 32900 31006
rect 32732 30772 32788 30782
rect 32732 30678 32788 30716
rect 32844 29876 32900 30940
rect 32732 29820 32900 29876
rect 32956 30548 33012 31892
rect 32732 29650 32788 29820
rect 32732 29598 32734 29650
rect 32786 29598 32788 29650
rect 32732 29586 32788 29598
rect 32508 29538 32676 29540
rect 32508 29486 32510 29538
rect 32562 29486 32676 29538
rect 32508 29484 32676 29486
rect 32508 29474 32564 29484
rect 32620 28532 32676 29484
rect 32620 28466 32676 28476
rect 32732 28980 32788 28990
rect 32508 28420 32564 28430
rect 32508 28326 32564 28364
rect 32396 28018 32452 28028
rect 32732 28082 32788 28924
rect 32956 28644 33012 30492
rect 33068 29988 33124 37884
rect 33292 37940 33348 37950
rect 33292 37846 33348 37884
rect 33404 37938 33460 38220
rect 33404 37886 33406 37938
rect 33458 37886 33460 37938
rect 33404 37874 33460 37886
rect 33292 37492 33348 37502
rect 33180 34916 33236 34926
rect 33180 34822 33236 34860
rect 33292 30772 33348 37436
rect 33516 37154 33572 38612
rect 33852 38276 33908 38286
rect 33628 37940 33684 37950
rect 33628 37846 33684 37884
rect 33516 37102 33518 37154
rect 33570 37102 33572 37154
rect 33404 36708 33460 36718
rect 33404 36482 33460 36652
rect 33404 36430 33406 36482
rect 33458 36430 33460 36482
rect 33404 36418 33460 36430
rect 33404 35700 33460 35710
rect 33404 34690 33460 35644
rect 33516 35476 33572 37102
rect 33740 37268 33796 37278
rect 33628 35476 33684 35486
rect 33516 35420 33628 35476
rect 33628 35382 33684 35420
rect 33404 34638 33406 34690
rect 33458 34638 33460 34690
rect 33404 33124 33460 34638
rect 33404 33030 33460 33068
rect 33516 35252 33572 35262
rect 33516 34802 33572 35196
rect 33516 34750 33518 34802
rect 33570 34750 33572 34802
rect 33516 34018 33572 34750
rect 33516 33966 33518 34018
rect 33570 33966 33572 34018
rect 33516 32340 33572 33966
rect 33628 34916 33684 34926
rect 33628 33124 33684 34860
rect 33740 33348 33796 37212
rect 33852 36482 33908 38220
rect 34412 38276 34468 38286
rect 34188 38052 34244 38062
rect 34188 37958 34244 37996
rect 34076 37826 34132 37838
rect 34076 37774 34078 37826
rect 34130 37774 34132 37826
rect 33964 36596 34020 36606
rect 34076 36596 34132 37774
rect 34300 37828 34356 37838
rect 34300 37734 34356 37772
rect 33964 36594 34132 36596
rect 33964 36542 33966 36594
rect 34018 36542 34132 36594
rect 33964 36540 34132 36542
rect 34188 37604 34244 37614
rect 33964 36530 34020 36540
rect 33852 36430 33854 36482
rect 33906 36430 33908 36482
rect 33852 36418 33908 36430
rect 34076 36372 34132 36382
rect 34188 36372 34244 37548
rect 34412 37378 34468 38220
rect 34524 37940 34580 37950
rect 34524 37846 34580 37884
rect 34412 37326 34414 37378
rect 34466 37326 34468 37378
rect 34412 37314 34468 37326
rect 34076 36370 34244 36372
rect 34076 36318 34078 36370
rect 34130 36318 34244 36370
rect 34076 36316 34244 36318
rect 34300 37266 34356 37278
rect 34300 37214 34302 37266
rect 34354 37214 34356 37266
rect 34300 36708 34356 37214
rect 33852 35924 33908 35934
rect 33852 35830 33908 35868
rect 33964 35700 34020 35710
rect 33964 35586 34020 35644
rect 33964 35534 33966 35586
rect 34018 35534 34020 35586
rect 33964 35522 34020 35534
rect 33740 33292 34020 33348
rect 33852 33124 33908 33134
rect 33628 33122 33908 33124
rect 33628 33070 33854 33122
rect 33906 33070 33908 33122
rect 33628 33068 33908 33070
rect 33628 32452 33684 32462
rect 33628 32358 33684 32396
rect 33516 32274 33572 32284
rect 33404 32228 33460 32238
rect 33404 31220 33460 32172
rect 33404 31154 33460 31164
rect 33516 31556 33572 31566
rect 33292 30716 33460 30772
rect 33292 30548 33348 30558
rect 33292 30210 33348 30492
rect 33292 30158 33294 30210
rect 33346 30158 33348 30210
rect 33292 30146 33348 30158
rect 33068 29932 33236 29988
rect 32956 28578 33012 28588
rect 33068 29764 33124 29774
rect 32732 28030 32734 28082
rect 32786 28030 32788 28082
rect 32508 27524 32564 27534
rect 32508 27076 32564 27468
rect 32508 27010 32564 27020
rect 32396 26964 32452 26974
rect 32284 26962 32452 26964
rect 32284 26910 32398 26962
rect 32450 26910 32452 26962
rect 32284 26908 32452 26910
rect 32172 26852 32340 26908
rect 32396 26898 32452 26908
rect 32508 26852 32564 26862
rect 32172 26514 32228 26852
rect 32508 26758 32564 26796
rect 32172 26462 32174 26514
rect 32226 26462 32228 26514
rect 32172 26450 32228 26462
rect 32732 25732 32788 28030
rect 32844 28532 32900 28542
rect 32844 27300 32900 28476
rect 33068 28420 33124 29708
rect 33180 28980 33236 29932
rect 33404 29764 33460 30716
rect 33404 29698 33460 29708
rect 33236 28924 33348 28980
rect 33180 28914 33236 28924
rect 32844 27234 32900 27244
rect 32956 28364 33124 28420
rect 33180 28418 33236 28430
rect 33180 28366 33182 28418
rect 33234 28366 33236 28418
rect 32060 25676 32340 25732
rect 31724 24658 31780 24668
rect 31836 25564 32228 25620
rect 31276 23940 31332 23950
rect 31388 23940 31444 24556
rect 31332 23884 31444 23940
rect 31164 23154 31220 23166
rect 31164 23102 31166 23154
rect 31218 23102 31220 23154
rect 31164 22708 31220 23102
rect 31164 22642 31220 22652
rect 30940 21026 31108 21028
rect 30940 20974 30942 21026
rect 30994 20974 31108 21026
rect 30940 20972 31108 20974
rect 30940 20962 30996 20972
rect 30716 19406 30718 19458
rect 30770 19406 30772 19458
rect 30716 19394 30772 19406
rect 30828 20242 30884 20254
rect 30828 20190 30830 20242
rect 30882 20190 30884 20242
rect 30604 18722 30660 18732
rect 30716 19012 30772 19022
rect 30492 18174 30494 18226
rect 30546 18174 30548 18226
rect 30044 17106 30212 17108
rect 30044 17054 30046 17106
rect 30098 17054 30212 17106
rect 30044 17052 30212 17054
rect 30268 17556 30324 17566
rect 30044 17042 30100 17052
rect 29484 16604 29708 16660
rect 29484 15988 29540 16604
rect 29708 16594 29764 16604
rect 30156 16882 30212 16894
rect 30156 16830 30158 16882
rect 30210 16830 30212 16882
rect 30156 16436 30212 16830
rect 29708 16380 30212 16436
rect 29708 16322 29764 16380
rect 29708 16270 29710 16322
rect 29762 16270 29764 16322
rect 29708 16258 29764 16270
rect 29596 16212 29652 16222
rect 29596 16118 29652 16156
rect 29484 15932 29764 15988
rect 29372 15876 29428 15886
rect 29372 15538 29428 15820
rect 29372 15486 29374 15538
rect 29426 15486 29428 15538
rect 29372 15474 29428 15486
rect 29596 15092 29652 15102
rect 29148 13918 29150 13970
rect 29202 13918 29204 13970
rect 29148 13906 29204 13918
rect 29484 14420 29540 14430
rect 28364 12646 28420 12684
rect 28700 12908 29036 12964
rect 28588 12628 28644 12638
rect 28028 12404 28084 12414
rect 27916 12402 28084 12404
rect 27916 12350 28030 12402
rect 28082 12350 28084 12402
rect 27916 12348 28084 12350
rect 28028 12338 28084 12348
rect 28588 12068 28644 12572
rect 28700 12402 28756 12908
rect 29036 12898 29092 12908
rect 28812 12738 28868 12750
rect 28812 12686 28814 12738
rect 28866 12686 28868 12738
rect 28812 12628 28868 12686
rect 28812 12562 28868 12572
rect 29484 12628 29540 14364
rect 29596 14084 29652 15036
rect 29596 13970 29652 14028
rect 29596 13918 29598 13970
rect 29650 13918 29652 13970
rect 29596 13906 29652 13918
rect 29708 14418 29764 15932
rect 29708 14366 29710 14418
rect 29762 14366 29764 14418
rect 29708 13522 29764 14366
rect 29820 13860 29876 16380
rect 30156 15092 30212 15102
rect 30044 15090 30212 15092
rect 30044 15038 30158 15090
rect 30210 15038 30212 15090
rect 30044 15036 30212 15038
rect 29932 14420 29988 14430
rect 29932 14326 29988 14364
rect 30044 14306 30100 15036
rect 30156 15026 30212 15036
rect 30268 15092 30324 17500
rect 30268 15026 30324 15036
rect 30380 16772 30436 16782
rect 30380 15986 30436 16716
rect 30492 16436 30548 18174
rect 30604 18452 30660 18462
rect 30604 17556 30660 18396
rect 30604 17424 30660 17500
rect 30604 16882 30660 16894
rect 30604 16830 30606 16882
rect 30658 16830 30660 16882
rect 30604 16770 30660 16830
rect 30604 16718 30606 16770
rect 30658 16718 30660 16770
rect 30604 16706 30660 16718
rect 30492 16370 30548 16380
rect 30604 16548 30660 16558
rect 30604 16322 30660 16492
rect 30604 16270 30606 16322
rect 30658 16270 30660 16322
rect 30604 16258 30660 16270
rect 30716 16212 30772 18956
rect 30828 17890 30884 20190
rect 30828 17838 30830 17890
rect 30882 17838 30884 17890
rect 30828 17556 30884 17838
rect 30828 17490 30884 17500
rect 30940 20018 30996 20030
rect 30940 19966 30942 20018
rect 30994 19966 30996 20018
rect 30940 19348 30996 19966
rect 30940 17108 30996 19292
rect 31052 18564 31108 20972
rect 31164 19460 31220 19470
rect 31164 19346 31220 19404
rect 31164 19294 31166 19346
rect 31218 19294 31220 19346
rect 31164 19282 31220 19294
rect 31052 18498 31108 18508
rect 31164 18788 31220 18798
rect 31052 18340 31108 18350
rect 31164 18340 31220 18732
rect 31276 18676 31332 23884
rect 31388 23154 31444 23166
rect 31388 23102 31390 23154
rect 31442 23102 31444 23154
rect 31388 22372 31444 23102
rect 31836 22596 31892 25564
rect 32172 25506 32228 25564
rect 32172 25454 32174 25506
rect 32226 25454 32228 25506
rect 32172 25442 32228 25454
rect 32060 25396 32116 25406
rect 32060 25302 32116 25340
rect 32284 25284 32340 25676
rect 32284 25218 32340 25228
rect 32396 25676 32788 25732
rect 32844 27076 32900 27086
rect 32844 25732 32900 27020
rect 32956 26514 33012 28364
rect 32956 26462 32958 26514
rect 33010 26462 33012 26514
rect 32956 26450 33012 26462
rect 33068 28196 33124 28206
rect 32844 25676 33012 25732
rect 31612 22540 31892 22596
rect 31948 25172 32004 25182
rect 31948 23938 32004 25116
rect 32172 25060 32228 25070
rect 32396 25060 32452 25676
rect 32844 25508 32900 25518
rect 32844 25414 32900 25452
rect 32228 25004 32452 25060
rect 32508 25284 32564 25294
rect 32060 24948 32116 24958
rect 32060 24854 32116 24892
rect 31948 23886 31950 23938
rect 32002 23886 32004 23938
rect 31612 22482 31668 22540
rect 31612 22430 31614 22482
rect 31666 22430 31668 22482
rect 31612 22418 31668 22430
rect 31388 21476 31444 22316
rect 31612 21476 31668 21486
rect 31388 21474 31668 21476
rect 31388 21422 31614 21474
rect 31666 21422 31668 21474
rect 31388 21420 31668 21422
rect 31276 18610 31332 18620
rect 31388 20132 31444 20142
rect 31052 18338 31220 18340
rect 31052 18286 31054 18338
rect 31106 18286 31220 18338
rect 31052 18284 31220 18286
rect 31052 18274 31108 18284
rect 31164 17444 31220 17454
rect 31164 17350 31220 17388
rect 31052 17108 31108 17118
rect 30940 17106 31108 17108
rect 30940 17054 31054 17106
rect 31106 17054 31108 17106
rect 30940 17052 31108 17054
rect 31052 17042 31108 17052
rect 31388 17106 31444 20076
rect 31500 18788 31556 21420
rect 31612 21410 31668 21420
rect 31612 21028 31668 21038
rect 31612 20934 31668 20972
rect 31724 20244 31780 22540
rect 31948 22484 32004 23886
rect 32172 23828 32228 25004
rect 32508 24610 32564 25228
rect 32956 25172 33012 25676
rect 33068 25508 33124 28140
rect 33180 28084 33236 28366
rect 33180 28018 33236 28028
rect 33180 25620 33236 25630
rect 33180 25526 33236 25564
rect 33068 25442 33124 25452
rect 32508 24558 32510 24610
rect 32562 24558 32564 24610
rect 32396 24162 32452 24174
rect 32396 24110 32398 24162
rect 32450 24110 32452 24162
rect 32396 24052 32452 24110
rect 32396 23986 32452 23996
rect 32172 23826 32340 23828
rect 32172 23774 32174 23826
rect 32226 23774 32340 23826
rect 32172 23772 32340 23774
rect 32172 23762 32228 23772
rect 31836 22428 32004 22484
rect 32060 23492 32116 23502
rect 32060 23378 32116 23436
rect 32060 23326 32062 23378
rect 32114 23326 32116 23378
rect 32060 22484 32116 23326
rect 32172 23268 32228 23306
rect 32172 23202 32228 23212
rect 31836 20804 31892 22428
rect 32060 22418 32116 22428
rect 32172 23042 32228 23054
rect 32172 22990 32174 23042
rect 32226 22990 32228 23042
rect 32172 21812 32228 22990
rect 32284 23044 32340 23772
rect 32396 23716 32452 23726
rect 32396 23492 32452 23660
rect 32396 23378 32452 23436
rect 32396 23326 32398 23378
rect 32450 23326 32452 23378
rect 32396 23314 32452 23326
rect 32284 22988 32452 23044
rect 32284 22820 32340 22830
rect 32284 22482 32340 22764
rect 32284 22430 32286 22482
rect 32338 22430 32340 22482
rect 32284 22418 32340 22430
rect 32396 22148 32452 22988
rect 32172 21746 32228 21756
rect 32284 22092 32452 22148
rect 31948 21700 32004 21710
rect 31948 21026 32004 21644
rect 31948 20974 31950 21026
rect 32002 20974 32004 21026
rect 31948 20962 32004 20974
rect 31836 20748 32004 20804
rect 31836 20578 31892 20590
rect 31836 20526 31838 20578
rect 31890 20526 31892 20578
rect 31836 20468 31892 20526
rect 31836 20402 31892 20412
rect 31612 20188 31780 20244
rect 31836 20244 31892 20254
rect 31948 20244 32004 20748
rect 31836 20242 32004 20244
rect 31836 20190 31838 20242
rect 31890 20190 32004 20242
rect 31836 20188 32004 20190
rect 31612 19236 31668 20188
rect 31836 20132 31892 20188
rect 31836 20066 31892 20076
rect 32060 20130 32116 20142
rect 32060 20078 32062 20130
rect 32114 20078 32116 20130
rect 31724 20020 31780 20030
rect 31724 19926 31780 19964
rect 32060 19796 32116 20078
rect 32060 19730 32116 19740
rect 32284 20020 32340 22092
rect 32508 22036 32564 24558
rect 32732 25060 32788 25070
rect 32732 23380 32788 25004
rect 32732 23314 32788 23324
rect 32844 24836 32900 24846
rect 32620 23154 32676 23166
rect 32620 23102 32622 23154
rect 32674 23102 32676 23154
rect 32620 22932 32676 23102
rect 32620 22866 32676 22876
rect 32844 22820 32900 24780
rect 32844 22754 32900 22764
rect 32956 22596 33012 25116
rect 32620 22540 33012 22596
rect 33292 25396 33348 28924
rect 33516 27972 33572 31500
rect 33740 31220 33796 31230
rect 33740 31106 33796 31164
rect 33740 31054 33742 31106
rect 33794 31054 33796 31106
rect 33628 30212 33684 30222
rect 33740 30212 33796 31054
rect 33684 30156 33796 30212
rect 33628 30080 33684 30156
rect 33852 30100 33908 33068
rect 33964 31948 34020 33292
rect 34076 32116 34132 36316
rect 34188 34690 34244 34702
rect 34188 34638 34190 34690
rect 34242 34638 34244 34690
rect 34188 34132 34244 34638
rect 34300 34468 34356 36652
rect 34524 36596 34580 36606
rect 34636 36596 34692 38612
rect 34524 36594 34692 36596
rect 34524 36542 34526 36594
rect 34578 36542 34692 36594
rect 34524 36540 34692 36542
rect 34524 35924 34580 36540
rect 34524 35858 34580 35868
rect 34636 35700 34692 35710
rect 34524 34916 34580 34954
rect 34524 34850 34580 34860
rect 34300 34402 34356 34412
rect 34524 34692 34580 34702
rect 34412 34132 34468 34142
rect 34188 34130 34468 34132
rect 34188 34078 34414 34130
rect 34466 34078 34468 34130
rect 34188 34076 34468 34078
rect 34412 34066 34468 34076
rect 34524 33572 34580 34636
rect 34636 34130 34692 35644
rect 34636 34078 34638 34130
rect 34690 34078 34692 34130
rect 34636 34066 34692 34078
rect 34076 32050 34132 32060
rect 34300 33516 34580 33572
rect 34748 33570 34804 39564
rect 34972 37940 35028 39564
rect 35084 39618 35140 39900
rect 35084 39566 35086 39618
rect 35138 39566 35140 39618
rect 35084 39554 35140 39566
rect 35532 38834 35588 40124
rect 35532 38782 35534 38834
rect 35586 38782 35588 38834
rect 35532 38770 35588 38782
rect 35196 38722 35252 38734
rect 35196 38670 35198 38722
rect 35250 38670 35252 38722
rect 35196 38668 35252 38670
rect 35644 38668 35700 40238
rect 35756 39956 35812 42588
rect 35868 41972 35924 41982
rect 35868 41878 35924 41916
rect 35980 41188 36036 41198
rect 35980 41094 36036 41132
rect 35980 40628 36036 40638
rect 35980 40534 36036 40572
rect 36092 40292 36148 43652
rect 36204 43652 36260 43662
rect 36204 42978 36260 43596
rect 36540 43428 36596 43438
rect 36204 42926 36206 42978
rect 36258 42926 36260 42978
rect 36204 42914 36260 42926
rect 36428 43426 36596 43428
rect 36428 43374 36542 43426
rect 36594 43374 36596 43426
rect 36428 43372 36596 43374
rect 36092 40226 36148 40236
rect 36204 42756 36260 42766
rect 36204 41186 36260 42700
rect 36204 41134 36206 41186
rect 36258 41134 36260 41186
rect 36204 40178 36260 41134
rect 36428 42532 36484 43372
rect 36540 43362 36596 43372
rect 36652 42756 36708 44940
rect 36652 42690 36708 42700
rect 36428 41300 36484 42476
rect 36540 42084 36596 42094
rect 36540 41990 36596 42028
rect 36428 41186 36484 41244
rect 36540 41300 36596 41310
rect 36764 41300 36820 45836
rect 36876 45668 36932 46396
rect 37100 45780 37156 48076
rect 36876 45602 36932 45612
rect 36988 45724 37100 45780
rect 36876 43426 36932 43438
rect 36876 43374 36878 43426
rect 36930 43374 36932 43426
rect 36876 41748 36932 43374
rect 36876 41682 36932 41692
rect 36988 41524 37044 45724
rect 37100 45714 37156 45724
rect 37100 45556 37156 45566
rect 37100 45330 37156 45500
rect 37100 45278 37102 45330
rect 37154 45278 37156 45330
rect 37100 45266 37156 45278
rect 36540 41298 36820 41300
rect 36540 41246 36542 41298
rect 36594 41246 36820 41298
rect 36540 41244 36820 41246
rect 36876 41468 37044 41524
rect 37100 42082 37156 42094
rect 37100 42030 37102 42082
rect 37154 42030 37156 42082
rect 36540 41234 36596 41244
rect 36428 41134 36430 41186
rect 36482 41134 36484 41186
rect 36428 41122 36484 41134
rect 36652 40962 36708 40974
rect 36652 40910 36654 40962
rect 36706 40910 36708 40962
rect 36204 40126 36206 40178
rect 36258 40126 36260 40178
rect 36204 40114 36260 40126
rect 36316 40740 36372 40750
rect 35756 39900 36260 39956
rect 36092 39620 36148 39630
rect 36092 39526 36148 39564
rect 35868 39508 35924 39518
rect 35868 38668 35924 39452
rect 35980 39394 36036 39406
rect 35980 39342 35982 39394
rect 36034 39342 36036 39394
rect 35980 38834 36036 39342
rect 35980 38782 35982 38834
rect 36034 38782 36036 38834
rect 35980 38770 36036 38782
rect 36204 38668 36260 39900
rect 36316 39058 36372 40684
rect 36428 40402 36484 40414
rect 36428 40350 36430 40402
rect 36482 40350 36484 40402
rect 36428 40292 36484 40350
rect 36652 40292 36708 40910
rect 36876 40516 36932 41468
rect 37100 41412 37156 42030
rect 37100 41346 37156 41356
rect 36484 40236 36596 40292
rect 36428 40226 36484 40236
rect 36428 40068 36484 40078
rect 36428 39618 36484 40012
rect 36428 39566 36430 39618
rect 36482 39566 36484 39618
rect 36428 39554 36484 39566
rect 36316 39006 36318 39058
rect 36370 39006 36372 39058
rect 36316 38994 36372 39006
rect 36540 39060 36596 40236
rect 36652 40226 36708 40236
rect 36764 40460 36932 40516
rect 36988 40964 37044 40974
rect 36540 38994 36596 39004
rect 36652 39060 36708 39070
rect 36764 39060 36820 40460
rect 36652 39058 36820 39060
rect 36652 39006 36654 39058
rect 36706 39006 36820 39058
rect 36652 39004 36820 39006
rect 36876 40290 36932 40302
rect 36876 40238 36878 40290
rect 36930 40238 36932 40290
rect 36876 40178 36932 40238
rect 36876 40126 36878 40178
rect 36930 40126 36932 40178
rect 36652 38668 36708 39004
rect 36876 38948 36932 40126
rect 34972 37874 35028 37884
rect 35084 38612 35700 38668
rect 35756 38612 35924 38668
rect 36092 38612 36260 38668
rect 36540 38612 36708 38668
rect 36764 38892 36932 38948
rect 35084 37268 35140 38612
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35756 38388 35812 38612
rect 35196 38378 35460 38388
rect 35532 38332 35812 38388
rect 35420 38276 35476 38286
rect 35532 38276 35588 38332
rect 35420 38274 35588 38276
rect 35420 38222 35422 38274
rect 35474 38222 35588 38274
rect 35420 38220 35588 38222
rect 35420 38210 35476 38220
rect 35196 38050 35252 38062
rect 35196 37998 35198 38050
rect 35250 37998 35252 38050
rect 35196 37940 35252 37998
rect 35196 37874 35252 37884
rect 35756 37826 35812 37838
rect 35756 37774 35758 37826
rect 35810 37774 35812 37826
rect 35308 37604 35364 37614
rect 35308 37490 35364 37548
rect 35308 37438 35310 37490
rect 35362 37438 35364 37490
rect 35308 37426 35364 37438
rect 35084 37202 35140 37212
rect 34860 37154 34916 37166
rect 34860 37102 34862 37154
rect 34914 37102 34916 37154
rect 34860 36484 34916 37102
rect 35756 37156 35812 37774
rect 35980 37156 36036 37166
rect 35756 37154 36036 37156
rect 35756 37102 35982 37154
rect 36034 37102 36036 37154
rect 35756 37100 36036 37102
rect 35980 37090 36036 37100
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35868 36596 35924 36606
rect 36092 36596 36148 38612
rect 36316 38164 36372 38174
rect 36316 38070 36372 38108
rect 35868 36594 36148 36596
rect 35868 36542 35870 36594
rect 35922 36542 36148 36594
rect 35868 36540 36148 36542
rect 36204 37828 36260 37838
rect 36204 37378 36260 37772
rect 36540 37828 36596 38612
rect 36540 37762 36596 37772
rect 36652 37826 36708 37838
rect 36652 37774 36654 37826
rect 36706 37774 36708 37826
rect 36204 37326 36206 37378
rect 36258 37326 36260 37378
rect 36204 37044 36260 37326
rect 35868 36530 35924 36540
rect 34860 36418 34916 36428
rect 35308 36484 35364 36494
rect 35308 36390 35364 36428
rect 35756 36258 35812 36270
rect 35756 36206 35758 36258
rect 35810 36206 35812 36258
rect 35756 36036 35812 36206
rect 35980 36260 36036 36270
rect 35980 36166 36036 36204
rect 35756 35970 35812 35980
rect 34972 35924 35028 35934
rect 34972 35830 35028 35868
rect 36204 35812 36260 36988
rect 36428 36708 36484 36718
rect 36652 36708 36708 37774
rect 36484 36652 36708 36708
rect 36428 36594 36484 36652
rect 36428 36542 36430 36594
rect 36482 36542 36484 36594
rect 36428 36530 36484 36542
rect 35980 35756 36260 35812
rect 36652 36260 36708 36270
rect 34860 35698 34916 35710
rect 34860 35646 34862 35698
rect 34914 35646 34916 35698
rect 34860 34916 34916 35646
rect 35084 35698 35140 35710
rect 35084 35646 35086 35698
rect 35138 35646 35140 35698
rect 35084 35588 35140 35646
rect 35308 35700 35364 35710
rect 35308 35698 35812 35700
rect 35308 35646 35310 35698
rect 35362 35646 35812 35698
rect 35308 35644 35812 35646
rect 35308 35634 35364 35644
rect 34860 34850 34916 34860
rect 34972 34914 35028 34926
rect 34972 34862 34974 34914
rect 35026 34862 35028 34914
rect 34748 33518 34750 33570
rect 34802 33518 34804 33570
rect 34300 33458 34356 33516
rect 34748 33460 34804 33518
rect 34300 33406 34302 33458
rect 34354 33406 34356 33458
rect 33964 31892 34244 31948
rect 34188 31890 34244 31892
rect 34188 31838 34190 31890
rect 34242 31838 34244 31890
rect 34188 31826 34244 31838
rect 34076 31778 34132 31790
rect 34076 31726 34078 31778
rect 34130 31726 34132 31778
rect 34076 31108 34132 31726
rect 34076 30210 34132 31052
rect 34188 30996 34244 31006
rect 34300 30996 34356 33406
rect 34524 33404 34804 33460
rect 34860 34468 34916 34478
rect 34524 32786 34580 33404
rect 34860 33348 34916 34412
rect 34972 34132 35028 34862
rect 35084 34802 35140 35532
rect 35756 35586 35812 35644
rect 35756 35534 35758 35586
rect 35810 35534 35812 35586
rect 35532 35476 35588 35486
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35084 34750 35086 34802
rect 35138 34750 35140 34802
rect 35084 34692 35140 34750
rect 35084 34626 35140 34636
rect 35196 34468 35252 34478
rect 35196 34244 35252 34412
rect 35308 34244 35364 34254
rect 35196 34242 35364 34244
rect 35196 34190 35310 34242
rect 35362 34190 35364 34242
rect 35196 34188 35364 34190
rect 35308 34178 35364 34188
rect 35084 34132 35140 34142
rect 34972 34076 35084 34132
rect 34748 33292 34916 33348
rect 34748 33236 34804 33292
rect 34524 32734 34526 32786
rect 34578 32734 34580 32786
rect 34524 32722 34580 32734
rect 34636 33234 34804 33236
rect 34636 33182 34750 33234
rect 34802 33182 34804 33234
rect 34636 33180 34804 33182
rect 34412 32564 34468 32574
rect 34636 32564 34692 33180
rect 34748 33170 34804 33180
rect 34412 32562 34692 32564
rect 34412 32510 34414 32562
rect 34466 32510 34692 32562
rect 34412 32508 34692 32510
rect 34748 32562 34804 32574
rect 34748 32510 34750 32562
rect 34802 32510 34804 32562
rect 34412 32228 34468 32508
rect 34412 32162 34468 32172
rect 34524 32340 34580 32350
rect 34412 31780 34468 31790
rect 34412 31686 34468 31724
rect 34188 30994 34356 30996
rect 34188 30942 34190 30994
rect 34242 30942 34356 30994
rect 34188 30940 34356 30942
rect 34188 30930 34244 30940
rect 34300 30884 34356 30940
rect 34300 30818 34356 30828
rect 34076 30158 34078 30210
rect 34130 30158 34132 30210
rect 34076 30146 34132 30158
rect 34300 30212 34356 30222
rect 33740 30044 33908 30100
rect 33628 29540 33684 29550
rect 33628 29446 33684 29484
rect 33740 28980 33796 30044
rect 33852 29764 33908 29774
rect 33852 29650 33908 29708
rect 33852 29598 33854 29650
rect 33906 29598 33908 29650
rect 33852 29586 33908 29598
rect 33964 29204 34020 29214
rect 33964 29202 34132 29204
rect 33964 29150 33966 29202
rect 34018 29150 34132 29202
rect 33964 29148 34132 29150
rect 33964 29138 34020 29148
rect 33740 28924 34020 28980
rect 33852 28756 33908 28766
rect 33852 28084 33908 28700
rect 33852 28018 33908 28028
rect 33628 27972 33684 27982
rect 33516 27970 33684 27972
rect 33516 27918 33630 27970
rect 33682 27918 33684 27970
rect 33516 27916 33684 27918
rect 33516 26908 33572 27916
rect 33628 27906 33684 27916
rect 33852 27634 33908 27646
rect 33852 27582 33854 27634
rect 33906 27582 33908 27634
rect 33852 27412 33908 27582
rect 33852 27346 33908 27356
rect 32620 22482 32676 22540
rect 32620 22430 32622 22482
rect 32674 22430 32676 22482
rect 32620 22418 32676 22430
rect 32732 22148 32788 22540
rect 33292 22484 33348 25340
rect 33404 26852 33572 26908
rect 33852 27076 33908 27086
rect 33404 24050 33460 26852
rect 33740 26292 33796 26302
rect 33404 23998 33406 24050
rect 33458 23998 33460 24050
rect 33404 23268 33460 23998
rect 33404 23202 33460 23212
rect 33516 25508 33572 25518
rect 33516 23044 33572 25452
rect 33740 24052 33796 26236
rect 33852 26290 33908 27020
rect 33964 26740 34020 28924
rect 34076 26908 34132 29148
rect 34188 28530 34244 28542
rect 34188 28478 34190 28530
rect 34242 28478 34244 28530
rect 34188 28308 34244 28478
rect 34188 28242 34244 28252
rect 34188 28084 34244 28094
rect 34188 27990 34244 28028
rect 34188 27076 34244 27086
rect 34300 27076 34356 30156
rect 34524 30100 34580 32284
rect 34524 29426 34580 30044
rect 34636 32116 34692 32126
rect 34636 30994 34692 32060
rect 34636 30942 34638 30994
rect 34690 30942 34692 30994
rect 34636 30212 34692 30942
rect 34748 30436 34804 32510
rect 34972 31668 35028 31678
rect 34972 30994 35028 31612
rect 34972 30942 34974 30994
rect 35026 30942 35028 30994
rect 34972 30548 35028 30942
rect 34972 30482 35028 30492
rect 35084 30436 35140 34076
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 33570 35252 33582
rect 35196 33518 35198 33570
rect 35250 33518 35252 33570
rect 35196 33458 35252 33518
rect 35196 33406 35198 33458
rect 35250 33406 35252 33458
rect 35196 33394 35252 33406
rect 35532 33012 35588 35420
rect 35756 35364 35812 35534
rect 35756 35298 35812 35308
rect 35868 34916 35924 34926
rect 35868 34822 35924 34860
rect 35756 34132 35812 34142
rect 35756 34038 35812 34076
rect 35980 33348 36036 35756
rect 36204 35588 36260 35598
rect 36204 35494 36260 35532
rect 36652 34916 36708 36204
rect 36764 35140 36820 38892
rect 36876 38612 36932 38622
rect 36876 37156 36932 38556
rect 36876 37090 36932 37100
rect 36876 36036 36932 36046
rect 36876 35698 36932 35980
rect 36876 35646 36878 35698
rect 36930 35646 36932 35698
rect 36876 35634 36932 35646
rect 36988 35476 37044 40908
rect 37100 39060 37156 39070
rect 37100 38724 37156 39004
rect 37100 38658 37156 38668
rect 37100 35588 37156 35598
rect 37100 35494 37156 35532
rect 36988 35410 37044 35420
rect 36764 35074 36820 35084
rect 36652 34860 36932 34916
rect 36092 34804 36148 34814
rect 36092 34020 36148 34748
rect 36204 34802 36260 34814
rect 36204 34750 36206 34802
rect 36258 34750 36260 34802
rect 36204 34244 36260 34750
rect 36764 34690 36820 34702
rect 36764 34638 36766 34690
rect 36818 34638 36820 34690
rect 36652 34356 36708 34366
rect 36652 34262 36708 34300
rect 36204 34178 36260 34188
rect 36764 34132 36820 34638
rect 36764 34066 36820 34076
rect 36204 34020 36260 34030
rect 36092 34018 36260 34020
rect 36092 33966 36206 34018
rect 36258 33966 36260 34018
rect 36092 33964 36260 33966
rect 36204 33954 36260 33964
rect 36876 34020 36932 34860
rect 37100 34020 37156 34030
rect 36876 34018 37156 34020
rect 36876 33966 37102 34018
rect 37154 33966 37156 34018
rect 36876 33964 37156 33966
rect 35980 33216 36036 33292
rect 36316 33236 36372 33246
rect 36316 33142 36372 33180
rect 36428 33124 36484 33134
rect 36428 33030 36484 33068
rect 36540 33122 36596 33134
rect 36540 33070 36542 33122
rect 36594 33070 36596 33122
rect 36540 33012 36596 33070
rect 36876 33012 36932 33964
rect 37100 33954 37156 33964
rect 35420 32956 35812 33012
rect 36540 32956 36932 33012
rect 35420 32674 35476 32956
rect 35420 32622 35422 32674
rect 35474 32622 35476 32674
rect 35420 32610 35476 32622
rect 35532 32788 35588 32798
rect 35308 32564 35364 32574
rect 35308 32470 35364 32508
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35532 32004 35588 32732
rect 35532 31938 35588 31948
rect 35644 32452 35700 32462
rect 35196 31892 35252 31902
rect 35196 31220 35252 31836
rect 35308 31220 35364 31230
rect 35196 31218 35364 31220
rect 35196 31166 35310 31218
rect 35362 31166 35364 31218
rect 35196 31164 35364 31166
rect 35308 31154 35364 31164
rect 35644 31106 35700 32396
rect 35644 31054 35646 31106
rect 35698 31054 35700 31106
rect 35644 31042 35700 31054
rect 35644 30772 35700 30782
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35532 30436 35588 30446
rect 35084 30380 35252 30436
rect 34748 30370 34804 30380
rect 34636 30156 35028 30212
rect 34636 29988 34692 30156
rect 34636 29922 34692 29932
rect 34972 29652 35028 30156
rect 34972 29586 35028 29596
rect 35084 29764 35140 29774
rect 34748 29428 34804 29438
rect 34524 29374 34526 29426
rect 34578 29374 34580 29426
rect 34524 29092 34580 29374
rect 34524 29026 34580 29036
rect 34636 29426 34804 29428
rect 34636 29374 34750 29426
rect 34802 29374 34804 29426
rect 34636 29372 34804 29374
rect 34524 28756 34580 28766
rect 34524 28530 34580 28700
rect 34524 28478 34526 28530
rect 34578 28478 34580 28530
rect 34524 28466 34580 28478
rect 34636 28532 34692 29372
rect 34748 29362 34804 29372
rect 34972 29428 35028 29438
rect 34860 29314 34916 29326
rect 34860 29262 34862 29314
rect 34914 29262 34916 29314
rect 34748 28980 34804 28990
rect 34748 28866 34804 28924
rect 34748 28814 34750 28866
rect 34802 28814 34804 28866
rect 34748 28802 34804 28814
rect 34636 28466 34692 28476
rect 34188 27074 34356 27076
rect 34188 27022 34190 27074
rect 34242 27022 34356 27074
rect 34188 27020 34356 27022
rect 34188 27010 34244 27020
rect 34076 26852 34244 26908
rect 33964 26674 34020 26684
rect 33964 26404 34020 26414
rect 33964 26310 34020 26348
rect 33852 26238 33854 26290
rect 33906 26238 33908 26290
rect 33852 24612 33908 26238
rect 34076 26290 34132 26302
rect 34076 26238 34078 26290
rect 34130 26238 34132 26290
rect 33964 25620 34020 25630
rect 34076 25620 34132 26238
rect 34020 25564 34132 25620
rect 34188 26290 34244 26852
rect 34188 26238 34190 26290
rect 34242 26238 34244 26290
rect 33964 25526 34020 25564
rect 34188 25506 34244 26238
rect 34300 25620 34356 27020
rect 34748 27748 34804 27758
rect 34748 27188 34804 27692
rect 34748 27074 34804 27132
rect 34748 27022 34750 27074
rect 34802 27022 34804 27074
rect 34748 27010 34804 27022
rect 34300 25554 34356 25564
rect 34412 26964 34468 26974
rect 34188 25454 34190 25506
rect 34242 25454 34244 25506
rect 34188 25442 34244 25454
rect 33964 25172 34020 25182
rect 33964 24834 34020 25116
rect 33964 24782 33966 24834
rect 34018 24782 34020 24834
rect 33964 24770 34020 24782
rect 34300 25172 34356 25182
rect 34188 24724 34244 24734
rect 33852 24556 34020 24612
rect 33852 24052 33908 24062
rect 33740 24050 33908 24052
rect 33740 23998 33854 24050
rect 33906 23998 33908 24050
rect 33740 23996 33908 23998
rect 33852 23986 33908 23996
rect 33628 23380 33684 23390
rect 33964 23380 34020 24556
rect 33628 23378 34020 23380
rect 33628 23326 33630 23378
rect 33682 23326 34020 23378
rect 33628 23324 34020 23326
rect 34076 23716 34132 23726
rect 33628 23314 33684 23324
rect 33964 23044 34020 23054
rect 33516 23042 34020 23044
rect 33516 22990 33966 23042
rect 34018 22990 34020 23042
rect 33516 22988 34020 22990
rect 32732 22082 32788 22092
rect 32844 22428 33348 22484
rect 31612 19180 31780 19236
rect 31612 19012 31668 19022
rect 31612 18918 31668 18956
rect 31500 18722 31556 18732
rect 31612 18676 31668 18686
rect 31500 18452 31556 18462
rect 31500 18358 31556 18396
rect 31388 17054 31390 17106
rect 31442 17054 31444 17106
rect 31388 17042 31444 17054
rect 31500 17444 31556 17454
rect 31612 17444 31668 18620
rect 31724 17668 31780 19180
rect 32060 19010 32116 19022
rect 32060 18958 32062 19010
rect 32114 18958 32116 19010
rect 32060 18788 32116 18958
rect 32060 18722 32116 18732
rect 32172 18564 32228 18574
rect 31724 17602 31780 17612
rect 31836 18228 31892 18238
rect 31612 17388 31780 17444
rect 31276 16658 31332 16670
rect 31276 16606 31278 16658
rect 31330 16606 31332 16658
rect 31276 16322 31332 16606
rect 31276 16270 31278 16322
rect 31330 16270 31332 16322
rect 31276 16258 31332 16270
rect 30716 16146 30772 16156
rect 30828 16156 31220 16212
rect 30380 15934 30382 15986
rect 30434 15934 30436 15986
rect 30156 14756 30212 14766
rect 30156 14662 30212 14700
rect 30380 14420 30436 15934
rect 30492 15874 30548 15886
rect 30492 15822 30494 15874
rect 30546 15822 30548 15874
rect 30492 15314 30548 15822
rect 30716 15540 30772 15550
rect 30828 15540 30884 16156
rect 31164 16098 31220 16156
rect 31164 16046 31166 16098
rect 31218 16046 31220 16098
rect 31164 16034 31220 16046
rect 31276 16100 31332 16110
rect 31276 15986 31332 16044
rect 31276 15934 31278 15986
rect 31330 15934 31332 15986
rect 31276 15922 31332 15934
rect 30716 15538 30884 15540
rect 30716 15486 30718 15538
rect 30770 15486 30884 15538
rect 30716 15484 30884 15486
rect 31052 15764 31108 15774
rect 30716 15474 30772 15484
rect 30492 15262 30494 15314
rect 30546 15262 30548 15314
rect 30492 15250 30548 15262
rect 30604 15314 30660 15326
rect 30604 15262 30606 15314
rect 30658 15262 30660 15314
rect 30604 14754 30660 15262
rect 30828 15314 30884 15326
rect 30828 15262 30830 15314
rect 30882 15262 30884 15314
rect 30828 15092 30884 15262
rect 30828 15026 30884 15036
rect 30604 14702 30606 14754
rect 30658 14702 30660 14754
rect 30380 14354 30436 14364
rect 30492 14644 30548 14654
rect 30492 14530 30548 14588
rect 30492 14478 30494 14530
rect 30546 14478 30548 14530
rect 30044 14254 30046 14306
rect 30098 14254 30100 14306
rect 30044 14242 30100 14254
rect 29820 13804 30212 13860
rect 30044 13636 30100 13646
rect 29708 13470 29710 13522
rect 29762 13470 29764 13522
rect 29708 13458 29764 13470
rect 29932 13634 30100 13636
rect 29932 13582 30046 13634
rect 30098 13582 30100 13634
rect 29932 13580 30100 13582
rect 29932 13522 29988 13580
rect 30044 13570 30100 13580
rect 29932 13470 29934 13522
rect 29986 13470 29988 13522
rect 29484 12562 29540 12572
rect 29708 12962 29764 12974
rect 29708 12910 29710 12962
rect 29762 12910 29764 12962
rect 28700 12350 28702 12402
rect 28754 12350 28756 12402
rect 28700 12338 28756 12350
rect 28812 12180 28868 12190
rect 29596 12180 29652 12190
rect 28812 12178 29652 12180
rect 28812 12126 28814 12178
rect 28866 12126 29598 12178
rect 29650 12126 29652 12178
rect 28812 12124 29652 12126
rect 28812 12114 28868 12124
rect 29596 12114 29652 12124
rect 28588 12002 28644 12012
rect 28924 11956 28980 11966
rect 29708 11956 29764 12910
rect 28924 11954 29764 11956
rect 28924 11902 28926 11954
rect 28978 11902 29764 11954
rect 28924 11900 29764 11902
rect 29820 12964 29876 12974
rect 28924 11890 28980 11900
rect 27468 11788 27860 11844
rect 27468 11394 27524 11788
rect 28364 11508 28420 11518
rect 28364 11414 28420 11452
rect 27468 11342 27470 11394
rect 27522 11342 27524 11394
rect 27468 11330 27524 11342
rect 27804 11170 27860 11182
rect 27804 11118 27806 11170
rect 27858 11118 27860 11170
rect 27804 11060 27860 11118
rect 27356 9998 27358 10050
rect 27410 9998 27412 10050
rect 27356 9986 27412 9998
rect 27468 10498 27524 10510
rect 27468 10446 27470 10498
rect 27522 10446 27524 10498
rect 26908 9828 26964 9838
rect 26796 9772 26908 9828
rect 26908 9604 26964 9772
rect 26908 9538 26964 9548
rect 27132 9716 27188 9726
rect 26236 9266 26740 9268
rect 26236 9214 26238 9266
rect 26290 9214 26686 9266
rect 26738 9214 26740 9266
rect 26236 9212 26740 9214
rect 26236 9202 26292 9212
rect 25452 8372 25956 8428
rect 25452 8370 25508 8372
rect 25452 8318 25454 8370
rect 25506 8318 25508 8370
rect 25452 8306 25508 8318
rect 25676 8036 25732 8046
rect 25676 7586 25732 7980
rect 25900 8036 25956 8372
rect 26012 8372 26068 8382
rect 26012 8258 26068 8316
rect 26012 8206 26014 8258
rect 26066 8206 26068 8258
rect 26012 8194 26068 8206
rect 26236 8146 26292 8158
rect 26236 8094 26238 8146
rect 26290 8094 26292 8146
rect 26236 8036 26292 8094
rect 25900 7980 26292 8036
rect 26348 8034 26404 8046
rect 26348 7982 26350 8034
rect 26402 7982 26404 8034
rect 25676 7534 25678 7586
rect 25730 7534 25732 7586
rect 25676 7522 25732 7534
rect 25788 7588 25844 7598
rect 25788 7494 25844 7532
rect 25788 6692 25844 6702
rect 25788 6598 25844 6636
rect 25452 6468 25508 6478
rect 25452 6374 25508 6412
rect 25900 6020 25956 7980
rect 26012 7476 26068 7486
rect 26348 7476 26404 7982
rect 26012 7474 26404 7476
rect 26012 7422 26014 7474
rect 26066 7422 26404 7474
rect 26012 7420 26404 7422
rect 26012 7410 26068 7420
rect 26460 6692 26516 6702
rect 26348 6690 26516 6692
rect 26348 6638 26462 6690
rect 26514 6638 26516 6690
rect 26348 6636 26516 6638
rect 26348 6468 26404 6636
rect 26460 6626 26516 6636
rect 26572 6692 26628 9212
rect 26684 9202 26740 9212
rect 27132 9266 27188 9660
rect 27468 9604 27524 10446
rect 27692 9716 27748 9726
rect 27692 9622 27748 9660
rect 27468 9510 27524 9548
rect 27132 9214 27134 9266
rect 27186 9214 27188 9266
rect 27132 9202 27188 9214
rect 27580 9044 27636 9054
rect 27580 8950 27636 8988
rect 26684 8258 26740 8270
rect 26684 8206 26686 8258
rect 26738 8206 26740 8258
rect 26684 7700 26740 8206
rect 27804 8258 27860 11004
rect 28028 11172 28084 11182
rect 27916 10498 27972 10510
rect 27916 10446 27918 10498
rect 27970 10446 27972 10498
rect 27916 9604 27972 10446
rect 28028 9828 28084 11116
rect 28924 11172 28980 11182
rect 28924 11078 28980 11116
rect 28476 10498 28532 10510
rect 28476 10446 28478 10498
rect 28530 10446 28532 10498
rect 28028 9826 28196 9828
rect 28028 9774 28030 9826
rect 28082 9774 28196 9826
rect 28028 9772 28196 9774
rect 28028 9762 28084 9772
rect 27916 9538 27972 9548
rect 28140 9044 28196 9772
rect 28476 9716 28532 10446
rect 28812 10498 28868 10510
rect 28812 10446 28814 10498
rect 28866 10446 28868 10498
rect 28588 9940 28644 9950
rect 28588 9846 28644 9884
rect 28532 9660 28644 9716
rect 28476 9584 28532 9660
rect 28140 9042 28308 9044
rect 28140 8990 28142 9042
rect 28194 8990 28308 9042
rect 28140 8988 28308 8990
rect 28140 8978 28196 8988
rect 28140 8820 28196 8830
rect 28140 8726 28196 8764
rect 27804 8206 27806 8258
rect 27858 8206 27860 8258
rect 27132 8146 27188 8158
rect 27132 8094 27134 8146
rect 27186 8094 27188 8146
rect 27132 7812 27188 8094
rect 27244 8036 27300 8046
rect 27244 7942 27300 7980
rect 27132 7746 27188 7756
rect 26684 7634 26740 7644
rect 27468 7700 27524 7710
rect 27468 7606 27524 7644
rect 27692 7700 27748 7710
rect 27356 7588 27412 7598
rect 27244 7532 27356 7588
rect 26796 7362 26852 7374
rect 26796 7310 26798 7362
rect 26850 7310 26852 7362
rect 26796 7252 26852 7310
rect 27244 7252 27300 7532
rect 27356 7494 27412 7532
rect 27580 7588 27636 7598
rect 27692 7588 27748 7644
rect 27580 7586 27748 7588
rect 27580 7534 27582 7586
rect 27634 7534 27748 7586
rect 27580 7532 27748 7534
rect 27580 7522 27636 7532
rect 26796 7186 26852 7196
rect 27020 7196 27300 7252
rect 27804 7252 27860 8206
rect 28252 8258 28308 8988
rect 28476 8818 28532 8830
rect 28476 8766 28478 8818
rect 28530 8766 28532 8818
rect 28476 8372 28532 8766
rect 28588 8484 28644 9660
rect 28700 9604 28756 9614
rect 28700 9380 28756 9548
rect 28812 9380 28868 10446
rect 29036 10276 29092 11900
rect 29260 10836 29316 10846
rect 29708 10836 29764 10846
rect 29820 10836 29876 12908
rect 29932 11172 29988 13470
rect 30044 13188 30100 13198
rect 30156 13188 30212 13804
rect 30044 13186 30212 13188
rect 30044 13134 30046 13186
rect 30098 13134 30212 13186
rect 30044 13132 30212 13134
rect 30044 13122 30100 13132
rect 30156 12852 30212 12862
rect 30156 12758 30212 12796
rect 29932 11106 29988 11116
rect 30044 12740 30100 12750
rect 30044 12178 30100 12684
rect 30492 12516 30548 14478
rect 30604 13412 30660 14702
rect 31052 14642 31108 15708
rect 31388 15540 31444 15578
rect 31388 15474 31444 15484
rect 31052 14590 31054 14642
rect 31106 14590 31108 14642
rect 31052 14578 31108 14590
rect 31388 15316 31444 15326
rect 31388 14642 31444 15260
rect 31388 14590 31390 14642
rect 31442 14590 31444 14642
rect 31388 14578 31444 14590
rect 31500 14532 31556 17388
rect 31612 15426 31668 15438
rect 31612 15374 31614 15426
rect 31666 15374 31668 15426
rect 31612 14754 31668 15374
rect 31612 14702 31614 14754
rect 31666 14702 31668 14754
rect 31612 14690 31668 14702
rect 31724 15314 31780 17388
rect 31836 17220 31892 18172
rect 31836 17106 31892 17164
rect 31836 17054 31838 17106
rect 31890 17054 31892 17106
rect 31836 16210 31892 17054
rect 31836 16158 31838 16210
rect 31890 16158 31892 16210
rect 31836 16146 31892 16158
rect 32172 16212 32228 18508
rect 32284 18450 32340 19964
rect 32396 21980 32564 22036
rect 32396 19348 32452 21980
rect 32844 21924 32900 22428
rect 33516 22372 33572 22382
rect 32508 21868 32900 21924
rect 32956 22370 33572 22372
rect 32956 22318 33518 22370
rect 33570 22318 33572 22370
rect 32956 22316 33572 22318
rect 32508 21698 32564 21868
rect 32508 21646 32510 21698
rect 32562 21646 32564 21698
rect 32508 21634 32564 21646
rect 32508 20916 32564 20926
rect 32508 20802 32564 20860
rect 32508 20750 32510 20802
rect 32562 20750 32564 20802
rect 32508 20738 32564 20750
rect 32508 19796 32564 19806
rect 32508 19702 32564 19740
rect 32620 19572 32676 21868
rect 32956 21812 33012 22316
rect 33516 22306 33572 22316
rect 32844 21756 33012 21812
rect 33068 22148 33124 22158
rect 33628 22148 33684 22988
rect 33964 22978 34020 22988
rect 32732 21700 32788 21710
rect 32732 21606 32788 21644
rect 32844 21474 32900 21756
rect 32844 21422 32846 21474
rect 32898 21422 32900 21474
rect 32844 21410 32900 21422
rect 32956 21588 33012 21598
rect 32956 20802 33012 21532
rect 32956 20750 32958 20802
rect 33010 20750 33012 20802
rect 32732 20244 32788 20254
rect 32732 20130 32788 20188
rect 32732 20078 32734 20130
rect 32786 20078 32788 20130
rect 32732 20066 32788 20078
rect 32956 20132 33012 20750
rect 32844 20020 32900 20030
rect 32844 19906 32900 19964
rect 32844 19854 32846 19906
rect 32898 19854 32900 19906
rect 32844 19842 32900 19854
rect 32396 19282 32452 19292
rect 32508 19516 32676 19572
rect 32508 19236 32564 19516
rect 32956 19346 33012 20076
rect 32956 19294 32958 19346
rect 33010 19294 33012 19346
rect 32956 19282 33012 19294
rect 32620 19236 32676 19246
rect 32508 19234 32676 19236
rect 32508 19182 32622 19234
rect 32674 19182 32676 19234
rect 32508 19180 32676 19182
rect 32620 19170 32676 19180
rect 33068 19124 33124 22092
rect 33516 22092 33684 22148
rect 33740 22820 33796 22830
rect 32284 18398 32286 18450
rect 32338 18398 32340 18450
rect 32284 18228 32340 18398
rect 32844 19068 33124 19124
rect 33292 21924 33348 21934
rect 32732 18340 32788 18350
rect 32732 18246 32788 18284
rect 32284 18162 32340 18172
rect 32284 17668 32340 17678
rect 32284 17554 32340 17612
rect 32284 17502 32286 17554
rect 32338 17502 32340 17554
rect 32284 17490 32340 17502
rect 32620 17668 32676 17678
rect 32620 16994 32676 17612
rect 32732 17556 32788 17566
rect 32732 17462 32788 17500
rect 32732 17108 32788 17118
rect 32844 17108 32900 19068
rect 32732 17106 32900 17108
rect 32732 17054 32734 17106
rect 32786 17054 32900 17106
rect 32732 17052 32900 17054
rect 32732 17042 32788 17052
rect 32620 16942 32622 16994
rect 32674 16942 32676 16994
rect 32284 16212 32340 16222
rect 32172 16210 32340 16212
rect 32172 16158 32286 16210
rect 32338 16158 32340 16210
rect 32172 16156 32340 16158
rect 32172 15764 32228 16156
rect 32284 16146 32340 16156
rect 32396 16212 32452 16222
rect 32172 15698 32228 15708
rect 32284 15540 32340 15550
rect 32396 15540 32452 16156
rect 32284 15538 32452 15540
rect 32284 15486 32286 15538
rect 32338 15486 32452 15538
rect 32284 15484 32452 15486
rect 32284 15474 32340 15484
rect 32620 15428 32676 16942
rect 32732 16212 32788 16222
rect 32732 16118 32788 16156
rect 32844 15988 32900 17052
rect 33068 18900 33124 18910
rect 33068 17890 33124 18844
rect 33068 17838 33070 17890
rect 33122 17838 33124 17890
rect 32956 16884 33012 16894
rect 32956 16790 33012 16828
rect 33068 16212 33124 17838
rect 33292 18340 33348 21868
rect 33404 20468 33460 20478
rect 33404 19346 33460 20412
rect 33516 20244 33572 22092
rect 33740 21924 33796 22764
rect 33852 22372 33908 22382
rect 33852 22278 33908 22316
rect 33964 22372 34020 22382
rect 34076 22372 34132 23660
rect 34188 22932 34244 24668
rect 34188 22866 34244 22876
rect 33964 22370 34132 22372
rect 33964 22318 33966 22370
rect 34018 22318 34132 22370
rect 33964 22316 34132 22318
rect 33964 22306 34020 22316
rect 34076 22146 34132 22158
rect 34076 22094 34078 22146
rect 34130 22094 34132 22146
rect 33740 21868 33908 21924
rect 33740 21700 33796 21710
rect 33516 20178 33572 20188
rect 33628 20804 33684 20814
rect 33404 19294 33406 19346
rect 33458 19294 33460 19346
rect 33404 19282 33460 19294
rect 33516 18676 33572 18686
rect 33516 18582 33572 18620
rect 33628 18452 33684 20748
rect 33628 18386 33684 18396
rect 33068 16146 33124 16156
rect 33180 17556 33236 17566
rect 33180 16996 33236 17500
rect 33180 16210 33236 16940
rect 33180 16158 33182 16210
rect 33234 16158 33236 16210
rect 32844 15922 32900 15932
rect 32620 15362 32676 15372
rect 31724 15262 31726 15314
rect 31778 15262 31780 15314
rect 31724 15092 31780 15262
rect 31500 14466 31556 14476
rect 31724 14308 31780 15036
rect 32172 15316 32228 15326
rect 31836 14308 31892 14318
rect 31724 14306 31892 14308
rect 31724 14254 31838 14306
rect 31890 14254 31892 14306
rect 31724 14252 31892 14254
rect 31500 13972 31556 13982
rect 31500 13878 31556 13916
rect 30828 13860 30884 13870
rect 30828 13766 30884 13804
rect 31164 13748 31220 13758
rect 30940 13522 30996 13534
rect 30940 13470 30942 13522
rect 30994 13470 30996 13522
rect 30940 13412 30996 13470
rect 30604 13356 30996 13412
rect 30716 12852 30772 12862
rect 30716 12758 30772 12796
rect 30268 12460 30548 12516
rect 30044 12126 30046 12178
rect 30098 12126 30100 12178
rect 29260 10834 29988 10836
rect 29260 10782 29262 10834
rect 29314 10782 29710 10834
rect 29762 10782 29988 10834
rect 29260 10780 29988 10782
rect 29260 10770 29316 10780
rect 29708 10770 29764 10780
rect 29036 10220 29764 10276
rect 29708 10050 29764 10220
rect 29708 9998 29710 10050
rect 29762 9998 29764 10050
rect 29708 9986 29764 9998
rect 29596 9940 29652 9950
rect 29596 9826 29652 9884
rect 29596 9774 29598 9826
rect 29650 9774 29652 9826
rect 29596 9762 29652 9774
rect 29708 9604 29764 9614
rect 29708 9510 29764 9548
rect 28700 9324 28980 9380
rect 28588 8418 28644 8428
rect 28476 8306 28532 8316
rect 28252 8206 28254 8258
rect 28306 8206 28308 8258
rect 28252 7588 28308 8206
rect 28812 8148 28868 8158
rect 28252 7456 28308 7532
rect 28588 8092 28812 8148
rect 27804 7196 28084 7252
rect 27020 6802 27076 7196
rect 27020 6750 27022 6802
rect 27074 6750 27076 6802
rect 27020 6738 27076 6750
rect 26684 6692 26740 6702
rect 26572 6690 26740 6692
rect 26572 6638 26686 6690
rect 26738 6638 26740 6690
rect 26572 6636 26740 6638
rect 26012 6132 26068 6142
rect 26012 6038 26068 6076
rect 25900 5954 25956 5964
rect 26348 5796 26404 6412
rect 26572 6132 26628 6636
rect 26684 6626 26740 6636
rect 26572 6066 26628 6076
rect 27020 6580 27076 6590
rect 27020 6130 27076 6524
rect 27580 6580 27636 6590
rect 27580 6486 27636 6524
rect 27020 6078 27022 6130
rect 27074 6078 27076 6130
rect 26460 6020 26516 6030
rect 26460 5926 26516 5964
rect 26348 5740 26516 5796
rect 26236 5684 26292 5694
rect 25900 5460 25956 5470
rect 25228 5234 25396 5236
rect 25228 5182 25230 5234
rect 25282 5182 25396 5234
rect 25228 5180 25396 5182
rect 25228 5170 25284 5180
rect 24668 4564 24724 4956
rect 24668 4498 24724 4508
rect 25004 4900 25060 4910
rect 25340 4900 25396 5180
rect 25452 5124 25508 5134
rect 25452 5030 25508 5068
rect 25340 4844 25620 4900
rect 25004 4562 25060 4844
rect 25004 4510 25006 4562
rect 25058 4510 25060 4562
rect 25004 4498 25060 4510
rect 23548 4398 23550 4450
rect 23602 4398 23604 4450
rect 23548 4386 23604 4398
rect 25564 4338 25620 4844
rect 25788 4564 25844 4574
rect 25788 4470 25844 4508
rect 25564 4286 25566 4338
rect 25618 4286 25620 4338
rect 25452 3778 25508 3790
rect 25452 3726 25454 3778
rect 25506 3726 25508 3778
rect 23772 3668 23828 3678
rect 23324 3666 23828 3668
rect 23324 3614 23326 3666
rect 23378 3614 23774 3666
rect 23826 3614 23828 3666
rect 23324 3612 23828 3614
rect 23324 3602 23380 3612
rect 23772 3602 23828 3612
rect 24220 3668 24276 3678
rect 24220 3574 24276 3612
rect 24668 3668 24724 3678
rect 24668 3574 24724 3612
rect 25452 3666 25508 3726
rect 25452 3614 25454 3666
rect 25506 3614 25508 3666
rect 25452 3602 25508 3614
rect 25564 3668 25620 4286
rect 25564 3602 25620 3612
rect 25900 3778 25956 5404
rect 26012 5124 26068 5134
rect 26012 4450 26068 5068
rect 26012 4398 26014 4450
rect 26066 4398 26068 4450
rect 26012 4386 26068 4398
rect 26236 4450 26292 5628
rect 26348 5460 26404 5470
rect 26348 5234 26404 5404
rect 26348 5182 26350 5234
rect 26402 5182 26404 5234
rect 26348 5170 26404 5182
rect 26236 4398 26238 4450
rect 26290 4398 26292 4450
rect 26236 4386 26292 4398
rect 26460 4340 26516 5740
rect 26908 5684 26964 5694
rect 26908 5346 26964 5628
rect 27020 5460 27076 6078
rect 27692 5794 27748 5806
rect 27692 5742 27694 5794
rect 27746 5742 27748 5794
rect 27580 5684 27636 5694
rect 27580 5590 27636 5628
rect 27020 5394 27076 5404
rect 27468 5460 27524 5470
rect 26908 5294 26910 5346
rect 26962 5294 26964 5346
rect 26908 5282 26964 5294
rect 27132 5348 27188 5358
rect 26460 4274 26516 4284
rect 26796 4340 26852 4350
rect 25900 3726 25902 3778
rect 25954 3726 25956 3778
rect 25900 3666 25956 3726
rect 25900 3614 25902 3666
rect 25954 3614 25956 3666
rect 25900 3602 25956 3614
rect 26348 4116 26404 4126
rect 26348 3666 26404 4060
rect 26348 3614 26350 3666
rect 26402 3614 26404 3666
rect 26348 3602 26404 3614
rect 26796 3666 26852 4284
rect 26908 4228 26964 4238
rect 26908 4134 26964 4172
rect 27132 4116 27188 5292
rect 27468 5122 27524 5404
rect 27468 5070 27470 5122
rect 27522 5070 27524 5122
rect 27468 5058 27524 5070
rect 27692 5124 27748 5742
rect 27804 5348 27860 7196
rect 28028 6802 28084 7196
rect 28588 6916 28644 8092
rect 28812 8054 28868 8092
rect 28924 8036 28980 9324
rect 29932 9044 29988 10780
rect 30044 10500 30100 12126
rect 30156 12292 30212 12302
rect 30156 11394 30212 12236
rect 30268 11508 30324 12460
rect 30492 12292 30548 12302
rect 30492 12198 30548 12236
rect 30828 12180 30884 13356
rect 31164 13074 31220 13692
rect 31164 13022 31166 13074
rect 31218 13022 31220 13074
rect 31164 13010 31220 13022
rect 31500 13748 31556 13758
rect 31388 12962 31444 12974
rect 31388 12910 31390 12962
rect 31442 12910 31444 12962
rect 30940 12850 30996 12862
rect 30940 12798 30942 12850
rect 30994 12798 30996 12850
rect 30940 12404 30996 12798
rect 30940 12338 30996 12348
rect 31052 12290 31108 12302
rect 31052 12238 31054 12290
rect 31106 12238 31108 12290
rect 31052 12180 31108 12238
rect 30828 12124 30996 12180
rect 30268 11442 30324 11452
rect 30380 12068 30436 12078
rect 30156 11342 30158 11394
rect 30210 11342 30212 11394
rect 30156 11330 30212 11342
rect 30156 10500 30212 10510
rect 30044 10498 30212 10500
rect 30044 10446 30158 10498
rect 30210 10446 30212 10498
rect 30044 10444 30212 10446
rect 30156 10388 30212 10444
rect 30156 10322 30212 10332
rect 30268 9604 30324 9614
rect 30044 9044 30100 9054
rect 29988 9042 30100 9044
rect 29988 8990 30046 9042
rect 30098 8990 30100 9042
rect 29988 8988 30100 8990
rect 29148 8932 29204 8942
rect 29148 8838 29204 8876
rect 29820 8930 29876 8942
rect 29820 8878 29822 8930
rect 29874 8878 29876 8930
rect 29932 8912 29988 8988
rect 28924 7970 28980 7980
rect 29036 8484 29092 8494
rect 28812 7474 28868 7486
rect 28812 7422 28814 7474
rect 28866 7422 28868 7474
rect 28812 7252 28868 7422
rect 28812 7186 28868 7196
rect 28028 6750 28030 6802
rect 28082 6750 28084 6802
rect 28028 6692 28084 6750
rect 28028 6626 28084 6636
rect 28476 6860 28644 6916
rect 28476 6468 28532 6860
rect 28588 6692 28644 6702
rect 28588 6598 28644 6636
rect 28700 6578 28756 6590
rect 28700 6526 28702 6578
rect 28754 6526 28756 6578
rect 28476 6412 28644 6468
rect 28588 6130 28644 6412
rect 28588 6078 28590 6130
rect 28642 6078 28644 6130
rect 28588 6066 28644 6078
rect 27916 5908 27972 5918
rect 27916 5906 28420 5908
rect 27916 5854 27918 5906
rect 27970 5854 28420 5906
rect 27916 5852 28420 5854
rect 27916 5842 27972 5852
rect 27804 5282 27860 5292
rect 28364 5234 28420 5852
rect 28364 5182 28366 5234
rect 28418 5182 28420 5234
rect 28364 5170 28420 5182
rect 28476 5460 28532 5470
rect 27692 5058 27748 5068
rect 28140 5122 28196 5134
rect 28140 5070 28142 5122
rect 28194 5070 28196 5122
rect 27356 5010 27412 5022
rect 27356 4958 27358 5010
rect 27410 4958 27412 5010
rect 27356 4452 27412 4958
rect 27580 5010 27636 5022
rect 27580 4958 27582 5010
rect 27634 4958 27636 5010
rect 27580 4900 27636 4958
rect 27580 4834 27636 4844
rect 28028 4452 28084 4462
rect 28140 4452 28196 5070
rect 28476 5122 28532 5404
rect 28476 5070 28478 5122
rect 28530 5070 28532 5122
rect 28476 5058 28532 5070
rect 27356 4450 28196 4452
rect 27356 4398 28030 4450
rect 28082 4398 28196 4450
rect 27356 4396 28196 4398
rect 28252 4788 28308 4798
rect 27244 4340 27300 4350
rect 27356 4340 27412 4396
rect 28028 4386 28084 4396
rect 27244 4338 27412 4340
rect 27244 4286 27246 4338
rect 27298 4286 27412 4338
rect 27244 4284 27412 4286
rect 27244 4274 27300 4284
rect 27468 4226 27524 4238
rect 27468 4174 27470 4226
rect 27522 4174 27524 4226
rect 27468 4116 27524 4174
rect 27132 4060 27524 4116
rect 28140 4228 28196 4238
rect 28252 4228 28308 4732
rect 28476 4452 28532 4462
rect 28364 4340 28420 4350
rect 28364 4246 28420 4284
rect 28476 4338 28532 4396
rect 28476 4286 28478 4338
rect 28530 4286 28532 4338
rect 28196 4172 28308 4228
rect 28140 4096 28196 4172
rect 26796 3614 26798 3666
rect 26850 3614 26852 3666
rect 26796 3602 26852 3614
rect 27692 3778 27748 3790
rect 27692 3726 27694 3778
rect 27746 3726 27748 3778
rect 27692 3666 27748 3726
rect 28476 3778 28532 4286
rect 28476 3726 28478 3778
rect 28530 3726 28532 3778
rect 28476 3714 28532 3726
rect 28588 4450 28644 4462
rect 28588 4398 28590 4450
rect 28642 4398 28644 4450
rect 27692 3614 27694 3666
rect 27746 3614 27748 3666
rect 27692 3602 27748 3614
rect 28588 3666 28644 4398
rect 28588 3614 28590 3666
rect 28642 3614 28644 3666
rect 28588 3602 28644 3614
rect 21644 3502 21646 3554
rect 21698 3502 21700 3554
rect 21644 3490 21700 3502
rect 28140 3556 28196 3566
rect 21532 3390 21534 3442
rect 21586 3390 21588 3442
rect 21532 3378 21588 3390
rect 27244 3444 27300 3482
rect 28140 3462 28196 3500
rect 28700 3556 28756 6526
rect 29036 6018 29092 8428
rect 29708 8484 29764 8494
rect 29820 8484 29876 8878
rect 29708 8482 29876 8484
rect 29708 8430 29710 8482
rect 29762 8430 29876 8482
rect 29708 8428 29876 8430
rect 29932 8484 29988 8494
rect 29708 8372 29764 8428
rect 29708 8306 29764 8316
rect 29820 8260 29876 8270
rect 29932 8260 29988 8428
rect 29820 8258 29988 8260
rect 29820 8206 29822 8258
rect 29874 8206 29988 8258
rect 29820 8204 29988 8206
rect 29820 8194 29876 8204
rect 29708 8036 29764 8046
rect 29708 7942 29764 7980
rect 29820 7700 29876 7710
rect 29820 7474 29876 7644
rect 29820 7422 29822 7474
rect 29874 7422 29876 7474
rect 29820 7410 29876 7422
rect 29932 7252 29988 7262
rect 30044 7252 30100 8988
rect 30268 9042 30324 9548
rect 30268 8990 30270 9042
rect 30322 8990 30324 9042
rect 30268 8372 30324 8990
rect 30268 8306 30324 8316
rect 30268 8034 30324 8046
rect 30268 7982 30270 8034
rect 30322 7982 30324 8034
rect 30268 7700 30324 7982
rect 30268 7634 30324 7644
rect 30380 7476 30436 12012
rect 30604 11620 30660 11630
rect 30604 11506 30660 11564
rect 30604 11454 30606 11506
rect 30658 11454 30660 11506
rect 30604 11442 30660 11454
rect 30828 11508 30884 11518
rect 30492 11396 30548 11406
rect 30492 11302 30548 11340
rect 30716 10498 30772 10510
rect 30716 10446 30718 10498
rect 30770 10446 30772 10498
rect 30716 9604 30772 10446
rect 30716 9538 30772 9548
rect 30604 8146 30660 8158
rect 30604 8094 30606 8146
rect 30658 8094 30660 8146
rect 30380 7410 30436 7420
rect 30492 8036 30548 8046
rect 30268 7364 30324 7374
rect 30268 7270 30324 7308
rect 29932 7250 30100 7252
rect 29932 7198 29934 7250
rect 29986 7198 30100 7250
rect 29932 7196 30100 7198
rect 30156 7252 30212 7262
rect 29596 6580 29652 6590
rect 29036 5966 29038 6018
rect 29090 5966 29092 6018
rect 28924 5124 28980 5134
rect 28812 5010 28868 5022
rect 28812 4958 28814 5010
rect 28866 4958 28868 5010
rect 28812 4900 28868 4958
rect 28812 4834 28868 4844
rect 28924 4450 28980 5068
rect 28924 4398 28926 4450
rect 28978 4398 28980 4450
rect 28924 4386 28980 4398
rect 29036 4340 29092 5966
rect 29372 6356 29428 6366
rect 29372 6132 29428 6300
rect 29372 6018 29428 6076
rect 29372 5966 29374 6018
rect 29426 5966 29428 6018
rect 29372 5954 29428 5966
rect 29036 4274 29092 4284
rect 29260 4338 29316 4350
rect 29260 4286 29262 4338
rect 29314 4286 29316 4338
rect 28700 3490 28756 3500
rect 29260 3556 29316 4286
rect 29596 4226 29652 6524
rect 29932 6580 29988 7196
rect 29932 6514 29988 6524
rect 29820 6466 29876 6478
rect 29820 6414 29822 6466
rect 29874 6414 29876 6466
rect 29708 6356 29764 6366
rect 29708 5124 29764 6300
rect 29708 4992 29764 5068
rect 29820 6356 29876 6414
rect 30156 6356 30212 7196
rect 30268 6468 30324 6478
rect 30492 6468 30548 7980
rect 30268 6466 30548 6468
rect 30268 6414 30270 6466
rect 30322 6414 30548 6466
rect 30268 6412 30548 6414
rect 30604 6804 30660 8094
rect 30716 6804 30772 6814
rect 30604 6802 30772 6804
rect 30604 6750 30718 6802
rect 30770 6750 30772 6802
rect 30604 6748 30772 6750
rect 30268 6402 30324 6412
rect 29820 6300 30212 6356
rect 29820 4452 29876 6300
rect 30268 5794 30324 5806
rect 30268 5742 30270 5794
rect 30322 5742 30324 5794
rect 30268 5572 30324 5742
rect 30268 5506 30324 5516
rect 30380 5010 30436 6412
rect 30604 6356 30660 6748
rect 30716 6738 30772 6748
rect 30604 6290 30660 6300
rect 30604 6132 30660 6142
rect 30604 6038 30660 6076
rect 30828 6130 30884 11452
rect 30940 9714 30996 12124
rect 31052 12114 31108 12124
rect 31276 12178 31332 12190
rect 31276 12126 31278 12178
rect 31330 12126 31332 12178
rect 31276 11620 31332 12126
rect 31276 11554 31332 11564
rect 31388 11396 31444 12910
rect 30940 9662 30942 9714
rect 30994 9662 30996 9714
rect 30940 9650 30996 9662
rect 31052 11284 31108 11294
rect 31052 11170 31108 11228
rect 31052 11118 31054 11170
rect 31106 11118 31108 11170
rect 31052 9492 31108 11118
rect 31388 10836 31444 11340
rect 31500 11284 31556 13692
rect 31724 13524 31780 14252
rect 31836 14242 31892 14252
rect 32172 13748 32228 15260
rect 32620 15204 32676 15214
rect 33180 15204 33236 16158
rect 32620 15202 33236 15204
rect 32620 15150 32622 15202
rect 32674 15150 33236 15202
rect 32620 15148 33236 15150
rect 32620 15138 32676 15148
rect 32508 15092 32564 15102
rect 31724 13074 31780 13468
rect 31724 13022 31726 13074
rect 31778 13022 31780 13074
rect 31724 13010 31780 13022
rect 32060 13746 32228 13748
rect 32060 13694 32174 13746
rect 32226 13694 32228 13746
rect 32060 13692 32228 13694
rect 31948 12404 32004 12414
rect 32060 12404 32116 13692
rect 32172 13682 32228 13692
rect 32284 14532 32340 14542
rect 32172 13076 32228 13086
rect 32284 13076 32340 14476
rect 32508 14530 32564 15036
rect 33068 15092 33236 15148
rect 33292 15148 33348 18284
rect 33404 17668 33460 17678
rect 33404 17574 33460 17612
rect 33740 16882 33796 21644
rect 33852 21586 33908 21868
rect 33852 21534 33854 21586
rect 33906 21534 33908 21586
rect 33852 20580 33908 21534
rect 33852 20514 33908 20524
rect 33964 21474 34020 21486
rect 33964 21422 33966 21474
rect 34018 21422 34020 21474
rect 33852 20132 33908 20142
rect 33852 20018 33908 20076
rect 33852 19966 33854 20018
rect 33906 19966 33908 20018
rect 33852 19954 33908 19966
rect 33852 19458 33908 19470
rect 33852 19406 33854 19458
rect 33906 19406 33908 19458
rect 33852 19346 33908 19406
rect 33852 19294 33854 19346
rect 33906 19294 33908 19346
rect 33852 19282 33908 19294
rect 33964 19348 34020 21422
rect 34076 21364 34132 22094
rect 34188 22146 34244 22158
rect 34188 22094 34190 22146
rect 34242 22094 34244 22146
rect 34188 21700 34244 22094
rect 34188 21634 34244 21644
rect 34076 21298 34132 21308
rect 34188 21028 34244 21038
rect 34300 21028 34356 25116
rect 34244 20972 34356 21028
rect 34412 21474 34468 26908
rect 34636 26516 34692 26526
rect 34524 24722 34580 24734
rect 34524 24670 34526 24722
rect 34578 24670 34580 24722
rect 34524 24612 34580 24670
rect 34524 22596 34580 24556
rect 34636 23716 34692 26460
rect 34860 26068 34916 29262
rect 34972 26908 35028 29372
rect 35084 29426 35140 29708
rect 35084 29374 35086 29426
rect 35138 29374 35140 29426
rect 35084 29204 35140 29374
rect 35196 29428 35252 30380
rect 35196 29362 35252 29372
rect 35420 29876 35476 29886
rect 35084 29138 35140 29148
rect 35420 29204 35476 29820
rect 35420 29138 35476 29148
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35084 28642 35140 28654
rect 35084 28590 35086 28642
rect 35138 28590 35140 28642
rect 35084 28532 35140 28590
rect 35084 27972 35140 28476
rect 35084 27916 35252 27972
rect 35196 27860 35252 27916
rect 35420 27860 35476 27870
rect 35196 27858 35476 27860
rect 35196 27806 35422 27858
rect 35474 27806 35476 27858
rect 35196 27804 35476 27806
rect 35532 27860 35588 30380
rect 35644 28308 35700 30716
rect 35756 29652 35812 32956
rect 36316 32452 36372 32462
rect 36092 32340 36148 32350
rect 35868 31668 35924 31678
rect 35868 31574 35924 31612
rect 36092 31444 36148 32284
rect 35980 31220 36036 31230
rect 36092 31220 36148 31388
rect 35980 31218 36148 31220
rect 35980 31166 35982 31218
rect 36034 31166 36148 31218
rect 35980 31164 36148 31166
rect 35980 31154 36036 31164
rect 35868 30996 35924 31006
rect 35868 30210 35924 30940
rect 36204 30772 36260 30782
rect 35868 30158 35870 30210
rect 35922 30158 35924 30210
rect 35868 30146 35924 30158
rect 36092 30212 36148 30222
rect 36092 30118 36148 30156
rect 36204 30210 36260 30716
rect 36204 30158 36206 30210
rect 36258 30158 36260 30210
rect 36204 30146 36260 30158
rect 35980 29986 36036 29998
rect 35980 29934 35982 29986
rect 36034 29934 36036 29986
rect 35980 29876 36036 29934
rect 35980 29810 36036 29820
rect 36316 29764 36372 32396
rect 36428 32340 36484 32350
rect 36428 32338 36820 32340
rect 36428 32286 36430 32338
rect 36482 32286 36820 32338
rect 36428 32284 36820 32286
rect 36428 32274 36484 32284
rect 36428 31778 36484 31790
rect 36428 31726 36430 31778
rect 36482 31726 36484 31778
rect 36428 31108 36484 31726
rect 36428 31042 36484 31052
rect 36540 31556 36596 31566
rect 36316 29708 36484 29764
rect 35868 29652 35924 29662
rect 35756 29650 36372 29652
rect 35756 29598 35870 29650
rect 35922 29598 36372 29650
rect 35756 29596 36372 29598
rect 35868 29586 35924 29596
rect 35756 29428 35812 29438
rect 36092 29428 36148 29438
rect 35812 29372 35924 29428
rect 35756 29296 35812 29372
rect 35868 28756 35924 29372
rect 36092 29426 36260 29428
rect 36092 29374 36094 29426
rect 36146 29374 36260 29426
rect 36092 29372 36260 29374
rect 36092 29362 36148 29372
rect 35868 28662 35924 28700
rect 36092 29204 36148 29214
rect 35756 28644 35812 28654
rect 35756 28420 35812 28588
rect 35980 28644 36036 28654
rect 35980 28550 36036 28588
rect 36092 28532 36148 29148
rect 35756 28364 36036 28420
rect 36092 28400 36148 28476
rect 35644 28252 35924 28308
rect 35644 27860 35700 27870
rect 35532 27858 35700 27860
rect 35532 27806 35646 27858
rect 35698 27806 35700 27858
rect 35532 27804 35700 27806
rect 35420 27794 35476 27804
rect 35644 27794 35700 27804
rect 35644 27524 35700 27534
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35308 27300 35364 27310
rect 34972 26852 35140 26908
rect 34972 26740 35028 26750
rect 34972 26402 35028 26684
rect 34972 26350 34974 26402
rect 35026 26350 35028 26402
rect 34972 26180 35028 26350
rect 34972 26114 35028 26124
rect 34860 26002 34916 26012
rect 34748 25620 34804 25630
rect 34748 25172 34804 25564
rect 34860 25396 34916 25406
rect 34860 25394 35028 25396
rect 34860 25342 34862 25394
rect 34914 25342 35028 25394
rect 34860 25340 35028 25342
rect 34860 25330 34916 25340
rect 34748 25116 34916 25172
rect 34636 23650 34692 23660
rect 34748 24946 34804 24958
rect 34748 24894 34750 24946
rect 34802 24894 34804 24946
rect 34748 24050 34804 24894
rect 34860 24946 34916 25116
rect 34860 24894 34862 24946
rect 34914 24894 34916 24946
rect 34860 24836 34916 24894
rect 34860 24770 34916 24780
rect 34972 24724 35028 25340
rect 35084 25172 35140 26852
rect 35196 26516 35252 26526
rect 35196 26422 35252 26460
rect 35308 26514 35364 27244
rect 35308 26462 35310 26514
rect 35362 26462 35364 26514
rect 35308 26450 35364 26462
rect 35532 26852 35588 26862
rect 35420 26292 35476 26302
rect 35420 26198 35476 26236
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35532 25394 35588 26796
rect 35532 25342 35534 25394
rect 35586 25342 35588 25394
rect 35084 25106 35140 25116
rect 35308 25284 35364 25294
rect 35308 24724 35364 25228
rect 34972 24658 35028 24668
rect 35084 24668 35364 24724
rect 34748 23998 34750 24050
rect 34802 23998 34804 24050
rect 34748 23604 34804 23998
rect 34636 23156 34692 23166
rect 34636 23062 34692 23100
rect 34748 23154 34804 23548
rect 34748 23102 34750 23154
rect 34802 23102 34804 23154
rect 34748 23090 34804 23102
rect 34972 23828 35028 23838
rect 35084 23828 35140 24668
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 34972 23826 35140 23828
rect 34972 23774 34974 23826
rect 35026 23774 35140 23826
rect 34972 23772 35140 23774
rect 34972 23044 35028 23772
rect 35196 23492 35252 23502
rect 35084 23268 35140 23278
rect 35084 23174 35140 23212
rect 35196 23044 35252 23436
rect 35532 23492 35588 25342
rect 35644 24948 35700 27468
rect 35868 26178 35924 28252
rect 35868 26126 35870 26178
rect 35922 26126 35924 26178
rect 35868 25844 35924 26126
rect 35980 26066 36036 28364
rect 36204 27074 36260 29372
rect 36316 28868 36372 29596
rect 36428 29650 36484 29708
rect 36428 29598 36430 29650
rect 36482 29598 36484 29650
rect 36428 29586 36484 29598
rect 36428 28868 36484 28878
rect 36316 28866 36484 28868
rect 36316 28814 36430 28866
rect 36482 28814 36484 28866
rect 36316 28812 36484 28814
rect 36428 28802 36484 28812
rect 36316 28084 36372 28094
rect 36316 27970 36372 28028
rect 36316 27918 36318 27970
rect 36370 27918 36372 27970
rect 36316 27906 36372 27918
rect 36540 27636 36596 31500
rect 36764 30996 36820 32284
rect 36876 31668 36932 32956
rect 36988 32564 37044 32574
rect 36988 32470 37044 32508
rect 36876 31602 36932 31612
rect 36652 30884 36708 30894
rect 36764 30864 36820 30940
rect 36876 31108 36932 31118
rect 36652 30212 36708 30828
rect 36764 30212 36820 30222
rect 36652 30210 36820 30212
rect 36652 30158 36766 30210
rect 36818 30158 36820 30210
rect 36652 30156 36820 30158
rect 36764 30146 36820 30156
rect 36652 28866 36708 28878
rect 36652 28814 36654 28866
rect 36706 28814 36708 28866
rect 36652 28754 36708 28814
rect 36652 28702 36654 28754
rect 36706 28702 36708 28754
rect 36652 27972 36708 28702
rect 36652 27906 36708 27916
rect 36764 28084 36820 28094
rect 36204 27022 36206 27074
rect 36258 27022 36260 27074
rect 36204 27010 36260 27022
rect 36316 27580 36596 27636
rect 36316 27074 36372 27580
rect 36316 27022 36318 27074
rect 36370 27022 36372 27074
rect 36316 27010 36372 27022
rect 36540 27412 36596 27422
rect 36540 27074 36596 27356
rect 36540 27022 36542 27074
rect 36594 27022 36596 27074
rect 36540 27010 36596 27022
rect 36652 26962 36708 26974
rect 36652 26910 36654 26962
rect 36706 26910 36708 26962
rect 36428 26850 36484 26862
rect 36428 26798 36430 26850
rect 36482 26798 36484 26850
rect 36428 26740 36484 26798
rect 35980 26014 35982 26066
rect 36034 26014 36036 26066
rect 35980 26002 36036 26014
rect 36204 26684 36484 26740
rect 36540 26852 36596 26862
rect 35868 25778 35924 25788
rect 35756 25284 35812 25294
rect 35756 25190 35812 25228
rect 35868 25282 35924 25294
rect 35868 25230 35870 25282
rect 35922 25230 35924 25282
rect 35644 24892 35812 24948
rect 35532 23156 35588 23436
rect 35644 24722 35700 24734
rect 35644 24670 35646 24722
rect 35698 24670 35700 24722
rect 35644 23268 35700 24670
rect 35644 23202 35700 23212
rect 35532 23090 35588 23100
rect 34636 22932 34692 22942
rect 34692 22876 34804 22932
rect 34636 22866 34692 22876
rect 34524 22540 34692 22596
rect 34636 21924 34692 22540
rect 34748 22484 34804 22876
rect 34972 22930 35028 22988
rect 34972 22878 34974 22930
rect 35026 22878 35028 22930
rect 34860 22484 34916 22494
rect 34748 22482 34916 22484
rect 34748 22430 34862 22482
rect 34914 22430 34916 22482
rect 34748 22428 34916 22430
rect 34860 22418 34916 22428
rect 34972 21924 35028 22878
rect 35084 22988 35252 23044
rect 35644 23044 35700 23054
rect 35084 22148 35140 22988
rect 35644 22950 35700 22988
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35644 22484 35700 22494
rect 35196 22148 35252 22158
rect 35084 22092 35196 22148
rect 35196 22054 35252 22092
rect 35644 22036 35700 22428
rect 35644 21970 35700 21980
rect 34636 21868 34916 21924
rect 34860 21810 34916 21868
rect 34972 21858 35028 21868
rect 35308 21924 35364 21934
rect 34860 21758 34862 21810
rect 34914 21758 34916 21810
rect 34860 21746 34916 21758
rect 35308 21810 35364 21868
rect 35308 21758 35310 21810
rect 35362 21758 35364 21810
rect 35308 21746 35364 21758
rect 35532 21812 35588 21822
rect 34412 21422 34414 21474
rect 34466 21422 34468 21474
rect 34076 20802 34132 20814
rect 34076 20750 34078 20802
rect 34130 20750 34132 20802
rect 34076 20468 34132 20750
rect 34188 20804 34244 20972
rect 34188 20672 34244 20748
rect 34132 20412 34356 20468
rect 34076 20402 34132 20412
rect 34188 19906 34244 19918
rect 34188 19854 34190 19906
rect 34242 19854 34244 19906
rect 33964 19282 34020 19292
rect 34076 19458 34132 19470
rect 34076 19406 34078 19458
rect 34130 19406 34132 19458
rect 34076 18676 34132 19406
rect 34188 19124 34244 19854
rect 34300 19346 34356 20412
rect 34412 19572 34468 21422
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 34748 21028 34804 21038
rect 34748 20934 34804 20972
rect 34860 20916 34916 20926
rect 34636 20804 34692 20814
rect 34636 20356 34692 20748
rect 34636 19906 34692 20300
rect 34636 19854 34638 19906
rect 34690 19854 34692 19906
rect 34412 19506 34468 19516
rect 34524 19796 34580 19806
rect 34300 19294 34302 19346
rect 34354 19294 34356 19346
rect 34300 19282 34356 19294
rect 34188 19068 34468 19124
rect 34076 18620 34356 18676
rect 34188 18452 34244 18462
rect 34188 18358 34244 18396
rect 33852 17668 33908 17678
rect 33852 17106 33908 17612
rect 34188 17668 34244 17678
rect 34188 17574 34244 17612
rect 33852 17054 33854 17106
rect 33906 17054 33908 17106
rect 33852 17042 33908 17054
rect 33964 17220 34020 17230
rect 33740 16830 33742 16882
rect 33794 16830 33796 16882
rect 33740 16818 33796 16830
rect 33964 16100 34020 17164
rect 34076 17108 34132 17118
rect 34076 17014 34132 17052
rect 34188 16996 34244 17006
rect 34188 16902 34244 16940
rect 34188 16770 34244 16782
rect 34188 16718 34190 16770
rect 34242 16718 34244 16770
rect 34188 16660 34244 16718
rect 34188 16594 34244 16604
rect 34076 16100 34132 16110
rect 33964 16044 34076 16100
rect 33628 15988 33684 15998
rect 34076 15968 34132 16044
rect 34188 15988 34244 15998
rect 33628 15538 33684 15932
rect 34188 15894 34244 15932
rect 33628 15486 33630 15538
rect 33682 15486 33684 15538
rect 33628 15474 33684 15486
rect 33516 15316 33572 15326
rect 33292 15092 33460 15148
rect 32508 14478 32510 14530
rect 32562 14478 32564 14530
rect 32508 13972 32564 14478
rect 32732 14532 32788 14542
rect 32732 14438 32788 14476
rect 32844 14308 32900 14318
rect 32508 13906 32564 13916
rect 32732 14306 32900 14308
rect 32732 14254 32846 14306
rect 32898 14254 32900 14306
rect 32732 14252 32900 14254
rect 32396 13748 32452 13758
rect 32396 13654 32452 13692
rect 32620 13746 32676 13758
rect 32620 13694 32622 13746
rect 32674 13694 32676 13746
rect 32508 13634 32564 13646
rect 32508 13582 32510 13634
rect 32562 13582 32564 13634
rect 32172 13074 32340 13076
rect 32172 13022 32174 13074
rect 32226 13022 32340 13074
rect 32172 13020 32340 13022
rect 32172 13010 32228 13020
rect 31948 12402 32116 12404
rect 31948 12350 31950 12402
rect 32002 12350 32116 12402
rect 31948 12348 32116 12350
rect 31948 12338 32004 12348
rect 32284 11954 32340 13020
rect 32396 13524 32452 13534
rect 32396 12402 32452 13468
rect 32396 12350 32398 12402
rect 32450 12350 32452 12402
rect 32396 12338 32452 12350
rect 32284 11902 32286 11954
rect 32338 11902 32340 11954
rect 32284 11890 32340 11902
rect 31500 11218 31556 11228
rect 32172 11284 32228 11294
rect 31500 10836 31556 10846
rect 31388 10834 31556 10836
rect 31388 10782 31502 10834
rect 31554 10782 31556 10834
rect 31388 10780 31556 10782
rect 31500 10770 31556 10780
rect 32172 10724 32228 11228
rect 32508 11172 32564 13582
rect 32620 13524 32676 13694
rect 32620 13458 32676 13468
rect 32732 13300 32788 14252
rect 32844 14242 32900 14252
rect 32956 14306 33012 14318
rect 32956 14254 32958 14306
rect 33010 14254 33012 14306
rect 32844 13746 32900 13758
rect 32844 13694 32846 13746
rect 32898 13694 32900 13746
rect 32844 13636 32900 13694
rect 32844 13570 32900 13580
rect 32956 13524 33012 14254
rect 32956 13458 33012 13468
rect 33068 14306 33124 15092
rect 33068 14254 33070 14306
rect 33122 14254 33124 14306
rect 32620 13244 32788 13300
rect 32620 11284 32676 13244
rect 32732 13076 32788 13086
rect 33068 13076 33124 14254
rect 32732 13074 33124 13076
rect 32732 13022 32734 13074
rect 32786 13022 33124 13074
rect 32732 13020 33124 13022
rect 32732 13010 32788 13020
rect 32956 12628 33012 12638
rect 32956 12402 33012 12572
rect 32956 12350 32958 12402
rect 33010 12350 33012 12402
rect 32956 12338 33012 12350
rect 32844 11954 32900 11966
rect 32844 11902 32846 11954
rect 32898 11902 32900 11954
rect 32620 11228 32788 11284
rect 32396 11116 32564 11172
rect 32396 10836 32452 11116
rect 32396 10770 32452 10780
rect 32172 10658 32228 10668
rect 32620 10724 32676 10734
rect 32620 10630 32676 10668
rect 31388 10610 31444 10622
rect 31388 10558 31390 10610
rect 31442 10558 31444 10610
rect 31388 9828 31444 10558
rect 31388 9762 31444 9772
rect 31500 10612 31556 10622
rect 31500 9826 31556 10556
rect 31612 10612 31668 10622
rect 31612 10610 31780 10612
rect 31612 10558 31614 10610
rect 31666 10558 31780 10610
rect 31612 10556 31780 10558
rect 31612 10546 31668 10556
rect 31500 9774 31502 9826
rect 31554 9774 31556 9826
rect 30940 9436 31108 9492
rect 30940 8932 30996 9436
rect 31052 9268 31108 9278
rect 31500 9268 31556 9774
rect 31052 9266 31556 9268
rect 31052 9214 31054 9266
rect 31106 9214 31556 9266
rect 31052 9212 31556 9214
rect 31052 9202 31108 9212
rect 31500 8932 31556 9212
rect 31724 9266 31780 10556
rect 32060 10610 32116 10622
rect 32060 10558 32062 10610
rect 32114 10558 32116 10610
rect 32060 10388 32116 10558
rect 32508 10612 32564 10622
rect 32508 10518 32564 10556
rect 32620 10388 32676 10398
rect 32060 10386 32676 10388
rect 32060 10334 32622 10386
rect 32674 10334 32676 10386
rect 32060 10332 32676 10334
rect 32620 10322 32676 10332
rect 32172 9828 32228 9838
rect 32732 9828 32788 11228
rect 32844 11172 32900 11902
rect 33404 11620 33460 15092
rect 33516 12962 33572 15260
rect 33964 15316 34020 15326
rect 33964 15222 34020 15260
rect 34300 15148 34356 18620
rect 34412 18564 34468 19068
rect 34412 18470 34468 18508
rect 34524 17666 34580 19740
rect 34636 18676 34692 19854
rect 34860 20018 34916 20860
rect 35532 20802 35588 21756
rect 35756 21700 35812 24892
rect 35868 24834 35924 25230
rect 35868 24782 35870 24834
rect 35922 24782 35924 24834
rect 35868 24770 35924 24782
rect 35980 25282 36036 25294
rect 35980 25230 35982 25282
rect 36034 25230 36036 25282
rect 35868 23604 35924 23614
rect 35980 23604 36036 25230
rect 36092 25172 36148 25182
rect 36092 24946 36148 25116
rect 36092 24894 36094 24946
rect 36146 24894 36148 24946
rect 36092 24882 36148 24894
rect 36204 24164 36260 26684
rect 36428 26178 36484 26190
rect 36428 26126 36430 26178
rect 36482 26126 36484 26178
rect 36428 26066 36484 26126
rect 36428 26014 36430 26066
rect 36482 26014 36484 26066
rect 36428 26002 36484 26014
rect 36428 25844 36484 25854
rect 36316 24724 36372 24734
rect 36316 24630 36372 24668
rect 36204 24108 36372 24164
rect 35924 23548 36036 23604
rect 36092 24052 36148 24062
rect 36092 23938 36148 23996
rect 36092 23886 36094 23938
rect 36146 23886 36148 23938
rect 35868 23154 35924 23548
rect 35868 23102 35870 23154
rect 35922 23102 35924 23154
rect 35868 23090 35924 23102
rect 36092 22484 36148 23886
rect 36204 23940 36260 23950
rect 36204 23378 36260 23884
rect 36204 23326 36206 23378
rect 36258 23326 36260 23378
rect 36204 23314 36260 23326
rect 36092 22482 36260 22484
rect 36092 22430 36094 22482
rect 36146 22430 36260 22482
rect 36092 22428 36260 22430
rect 36092 22418 36148 22428
rect 35532 20750 35534 20802
rect 35586 20750 35588 20802
rect 35532 20738 35588 20750
rect 35644 21644 35812 21700
rect 36204 21812 36260 22428
rect 36316 21924 36372 24108
rect 36316 21858 36372 21868
rect 36204 21700 36260 21756
rect 36316 21700 36372 21710
rect 36204 21698 36372 21700
rect 36204 21646 36318 21698
rect 36370 21646 36372 21698
rect 36204 21644 36372 21646
rect 35532 20244 35588 20254
rect 34860 19966 34862 20018
rect 34914 19966 34916 20018
rect 34860 19460 34916 19966
rect 35084 20132 35140 20142
rect 34972 19796 35028 19806
rect 34972 19702 35028 19740
rect 34860 19458 35028 19460
rect 34860 19406 34862 19458
rect 34914 19406 35028 19458
rect 34860 19404 35028 19406
rect 34860 19394 34916 19404
rect 34748 19348 34804 19358
rect 34748 19254 34804 19292
rect 34860 19236 34916 19246
rect 34636 18610 34692 18620
rect 34748 18900 34804 18910
rect 34748 18562 34804 18844
rect 34748 18510 34750 18562
rect 34802 18510 34804 18562
rect 34748 18498 34804 18510
rect 34524 17614 34526 17666
rect 34578 17614 34580 17666
rect 34524 17602 34580 17614
rect 34636 18338 34692 18350
rect 34636 18286 34638 18338
rect 34690 18286 34692 18338
rect 34636 17668 34692 18286
rect 34636 17602 34692 17612
rect 34748 18340 34804 18350
rect 34524 17108 34580 17118
rect 34076 15092 34356 15148
rect 34412 15874 34468 15886
rect 34412 15822 34414 15874
rect 34466 15822 34468 15874
rect 33852 14754 33908 14766
rect 33852 14702 33854 14754
rect 33906 14702 33908 14754
rect 33516 12910 33518 12962
rect 33570 12910 33572 12962
rect 33516 12628 33572 12910
rect 33516 12562 33572 12572
rect 33628 14084 33684 14094
rect 33516 12404 33572 12414
rect 33628 12404 33684 14028
rect 33740 13748 33796 13758
rect 33740 13074 33796 13692
rect 33852 13636 33908 14702
rect 34076 14530 34132 15092
rect 34076 14478 34078 14530
rect 34130 14478 34132 14530
rect 34076 14308 34132 14478
rect 33852 13570 33908 13580
rect 33964 14252 34132 14308
rect 33964 13860 34020 14252
rect 33740 13022 33742 13074
rect 33794 13022 33796 13074
rect 33740 13010 33796 13022
rect 33516 12402 33796 12404
rect 33516 12350 33518 12402
rect 33570 12350 33796 12402
rect 33516 12348 33796 12350
rect 33516 12338 33572 12348
rect 33516 11620 33572 11630
rect 32956 11618 33572 11620
rect 32956 11566 33518 11618
rect 33570 11566 33572 11618
rect 32956 11564 33572 11566
rect 32956 11506 33012 11564
rect 32956 11454 32958 11506
rect 33010 11454 33012 11506
rect 32956 11442 33012 11454
rect 32844 11116 33460 11172
rect 32956 10836 33012 10846
rect 32228 9772 32340 9828
rect 32732 9772 32900 9828
rect 32172 9734 32228 9772
rect 31724 9214 31726 9266
rect 31778 9214 31780 9266
rect 31724 9202 31780 9214
rect 31612 9156 31668 9166
rect 31612 9062 31668 9100
rect 31836 8932 31892 8942
rect 31500 8930 31892 8932
rect 31500 8878 31838 8930
rect 31890 8878 31892 8930
rect 31500 8876 31892 8878
rect 30940 8866 30996 8876
rect 31836 8866 31892 8876
rect 31164 8372 31220 8382
rect 31164 8034 31220 8316
rect 32284 8370 32340 9772
rect 32732 9602 32788 9614
rect 32732 9550 32734 9602
rect 32786 9550 32788 9602
rect 32396 9154 32452 9166
rect 32396 9102 32398 9154
rect 32450 9102 32452 9154
rect 32396 8708 32452 9102
rect 32732 9154 32788 9550
rect 32844 9604 32900 9772
rect 32844 9538 32900 9548
rect 32732 9102 32734 9154
rect 32786 9102 32788 9154
rect 32732 9090 32788 9102
rect 32396 8642 32452 8652
rect 32284 8318 32286 8370
rect 32338 8318 32340 8370
rect 32284 8306 32340 8318
rect 31164 7982 31166 8034
rect 31218 7982 31220 8034
rect 31164 7252 31220 7982
rect 31948 8258 32004 8270
rect 31948 8206 31950 8258
rect 32002 8206 32004 8258
rect 31612 7476 31668 7486
rect 31276 7364 31332 7374
rect 31276 7270 31332 7308
rect 31164 7186 31220 7196
rect 30828 6078 30830 6130
rect 30882 6078 30884 6130
rect 30380 4958 30382 5010
rect 30434 4958 30436 5010
rect 30380 4788 30436 4958
rect 30380 4722 30436 4732
rect 30828 5796 30884 6078
rect 31612 6690 31668 7420
rect 31836 7364 31892 7374
rect 31836 6914 31892 7308
rect 31836 6862 31838 6914
rect 31890 6862 31892 6914
rect 31836 6850 31892 6862
rect 31612 6638 31614 6690
rect 31666 6638 31668 6690
rect 30380 4564 30436 4574
rect 30380 4470 30436 4508
rect 30828 4564 30884 5740
rect 30940 5906 30996 5918
rect 30940 5854 30942 5906
rect 30994 5854 30996 5906
rect 30940 4900 30996 5854
rect 31612 5572 31668 6638
rect 31948 6692 32004 8206
rect 32172 8258 32228 8270
rect 32172 8206 32174 8258
rect 32226 8206 32228 8258
rect 32172 7364 32228 8206
rect 32508 8260 32564 8270
rect 32508 8258 32788 8260
rect 32508 8206 32510 8258
rect 32562 8206 32788 8258
rect 32508 8204 32788 8206
rect 32508 8194 32564 8204
rect 32620 7476 32676 7486
rect 32620 7382 32676 7420
rect 32172 7362 32340 7364
rect 32172 7310 32174 7362
rect 32226 7310 32340 7362
rect 32172 7308 32340 7310
rect 32172 7298 32228 7308
rect 32172 6692 32228 6702
rect 31948 6690 32228 6692
rect 31948 6638 32174 6690
rect 32226 6638 32228 6690
rect 31948 6636 32228 6638
rect 32172 6626 32228 6636
rect 32060 5908 32116 5918
rect 32284 5908 32340 7308
rect 32732 6804 32788 8204
rect 32844 8036 32900 8046
rect 32844 7942 32900 7980
rect 32844 6804 32900 6814
rect 32060 5906 32340 5908
rect 32060 5854 32062 5906
rect 32114 5854 32340 5906
rect 32060 5852 32340 5854
rect 32396 6802 32900 6804
rect 32396 6750 32846 6802
rect 32898 6750 32900 6802
rect 32396 6748 32900 6750
rect 32396 5906 32452 6748
rect 32844 6738 32900 6748
rect 32956 6692 33012 10780
rect 33404 9268 33460 11116
rect 33516 10612 33572 11564
rect 33628 11172 33684 11182
rect 33628 10836 33684 11116
rect 33740 11060 33796 12348
rect 33964 12402 34020 13804
rect 34300 14084 34356 14094
rect 34300 13858 34356 14028
rect 34300 13806 34302 13858
rect 34354 13806 34356 13858
rect 34300 13794 34356 13806
rect 34076 13636 34132 13646
rect 34076 13542 34132 13580
rect 34412 13076 34468 15822
rect 34524 15538 34580 17052
rect 34748 17106 34804 18284
rect 34860 17220 34916 19180
rect 34972 18226 35028 19404
rect 35084 19012 35140 20076
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35084 18956 35252 19012
rect 35196 18452 35252 18956
rect 35308 18676 35364 18686
rect 35532 18676 35588 20188
rect 35308 18674 35588 18676
rect 35308 18622 35310 18674
rect 35362 18622 35588 18674
rect 35308 18620 35588 18622
rect 35308 18610 35364 18620
rect 35644 18564 35700 21644
rect 36316 21634 36372 21644
rect 35868 21588 35924 21598
rect 35756 21532 35868 21588
rect 35756 21028 35812 21532
rect 35868 21456 35924 21532
rect 36092 21588 36148 21598
rect 36092 21586 36260 21588
rect 36092 21534 36094 21586
rect 36146 21534 36260 21586
rect 36092 21532 36260 21534
rect 36092 21522 36148 21532
rect 35756 20802 35812 20972
rect 36092 20916 36148 20926
rect 36092 20822 36148 20860
rect 35756 20750 35758 20802
rect 35810 20750 35812 20802
rect 35756 20738 35812 20750
rect 35868 20580 35924 20590
rect 35868 20130 35924 20524
rect 35868 20078 35870 20130
rect 35922 20078 35924 20130
rect 35868 20066 35924 20078
rect 35980 20578 36036 20590
rect 35980 20526 35982 20578
rect 36034 20526 36036 20578
rect 35980 20132 36036 20526
rect 35980 20066 36036 20076
rect 36092 20580 36148 20590
rect 36204 20580 36260 21532
rect 36428 21476 36484 25788
rect 36540 25618 36596 26796
rect 36652 26740 36708 26910
rect 36652 26674 36708 26684
rect 36540 25566 36542 25618
rect 36594 25566 36596 25618
rect 36540 25554 36596 25566
rect 36652 26180 36708 26190
rect 36652 24946 36708 26124
rect 36652 24894 36654 24946
rect 36706 24894 36708 24946
rect 36652 24882 36708 24894
rect 36764 24388 36820 28028
rect 36876 27524 36932 31052
rect 36988 30994 37044 31006
rect 36988 30942 36990 30994
rect 37042 30942 37044 30994
rect 36988 30100 37044 30942
rect 36988 30034 37044 30044
rect 36988 27970 37044 27982
rect 36988 27918 36990 27970
rect 37042 27918 37044 27970
rect 36988 27860 37044 27918
rect 36988 27794 37044 27804
rect 37100 27858 37156 27870
rect 37100 27806 37102 27858
rect 37154 27806 37156 27858
rect 37100 27636 37156 27806
rect 37100 27570 37156 27580
rect 36876 27458 36932 27468
rect 36876 27188 36932 27198
rect 36876 26908 36932 27132
rect 37212 26908 37268 56588
rect 37548 55522 37604 57372
rect 38108 57204 38164 57822
rect 38892 57876 38948 58158
rect 38892 57810 38948 57820
rect 39116 58156 39396 58212
rect 38108 57138 38164 57148
rect 38220 57650 38276 57662
rect 38220 57598 38222 57650
rect 38274 57598 38276 57650
rect 38220 57092 38276 57598
rect 38444 57650 38500 57662
rect 38444 57598 38446 57650
rect 38498 57598 38500 57650
rect 38220 57026 38276 57036
rect 38332 57538 38388 57550
rect 38332 57486 38334 57538
rect 38386 57486 38388 57538
rect 37772 56980 37828 56990
rect 37660 56644 37716 56654
rect 37772 56644 37828 56924
rect 38332 56868 38388 57486
rect 38444 57092 38500 57598
rect 38668 57650 38724 57662
rect 38668 57598 38670 57650
rect 38722 57598 38724 57650
rect 38668 57316 38724 57598
rect 38668 57204 38724 57260
rect 38444 57026 38500 57036
rect 38556 57148 38724 57204
rect 38780 57652 38836 57662
rect 39116 57652 39172 58156
rect 39676 57874 39732 59724
rect 42924 59778 42980 59790
rect 42924 59726 42926 59778
rect 42978 59726 42980 59778
rect 40796 59556 40852 59566
rect 40572 59332 40628 59342
rect 40572 59218 40628 59276
rect 40572 59166 40574 59218
rect 40626 59166 40628 59218
rect 40572 59154 40628 59166
rect 40012 58994 40068 59006
rect 40012 58942 40014 58994
rect 40066 58942 40068 58994
rect 40012 58434 40068 58942
rect 40348 58996 40404 59006
rect 40348 58902 40404 58940
rect 40572 58884 40628 58894
rect 40572 58658 40628 58828
rect 40572 58606 40574 58658
rect 40626 58606 40628 58658
rect 40572 58594 40628 58606
rect 40796 58548 40852 59500
rect 42924 59444 42980 59726
rect 42252 59388 43428 59444
rect 42028 59332 42084 59342
rect 41468 59220 41524 59230
rect 41468 59126 41524 59164
rect 41804 58996 41860 59006
rect 41580 58772 41636 58782
rect 40796 58482 40852 58492
rect 41244 58660 41300 58670
rect 41244 58546 41300 58604
rect 41244 58494 41246 58546
rect 41298 58494 41300 58546
rect 41244 58482 41300 58494
rect 40012 58382 40014 58434
rect 40066 58382 40068 58434
rect 40012 58370 40068 58382
rect 40348 58436 40404 58446
rect 40236 58324 40292 58334
rect 40236 58230 40292 58268
rect 39676 57822 39678 57874
rect 39730 57822 39732 57874
rect 39676 57810 39732 57822
rect 40124 58210 40180 58222
rect 40124 58158 40126 58210
rect 40178 58158 40180 58210
rect 38556 56980 38612 57148
rect 38780 57092 38836 57596
rect 38556 56914 38612 56924
rect 38668 57036 38836 57092
rect 38892 57596 39172 57652
rect 39228 57650 39284 57662
rect 39228 57598 39230 57650
rect 39282 57598 39284 57650
rect 38332 56802 38388 56812
rect 38668 56866 38724 57036
rect 38668 56814 38670 56866
rect 38722 56814 38724 56866
rect 38668 56802 38724 56814
rect 38780 56868 38836 56878
rect 38780 56774 38836 56812
rect 38556 56756 38612 56766
rect 38556 56662 38612 56700
rect 37660 56642 37828 56644
rect 37660 56590 37662 56642
rect 37714 56590 37828 56642
rect 37660 56588 37828 56590
rect 37660 56578 37716 56588
rect 37548 55470 37550 55522
rect 37602 55470 37604 55522
rect 37548 55458 37604 55470
rect 37548 53620 37604 53630
rect 37548 52946 37604 53564
rect 37548 52894 37550 52946
rect 37602 52894 37604 52946
rect 37548 52882 37604 52894
rect 37548 51604 37604 51614
rect 37548 51510 37604 51548
rect 37324 51380 37380 51390
rect 37324 51286 37380 51324
rect 37660 51154 37716 51166
rect 37660 51102 37662 51154
rect 37714 51102 37716 51154
rect 37660 51044 37716 51102
rect 37660 50978 37716 50988
rect 37660 50708 37716 50718
rect 37660 50614 37716 50652
rect 37548 49698 37604 49710
rect 37548 49646 37550 49698
rect 37602 49646 37604 49698
rect 37548 49140 37604 49646
rect 37548 49074 37604 49084
rect 37548 48802 37604 48814
rect 37548 48750 37550 48802
rect 37602 48750 37604 48802
rect 37436 47460 37492 47470
rect 37436 47366 37492 47404
rect 37548 47348 37604 48750
rect 37548 47282 37604 47292
rect 37772 47236 37828 56588
rect 38220 56420 38276 56430
rect 38220 56306 38276 56364
rect 38220 56254 38222 56306
rect 38274 56254 38276 56306
rect 38220 56242 38276 56254
rect 38556 55972 38612 55982
rect 38668 55972 38724 55982
rect 38556 55970 38668 55972
rect 38556 55918 38558 55970
rect 38610 55918 38668 55970
rect 38556 55916 38668 55918
rect 38556 55524 38612 55916
rect 38668 55906 38724 55916
rect 38556 55458 38612 55468
rect 38780 55524 38836 55534
rect 38892 55524 38948 57596
rect 39116 56756 39172 56766
rect 39004 56642 39060 56654
rect 39004 56590 39006 56642
rect 39058 56590 39060 56642
rect 39004 56532 39060 56590
rect 39004 56466 39060 56476
rect 39116 56082 39172 56700
rect 39116 56030 39118 56082
rect 39170 56030 39172 56082
rect 39116 56018 39172 56030
rect 39228 55972 39284 57598
rect 39452 57652 39508 57662
rect 39452 57558 39508 57596
rect 39788 57650 39844 57662
rect 39788 57598 39790 57650
rect 39842 57598 39844 57650
rect 39340 56868 39396 56878
rect 39340 56774 39396 56812
rect 39452 56866 39508 56878
rect 39452 56814 39454 56866
rect 39506 56814 39508 56866
rect 39452 56196 39508 56814
rect 39788 56420 39844 57598
rect 40012 56868 40068 56878
rect 40124 56868 40180 58158
rect 40348 57762 40404 58380
rect 40572 58434 40628 58446
rect 40572 58382 40574 58434
rect 40626 58382 40628 58434
rect 40460 57876 40516 57886
rect 40572 57876 40628 58382
rect 40460 57874 40628 57876
rect 40460 57822 40462 57874
rect 40514 57822 40628 57874
rect 40460 57820 40628 57822
rect 40460 57810 40516 57820
rect 40348 57710 40350 57762
rect 40402 57710 40404 57762
rect 40348 57698 40404 57710
rect 40684 57540 40740 57550
rect 41580 57540 41636 58716
rect 41804 57650 41860 58940
rect 42028 58434 42084 59276
rect 42252 59330 42308 59388
rect 42252 59278 42254 59330
rect 42306 59278 42308 59330
rect 42252 59266 42308 59278
rect 42028 58382 42030 58434
rect 42082 58382 42084 58434
rect 42028 57876 42084 58382
rect 42364 59220 42420 59230
rect 42364 58434 42420 59164
rect 42700 59220 42756 59230
rect 43036 59220 43092 59230
rect 42700 59218 43092 59220
rect 42700 59166 42702 59218
rect 42754 59166 43038 59218
rect 43090 59166 43092 59218
rect 42700 59164 43092 59166
rect 43372 59220 43428 59388
rect 43484 59220 43540 59230
rect 43372 59218 43652 59220
rect 43372 59166 43486 59218
rect 43538 59166 43652 59218
rect 43372 59164 43652 59166
rect 42700 59154 42756 59164
rect 42476 59106 42532 59118
rect 42476 59054 42478 59106
rect 42530 59054 42532 59106
rect 42476 58884 42532 59054
rect 42476 58818 42532 58828
rect 42812 58548 42868 58558
rect 42812 58454 42868 58492
rect 42364 58382 42366 58434
rect 42418 58382 42420 58434
rect 42364 58370 42420 58382
rect 43036 58212 43092 59164
rect 43484 59154 43540 59164
rect 43260 59108 43316 59118
rect 43260 59106 43428 59108
rect 43260 59054 43262 59106
rect 43314 59054 43428 59106
rect 43260 59052 43428 59054
rect 43260 59042 43316 59052
rect 43148 58548 43204 58558
rect 43148 58322 43204 58492
rect 43148 58270 43150 58322
rect 43202 58270 43204 58322
rect 43148 58258 43204 58270
rect 43036 58146 43092 58156
rect 42140 57876 42196 57886
rect 42028 57874 42196 57876
rect 42028 57822 42142 57874
rect 42194 57822 42196 57874
rect 42028 57820 42196 57822
rect 42140 57810 42196 57820
rect 43260 57876 43316 57886
rect 43372 57876 43428 59052
rect 43596 58548 43652 59164
rect 43708 59218 43764 59838
rect 43820 59780 43876 59790
rect 44940 59780 44996 59790
rect 49868 59780 49924 59790
rect 43820 59778 44212 59780
rect 43820 59726 43822 59778
rect 43874 59726 44212 59778
rect 43820 59724 44212 59726
rect 43820 59714 43876 59724
rect 43708 59166 43710 59218
rect 43762 59166 43764 59218
rect 43708 58772 43764 59166
rect 43708 58706 43764 58716
rect 43596 58482 43652 58492
rect 43484 58434 43540 58446
rect 43484 58382 43486 58434
rect 43538 58382 43540 58434
rect 43484 58212 43540 58382
rect 43484 58146 43540 58156
rect 44156 58434 44212 59724
rect 44940 59778 45108 59780
rect 44940 59726 44942 59778
rect 44994 59726 45108 59778
rect 44940 59724 45108 59726
rect 44940 59714 44996 59724
rect 44268 59218 44324 59230
rect 44268 59166 44270 59218
rect 44322 59166 44324 59218
rect 44268 58660 44324 59166
rect 44492 59220 44548 59230
rect 44940 59220 44996 59230
rect 44492 59218 44660 59220
rect 44492 59166 44494 59218
rect 44546 59166 44660 59218
rect 44492 59164 44660 59166
rect 44492 59154 44548 59164
rect 44380 59106 44436 59118
rect 44380 59054 44382 59106
rect 44434 59054 44436 59106
rect 44380 58884 44436 59054
rect 44380 58828 44548 58884
rect 44380 58660 44436 58670
rect 44268 58658 44436 58660
rect 44268 58606 44382 58658
rect 44434 58606 44436 58658
rect 44268 58604 44436 58606
rect 44156 58382 44158 58434
rect 44210 58382 44212 58434
rect 43316 57820 43428 57876
rect 43484 57876 43540 57886
rect 41804 57598 41806 57650
rect 41858 57598 41860 57650
rect 41804 57586 41860 57598
rect 42812 57650 42868 57662
rect 42812 57598 42814 57650
rect 42866 57598 42868 57650
rect 40012 56866 40180 56868
rect 40012 56814 40014 56866
rect 40066 56814 40180 56866
rect 40012 56812 40180 56814
rect 40348 56868 40404 56878
rect 40012 56802 40068 56812
rect 39788 56354 39844 56364
rect 40124 56642 40180 56654
rect 40124 56590 40126 56642
rect 40178 56590 40180 56642
rect 40012 56306 40068 56318
rect 40012 56254 40014 56306
rect 40066 56254 40068 56306
rect 40012 56196 40068 56254
rect 39452 56140 40068 56196
rect 39340 56084 39396 56094
rect 40124 56084 40180 56590
rect 40236 56644 40292 56654
rect 40236 56550 40292 56588
rect 39340 56082 40180 56084
rect 39340 56030 39342 56082
rect 39394 56030 40180 56082
rect 39340 56028 40180 56030
rect 39340 56018 39396 56028
rect 39228 55906 39284 55916
rect 40348 55970 40404 56812
rect 40684 56866 40740 57484
rect 40684 56814 40686 56866
rect 40738 56814 40740 56866
rect 40684 56802 40740 56814
rect 41468 57538 41636 57540
rect 41468 57486 41582 57538
rect 41634 57486 41636 57538
rect 41468 57484 41636 57486
rect 41020 56644 41076 56654
rect 41020 56550 41076 56588
rect 40348 55918 40350 55970
rect 40402 55918 40404 55970
rect 39564 55860 39620 55870
rect 39564 55766 39620 55804
rect 40348 55748 40404 55918
rect 40348 55682 40404 55692
rect 38780 55522 38948 55524
rect 38780 55470 38782 55522
rect 38834 55470 38948 55522
rect 38780 55468 38948 55470
rect 38780 55458 38836 55468
rect 41356 55412 41412 55422
rect 41468 55412 41524 57484
rect 41580 57474 41636 57484
rect 42588 57316 42644 57326
rect 42812 57316 42868 57598
rect 42644 57260 42868 57316
rect 42588 56978 42644 57260
rect 42588 56926 42590 56978
rect 42642 56926 42644 56978
rect 42588 56914 42644 56926
rect 42812 56308 42868 57260
rect 43260 56978 43316 57820
rect 43372 57540 43428 57550
rect 43372 57446 43428 57484
rect 43484 57090 43540 57820
rect 44156 57874 44212 58382
rect 44156 57822 44158 57874
rect 44210 57822 44212 57874
rect 44156 57810 44212 57822
rect 44268 58210 44324 58222
rect 44268 58158 44270 58210
rect 44322 58158 44324 58210
rect 44268 57876 44324 58158
rect 44380 57988 44436 58604
rect 44492 58660 44548 58828
rect 44492 58594 44548 58604
rect 44604 58436 44660 59164
rect 44940 59126 44996 59164
rect 45052 58548 45108 59724
rect 49868 59686 49924 59724
rect 50428 59780 50484 59950
rect 50428 59714 50484 59724
rect 50556 59612 50820 59622
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50556 59546 50820 59556
rect 45500 59332 45556 59342
rect 45500 59238 45556 59276
rect 45388 59220 45444 59230
rect 45388 59126 45444 59164
rect 44604 58434 44772 58436
rect 44604 58382 44606 58434
rect 44658 58382 44772 58434
rect 44604 58380 44772 58382
rect 44604 58370 44660 58380
rect 44380 57922 44436 57932
rect 44492 58324 44548 58334
rect 44268 57810 44324 57820
rect 44492 57874 44548 58268
rect 44492 57822 44494 57874
rect 44546 57822 44548 57874
rect 44492 57810 44548 57822
rect 44604 57988 44660 57998
rect 44604 57874 44660 57932
rect 44604 57822 44606 57874
rect 44658 57822 44660 57874
rect 44604 57810 44660 57822
rect 44380 57650 44436 57662
rect 44380 57598 44382 57650
rect 44434 57598 44436 57650
rect 44380 57540 44436 57598
rect 44716 57540 44772 58380
rect 45052 58212 45108 58492
rect 45948 59106 46004 59118
rect 45948 59054 45950 59106
rect 46002 59054 46004 59106
rect 45388 58212 45444 58222
rect 45052 58210 45444 58212
rect 45052 58158 45390 58210
rect 45442 58158 45444 58210
rect 45052 58156 45444 58158
rect 45388 57876 45444 58156
rect 45388 57810 45444 57820
rect 45052 57540 45108 57550
rect 45500 57540 45556 57550
rect 44380 57538 45556 57540
rect 44380 57486 45054 57538
rect 45106 57486 45502 57538
rect 45554 57486 45556 57538
rect 44380 57484 45556 57486
rect 45052 57474 45108 57484
rect 43484 57038 43486 57090
rect 43538 57038 43540 57090
rect 43484 57026 43540 57038
rect 43820 57092 43876 57102
rect 43820 56998 43876 57036
rect 44156 57092 44212 57102
rect 43260 56926 43262 56978
rect 43314 56926 43316 56978
rect 43260 56914 43316 56926
rect 42812 56176 42868 56252
rect 43932 56308 43988 56318
rect 43932 56214 43988 56252
rect 44156 56306 44212 57036
rect 45500 57092 45556 57484
rect 45500 57026 45556 57036
rect 45948 57092 46004 59054
rect 46396 58548 46452 58558
rect 46396 58454 46452 58492
rect 46732 58548 46788 58558
rect 46620 58436 46676 58446
rect 46620 58342 46676 58380
rect 46060 58210 46116 58222
rect 46060 58158 46062 58210
rect 46114 58158 46116 58210
rect 46060 57988 46116 58158
rect 46060 57922 46116 57932
rect 46732 57874 46788 58492
rect 47180 58548 47236 58558
rect 47180 58454 47236 58492
rect 50652 58548 50708 58558
rect 51212 58548 51268 58558
rect 50652 58546 51268 58548
rect 50652 58494 50654 58546
rect 50706 58494 51214 58546
rect 51266 58494 51268 58546
rect 50652 58492 51268 58494
rect 50652 58482 50708 58492
rect 47516 58436 47572 58446
rect 47516 58342 47572 58380
rect 50092 58436 50148 58446
rect 50092 58342 50148 58380
rect 50428 58434 50484 58446
rect 50428 58382 50430 58434
rect 50482 58382 50484 58434
rect 47292 58212 47348 58222
rect 47292 58118 47348 58156
rect 46732 57822 46734 57874
rect 46786 57822 46788 57874
rect 46732 57810 46788 57822
rect 50428 57764 50484 58382
rect 50556 58044 50820 58054
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50556 57978 50820 57988
rect 50204 57708 50484 57764
rect 51212 57762 51268 58492
rect 51548 58322 51604 58334
rect 51548 58270 51550 58322
rect 51602 58270 51604 58322
rect 51324 58212 51380 58222
rect 51324 58210 51492 58212
rect 51324 58158 51326 58210
rect 51378 58158 51492 58210
rect 51324 58156 51492 58158
rect 51324 58146 51380 58156
rect 51212 57710 51214 57762
rect 51266 57710 51268 57762
rect 45948 57026 46004 57036
rect 46284 57650 46340 57662
rect 46508 57652 46564 57662
rect 46284 57598 46286 57650
rect 46338 57598 46340 57650
rect 44156 56254 44158 56306
rect 44210 56254 44212 56306
rect 44156 56242 44212 56254
rect 46284 56978 46340 57598
rect 46284 56926 46286 56978
rect 46338 56926 46340 56978
rect 44604 56084 44660 56094
rect 44604 55990 44660 56028
rect 43372 55972 43428 55982
rect 43260 55524 43316 55534
rect 43260 55430 43316 55468
rect 41356 55410 41524 55412
rect 41356 55358 41358 55410
rect 41410 55358 41524 55410
rect 41356 55356 41524 55358
rect 42588 55410 42644 55422
rect 42588 55358 42590 55410
rect 42642 55358 42644 55410
rect 41356 55346 41412 55356
rect 37884 55298 37940 55310
rect 37884 55246 37886 55298
rect 37938 55246 37940 55298
rect 37884 55188 37940 55246
rect 38108 55300 38164 55310
rect 39452 55300 39508 55310
rect 38108 55206 38164 55244
rect 39340 55244 39452 55300
rect 37884 55122 37940 55132
rect 38668 55188 38724 55198
rect 38668 55094 38724 55132
rect 38780 55074 38836 55086
rect 38780 55022 38782 55074
rect 38834 55022 38836 55074
rect 38780 54740 38836 55022
rect 38780 54674 38836 54684
rect 39340 54402 39396 55244
rect 39452 55206 39508 55244
rect 39676 55300 39732 55310
rect 39676 55206 39732 55244
rect 40460 55300 40516 55310
rect 40460 55206 40516 55244
rect 40684 55298 40740 55310
rect 40684 55246 40686 55298
rect 40738 55246 40740 55298
rect 39788 55186 39844 55198
rect 39788 55134 39790 55186
rect 39842 55134 39844 55186
rect 39788 54740 39844 55134
rect 40684 55188 40740 55246
rect 40684 55122 40740 55132
rect 41580 55300 41636 55310
rect 39788 54674 39844 54684
rect 40460 55076 40516 55086
rect 39452 54628 39508 54638
rect 39452 54626 39620 54628
rect 39452 54574 39454 54626
rect 39506 54574 39620 54626
rect 39452 54572 39620 54574
rect 39452 54562 39508 54572
rect 39340 54350 39342 54402
rect 39394 54350 39396 54402
rect 39340 54338 39396 54350
rect 38332 53732 38388 53742
rect 38332 53058 38388 53676
rect 39564 53732 39620 54572
rect 39564 53638 39620 53676
rect 39676 54290 39732 54302
rect 39676 54238 39678 54290
rect 39730 54238 39732 54290
rect 39676 53842 39732 54238
rect 40348 53956 40404 53966
rect 40348 53862 40404 53900
rect 39676 53790 39678 53842
rect 39730 53790 39732 53842
rect 39564 53172 39620 53182
rect 39676 53172 39732 53790
rect 39564 53170 39732 53172
rect 39564 53118 39566 53170
rect 39618 53118 39732 53170
rect 39564 53116 39732 53118
rect 39564 53106 39620 53116
rect 38332 53006 38334 53058
rect 38386 53006 38388 53058
rect 38332 52994 38388 53006
rect 39340 52946 39396 52958
rect 39340 52894 39342 52946
rect 39394 52894 39396 52946
rect 39340 52276 39396 52894
rect 39228 52164 39284 52174
rect 39004 51380 39060 51390
rect 39004 51378 39172 51380
rect 39004 51326 39006 51378
rect 39058 51326 39172 51378
rect 39004 51324 39172 51326
rect 39004 51314 39060 51324
rect 38556 50708 38612 50718
rect 38556 50614 38612 50652
rect 37884 50596 37940 50606
rect 37884 50502 37940 50540
rect 39116 50594 39172 51324
rect 39116 50542 39118 50594
rect 39170 50542 39172 50594
rect 38556 50484 38612 50494
rect 38332 49140 38388 49150
rect 38332 49046 38388 49084
rect 37884 48802 37940 48814
rect 37884 48750 37886 48802
rect 37938 48750 37940 48802
rect 37884 48692 37940 48750
rect 37884 48626 37940 48636
rect 37884 48244 37940 48254
rect 37884 48150 37940 48188
rect 38108 48242 38164 48254
rect 38108 48190 38110 48242
rect 38162 48190 38164 48242
rect 37772 47170 37828 47180
rect 37996 47234 38052 47246
rect 37996 47182 37998 47234
rect 38050 47182 38052 47234
rect 37996 47124 38052 47182
rect 37996 47058 38052 47068
rect 38108 47236 38164 48190
rect 38444 48244 38500 48254
rect 38444 47458 38500 48188
rect 38556 47570 38612 50428
rect 39116 50484 39172 50542
rect 39116 50418 39172 50428
rect 39228 50260 39284 52108
rect 39340 51604 39396 52220
rect 39564 52946 39620 52958
rect 39564 52894 39566 52946
rect 39618 52894 39620 52946
rect 39564 52836 39620 52894
rect 39564 52164 39620 52780
rect 39788 52946 39844 52958
rect 39788 52894 39790 52946
rect 39842 52894 39844 52946
rect 39788 52388 39844 52894
rect 40348 52836 40404 52846
rect 40348 52742 40404 52780
rect 39564 52098 39620 52108
rect 39676 52332 39844 52388
rect 39340 51548 39508 51604
rect 39452 51490 39508 51548
rect 39452 51438 39454 51490
rect 39506 51438 39508 51490
rect 39452 51426 39508 51438
rect 39340 51378 39396 51390
rect 39340 51326 39342 51378
rect 39394 51326 39396 51378
rect 39340 50818 39396 51326
rect 39340 50766 39342 50818
rect 39394 50766 39396 50818
rect 39340 50708 39396 50766
rect 39676 50818 39732 52332
rect 39900 52276 39956 52286
rect 39900 52182 39956 52220
rect 39788 52164 39844 52174
rect 39788 52070 39844 52108
rect 39900 51266 39956 51278
rect 39900 51214 39902 51266
rect 39954 51214 39956 51266
rect 39676 50766 39678 50818
rect 39730 50766 39732 50818
rect 39676 50754 39732 50766
rect 39788 51044 39844 51054
rect 39340 50642 39396 50652
rect 39004 50204 39284 50260
rect 38780 48132 38836 48142
rect 38780 48038 38836 48076
rect 38556 47518 38558 47570
rect 38610 47518 38612 47570
rect 38556 47506 38612 47518
rect 38444 47406 38446 47458
rect 38498 47406 38500 47458
rect 38444 47394 38500 47406
rect 38108 46898 38164 47180
rect 38668 47236 38724 47246
rect 38668 47142 38724 47180
rect 38108 46846 38110 46898
rect 38162 46846 38164 46898
rect 38108 46834 38164 46846
rect 38444 46900 38500 46910
rect 38444 46806 38500 46844
rect 37884 46786 37940 46798
rect 37884 46734 37886 46786
rect 37938 46734 37940 46786
rect 37772 46674 37828 46686
rect 37772 46622 37774 46674
rect 37826 46622 37828 46674
rect 37772 46116 37828 46622
rect 37772 46050 37828 46060
rect 37772 45892 37828 45902
rect 37884 45892 37940 46734
rect 38556 46116 38612 46126
rect 38556 46022 38612 46060
rect 37996 46004 38052 46014
rect 37996 45910 38052 45948
rect 37828 45836 37940 45892
rect 37772 45798 37828 45836
rect 38668 45780 38724 45790
rect 38444 45668 38500 45678
rect 38444 45330 38500 45612
rect 38444 45278 38446 45330
rect 38498 45278 38500 45330
rect 38444 45266 38500 45278
rect 38220 45220 38276 45230
rect 38108 45106 38164 45118
rect 38108 45054 38110 45106
rect 38162 45054 38164 45106
rect 37548 44996 37604 45006
rect 37548 43764 37604 44940
rect 37548 43698 37604 43708
rect 37884 44436 37940 44446
rect 38108 44436 38164 45054
rect 37884 44434 38164 44436
rect 37884 44382 37886 44434
rect 37938 44382 38164 44434
rect 37884 44380 38164 44382
rect 37884 43652 37940 44380
rect 38220 44322 38276 45164
rect 38220 44270 38222 44322
rect 38274 44270 38276 44322
rect 38220 44258 38276 44270
rect 37884 43586 37940 43596
rect 38108 44212 38164 44222
rect 37324 43540 37380 43550
rect 37324 43446 37380 43484
rect 37884 43428 37940 43438
rect 37548 43426 37940 43428
rect 37548 43374 37886 43426
rect 37938 43374 37940 43426
rect 37548 43372 37940 43374
rect 37548 42420 37604 43372
rect 37884 43362 37940 43372
rect 38108 42754 38164 44156
rect 38220 43764 38276 43774
rect 38276 43708 38388 43764
rect 38220 43670 38276 43708
rect 38108 42702 38110 42754
rect 38162 42702 38164 42754
rect 38108 42690 38164 42702
rect 37436 42196 37492 42206
rect 37436 42102 37492 42140
rect 37548 42194 37604 42364
rect 37772 42642 37828 42654
rect 37772 42590 37774 42642
rect 37826 42590 37828 42642
rect 37548 42142 37550 42194
rect 37602 42142 37604 42194
rect 37548 42130 37604 42142
rect 37660 42308 37716 42318
rect 37660 42194 37716 42252
rect 37660 42142 37662 42194
rect 37714 42142 37716 42194
rect 37660 42130 37716 42142
rect 37324 42082 37380 42094
rect 37324 42030 37326 42082
rect 37378 42030 37380 42082
rect 37324 41972 37380 42030
rect 37324 41906 37380 41916
rect 37772 41412 37828 42590
rect 37996 42644 38052 42654
rect 37660 41356 37828 41412
rect 37884 42530 37940 42542
rect 37884 42478 37886 42530
rect 37938 42478 37940 42530
rect 37884 42084 37940 42478
rect 37660 41186 37716 41356
rect 37660 41134 37662 41186
rect 37714 41134 37716 41186
rect 37324 40402 37380 40414
rect 37324 40350 37326 40402
rect 37378 40350 37380 40402
rect 37324 40292 37380 40350
rect 37660 40404 37716 41134
rect 37660 40338 37716 40348
rect 37772 41188 37828 41198
rect 37772 40626 37828 41132
rect 37884 41186 37940 42028
rect 37884 41134 37886 41186
rect 37938 41134 37940 41186
rect 37884 41122 37940 41134
rect 37996 41636 38052 42588
rect 38332 42082 38388 43708
rect 38668 43708 38724 45724
rect 38780 45332 38836 45342
rect 38780 45238 38836 45276
rect 38780 44436 38836 44446
rect 38780 44322 38836 44380
rect 38780 44270 38782 44322
rect 38834 44270 38836 44322
rect 38780 44258 38836 44270
rect 39004 43708 39060 50204
rect 39788 50034 39844 50988
rect 39900 50820 39956 51214
rect 39900 50754 39956 50764
rect 40348 50820 40404 50830
rect 40236 50706 40292 50718
rect 40236 50654 40238 50706
rect 40290 50654 40292 50706
rect 40236 50428 40292 50654
rect 39788 49982 39790 50034
rect 39842 49982 39844 50034
rect 39788 49970 39844 49982
rect 39900 50372 40292 50428
rect 40348 50484 40404 50764
rect 40348 50418 40404 50428
rect 40460 50428 40516 55020
rect 41580 54514 41636 55244
rect 42476 55300 42532 55310
rect 42476 55206 42532 55244
rect 41804 54740 41860 54750
rect 41804 54646 41860 54684
rect 41916 54628 41972 54638
rect 41916 54534 41972 54572
rect 42588 54628 42644 55358
rect 43372 55076 43428 55916
rect 44044 55970 44100 55982
rect 44044 55918 44046 55970
rect 44098 55918 44100 55970
rect 44044 55860 44100 55918
rect 44380 55972 44436 55982
rect 44380 55878 44436 55916
rect 44828 55972 44884 55982
rect 44828 55878 44884 55916
rect 44044 55794 44100 55804
rect 46284 55524 46340 56926
rect 46284 55458 46340 55468
rect 46396 57650 46564 57652
rect 46396 57598 46510 57650
rect 46562 57598 46564 57650
rect 46396 57596 46564 57598
rect 46396 56866 46452 57596
rect 46508 57586 46564 57596
rect 46956 57652 47012 57662
rect 46956 57558 47012 57596
rect 47516 57650 47572 57662
rect 47516 57598 47518 57650
rect 47570 57598 47572 57650
rect 47068 57428 47124 57438
rect 47068 57090 47124 57372
rect 47516 57428 47572 57598
rect 47740 57652 47796 57662
rect 47740 57558 47796 57596
rect 48076 57652 48132 57662
rect 48412 57652 48468 57662
rect 48076 57650 48244 57652
rect 48076 57598 48078 57650
rect 48130 57598 48244 57650
rect 48076 57596 48244 57598
rect 48076 57586 48132 57596
rect 47516 57362 47572 57372
rect 47852 57538 47908 57550
rect 47852 57486 47854 57538
rect 47906 57486 47908 57538
rect 47068 57038 47070 57090
rect 47122 57038 47124 57090
rect 47068 57026 47124 57038
rect 46396 56814 46398 56866
rect 46450 56814 46452 56866
rect 43372 55010 43428 55020
rect 46396 54738 46452 56814
rect 46508 56644 46564 56654
rect 46508 56194 46564 56588
rect 47740 56644 47796 56654
rect 47740 56550 47796 56588
rect 46508 56142 46510 56194
rect 46562 56142 46564 56194
rect 46508 56084 46564 56142
rect 46508 56018 46564 56028
rect 46732 56084 46788 56094
rect 46732 55990 46788 56028
rect 47852 56084 47908 57486
rect 48188 56868 48244 57596
rect 48188 56774 48244 56812
rect 48300 57428 48356 57438
rect 48300 56866 48356 57372
rect 48300 56814 48302 56866
rect 48354 56814 48356 56866
rect 48300 56802 48356 56814
rect 48412 56754 48468 57596
rect 50204 57650 50260 57708
rect 51212 57698 51268 57710
rect 50204 57598 50206 57650
rect 50258 57598 50260 57650
rect 49980 57540 50036 57550
rect 49980 56866 50036 57484
rect 49980 56814 49982 56866
rect 50034 56814 50036 56866
rect 49980 56802 50036 56814
rect 50092 56868 50148 56878
rect 50092 56774 50148 56812
rect 48412 56702 48414 56754
rect 48466 56702 48468 56754
rect 48412 56420 48468 56702
rect 47852 56018 47908 56028
rect 48188 56364 48468 56420
rect 50204 56642 50260 57598
rect 50204 56590 50206 56642
rect 50258 56590 50260 56642
rect 46508 55860 46564 55870
rect 46508 55412 46564 55804
rect 47068 55860 47124 55870
rect 47068 55858 47348 55860
rect 47068 55806 47070 55858
rect 47122 55806 47348 55858
rect 47068 55804 47348 55806
rect 47068 55794 47124 55804
rect 46508 55410 47012 55412
rect 46508 55358 46510 55410
rect 46562 55358 47012 55410
rect 46508 55356 47012 55358
rect 46508 55346 46564 55356
rect 46956 55298 47012 55356
rect 46956 55246 46958 55298
rect 47010 55246 47012 55298
rect 46956 55234 47012 55246
rect 47292 55298 47348 55804
rect 47852 55748 47908 55758
rect 47852 55410 47908 55692
rect 47852 55358 47854 55410
rect 47906 55358 47908 55410
rect 47852 55346 47908 55358
rect 47516 55300 47572 55310
rect 47292 55246 47294 55298
rect 47346 55246 47348 55298
rect 47292 55234 47348 55246
rect 47404 55298 47572 55300
rect 47404 55246 47518 55298
rect 47570 55246 47572 55298
rect 47404 55244 47572 55246
rect 46396 54686 46398 54738
rect 46450 54686 46452 54738
rect 46396 54674 46452 54686
rect 47404 54738 47460 55244
rect 47516 55234 47572 55244
rect 47740 55300 47796 55310
rect 47740 55206 47796 55244
rect 47404 54686 47406 54738
rect 47458 54686 47460 54738
rect 47404 54674 47460 54686
rect 47964 55186 48020 55198
rect 47964 55134 47966 55186
rect 48018 55134 48020 55186
rect 47964 54740 48020 55134
rect 47964 54674 48020 54684
rect 48076 55188 48132 55198
rect 42644 54572 42868 54628
rect 42588 54562 42644 54572
rect 41580 54462 41582 54514
rect 41634 54462 41636 54514
rect 41580 53956 41636 54462
rect 41580 53890 41636 53900
rect 41692 54292 41748 54302
rect 40572 53844 40628 53854
rect 40572 52386 40628 53788
rect 41692 53844 41748 54236
rect 41692 53730 41748 53788
rect 41692 53678 41694 53730
rect 41746 53678 41748 53730
rect 41692 53666 41748 53678
rect 42700 53842 42756 53854
rect 42700 53790 42702 53842
rect 42754 53790 42756 53842
rect 41804 53506 41860 53518
rect 41804 53454 41806 53506
rect 41858 53454 41860 53506
rect 41804 53284 41860 53454
rect 42028 53508 42084 53518
rect 42028 53506 42644 53508
rect 42028 53454 42030 53506
rect 42082 53454 42644 53506
rect 42028 53452 42644 53454
rect 42028 53442 42084 53452
rect 42140 53284 42196 53294
rect 41804 53228 42140 53284
rect 40572 52334 40574 52386
rect 40626 52334 40628 52386
rect 40572 52322 40628 52334
rect 41132 52164 41188 52174
rect 41132 52070 41188 52108
rect 42140 51602 42196 53228
rect 42588 52946 42644 53452
rect 42700 53284 42756 53790
rect 42700 53218 42756 53228
rect 42812 53170 42868 54572
rect 42924 54626 42980 54638
rect 42924 54574 42926 54626
rect 42978 54574 42980 54626
rect 42924 53284 42980 54574
rect 46172 54628 46228 54638
rect 46172 54626 46340 54628
rect 46172 54574 46174 54626
rect 46226 54574 46340 54626
rect 46172 54572 46340 54574
rect 46172 54562 46228 54572
rect 46060 54516 46116 54526
rect 45948 54514 46116 54516
rect 45948 54462 46062 54514
rect 46114 54462 46116 54514
rect 45948 54460 46116 54462
rect 43036 54402 43092 54414
rect 43036 54350 43038 54402
rect 43090 54350 43092 54402
rect 43036 53956 43092 54350
rect 43148 54292 43204 54302
rect 43148 54198 43204 54236
rect 44044 54292 44100 54302
rect 43036 53900 43316 53956
rect 42924 53218 42980 53228
rect 43036 53618 43092 53630
rect 43036 53566 43038 53618
rect 43090 53566 43092 53618
rect 42812 53118 42814 53170
rect 42866 53118 42868 53170
rect 42812 53106 42868 53118
rect 42588 52894 42590 52946
rect 42642 52894 42644 52946
rect 42588 52882 42644 52894
rect 43036 52946 43092 53566
rect 43260 53058 43316 53900
rect 44044 53730 44100 54236
rect 44716 53844 44772 53854
rect 44716 53750 44772 53788
rect 45948 53844 46004 54460
rect 46060 54450 46116 54460
rect 45948 53750 46004 53788
rect 46172 53732 46228 53742
rect 46284 53732 46340 54572
rect 47292 54626 47348 54638
rect 47292 54574 47294 54626
rect 47346 54574 47348 54626
rect 47292 54516 47348 54574
rect 48076 54516 48132 55132
rect 47292 54514 48132 54516
rect 47292 54462 48078 54514
rect 48130 54462 48132 54514
rect 47292 54460 48132 54462
rect 44044 53678 44046 53730
rect 44098 53678 44100 53730
rect 44044 53666 44100 53678
rect 46060 53730 46340 53732
rect 46060 53678 46174 53730
rect 46226 53678 46340 53730
rect 46060 53676 46340 53678
rect 46844 53732 46900 53742
rect 43260 53006 43262 53058
rect 43314 53006 43316 53058
rect 43260 52994 43316 53006
rect 45276 53396 45332 53406
rect 43036 52894 43038 52946
rect 43090 52894 43092 52946
rect 42140 51550 42142 51602
rect 42194 51550 42196 51602
rect 42140 51538 42196 51550
rect 42252 51490 42308 51502
rect 42252 51438 42254 51490
rect 42306 51438 42308 51490
rect 42028 51156 42084 51166
rect 41804 51154 42084 51156
rect 41804 51102 42030 51154
rect 42082 51102 42084 51154
rect 41804 51100 42084 51102
rect 41804 50706 41860 51100
rect 42028 51090 42084 51100
rect 41916 50820 41972 50830
rect 41916 50726 41972 50764
rect 41804 50654 41806 50706
rect 41858 50654 41860 50706
rect 41804 50642 41860 50654
rect 40572 50596 40628 50606
rect 41020 50596 41076 50606
rect 40572 50594 41076 50596
rect 40572 50542 40574 50594
rect 40626 50542 41022 50594
rect 41074 50542 41076 50594
rect 40572 50540 41076 50542
rect 40572 50530 40628 50540
rect 40908 50428 40964 50438
rect 40460 50372 40740 50428
rect 39676 49924 39732 49934
rect 39676 49830 39732 49868
rect 39900 49922 39956 50372
rect 39900 49870 39902 49922
rect 39954 49870 39956 49922
rect 39900 49858 39956 49870
rect 40348 49924 40404 49934
rect 40348 49830 40404 49868
rect 39564 48916 39620 48926
rect 40460 48916 40516 48926
rect 39564 48914 39732 48916
rect 39564 48862 39566 48914
rect 39618 48862 39732 48914
rect 39564 48860 39732 48862
rect 39564 48850 39620 48860
rect 39228 48802 39284 48814
rect 39228 48750 39230 48802
rect 39282 48750 39284 48802
rect 39116 47460 39172 47470
rect 39228 47460 39284 48750
rect 39452 48802 39508 48814
rect 39452 48750 39454 48802
rect 39506 48750 39508 48802
rect 39452 48244 39508 48750
rect 39564 48244 39620 48254
rect 39452 48242 39620 48244
rect 39452 48190 39566 48242
rect 39618 48190 39620 48242
rect 39452 48188 39620 48190
rect 39116 47458 39284 47460
rect 39116 47406 39118 47458
rect 39170 47406 39284 47458
rect 39116 47404 39284 47406
rect 39116 47394 39172 47404
rect 39452 47348 39508 47358
rect 39452 47254 39508 47292
rect 39564 46900 39620 48188
rect 39676 48132 39732 48860
rect 40460 48354 40516 48860
rect 40460 48302 40462 48354
rect 40514 48302 40516 48354
rect 40460 48290 40516 48302
rect 40684 48356 40740 50372
rect 41020 50428 41076 50540
rect 41580 50596 41636 50606
rect 41580 50502 41636 50540
rect 41020 50372 41188 50428
rect 40684 48290 40740 48300
rect 40796 48804 40852 48814
rect 39676 48038 39732 48076
rect 40796 47570 40852 48748
rect 40796 47518 40798 47570
rect 40850 47518 40852 47570
rect 40796 47506 40852 47518
rect 40012 47460 40068 47470
rect 39116 46844 39620 46900
rect 39676 47348 39732 47358
rect 39116 45780 39172 46844
rect 39564 46674 39620 46686
rect 39564 46622 39566 46674
rect 39618 46622 39620 46674
rect 39228 46562 39284 46574
rect 39228 46510 39230 46562
rect 39282 46510 39284 46562
rect 39228 46116 39284 46510
rect 39340 46116 39396 46126
rect 39284 46114 39396 46116
rect 39284 46062 39342 46114
rect 39394 46062 39396 46114
rect 39284 46060 39396 46062
rect 39228 45984 39284 46060
rect 39340 46050 39396 46060
rect 39452 46004 39508 46014
rect 39116 45724 39396 45780
rect 38668 43652 38948 43708
rect 39004 43652 39284 43708
rect 38668 43428 38724 43438
rect 38444 43426 38724 43428
rect 38444 43374 38670 43426
rect 38722 43374 38724 43426
rect 38444 43372 38724 43374
rect 38444 42532 38500 43372
rect 38668 43362 38724 43372
rect 38444 42194 38500 42476
rect 38444 42142 38446 42194
rect 38498 42142 38500 42194
rect 38444 42130 38500 42142
rect 38780 43314 38836 43326
rect 38780 43262 38782 43314
rect 38834 43262 38836 43314
rect 38332 42030 38334 42082
rect 38386 42030 38388 42082
rect 38332 42018 38388 42030
rect 38668 41972 38724 41982
rect 38668 41878 38724 41916
rect 37772 40574 37774 40626
rect 37826 40574 37828 40626
rect 37324 38948 37380 40236
rect 37548 39172 37604 39182
rect 37548 39058 37604 39116
rect 37548 39006 37550 39058
rect 37602 39006 37604 39058
rect 37548 38994 37604 39006
rect 37324 38668 37380 38892
rect 37324 38612 37716 38668
rect 37436 37826 37492 37838
rect 37436 37774 37438 37826
rect 37490 37774 37492 37826
rect 37436 37268 37492 37774
rect 37436 37174 37492 37212
rect 37436 36260 37492 36270
rect 37436 36166 37492 36204
rect 37324 35700 37380 35710
rect 37324 34356 37380 35644
rect 37548 35698 37604 35710
rect 37548 35646 37550 35698
rect 37602 35646 37604 35698
rect 37436 35586 37492 35598
rect 37436 35534 37438 35586
rect 37490 35534 37492 35586
rect 37436 34916 37492 35534
rect 37548 35140 37604 35646
rect 37548 35074 37604 35084
rect 37548 34916 37604 34926
rect 37436 34914 37604 34916
rect 37436 34862 37550 34914
rect 37602 34862 37604 34914
rect 37436 34860 37604 34862
rect 37548 34850 37604 34860
rect 37324 34290 37380 34300
rect 37548 34244 37604 34254
rect 37548 34018 37604 34188
rect 37548 33966 37550 34018
rect 37602 33966 37604 34018
rect 37548 33684 37604 33966
rect 37548 33618 37604 33628
rect 37436 33348 37492 33358
rect 37436 33254 37492 33292
rect 37436 32450 37492 32462
rect 37436 32398 37438 32450
rect 37490 32398 37492 32450
rect 37436 32340 37492 32398
rect 37436 32274 37492 32284
rect 37660 31780 37716 38612
rect 37772 38612 37828 40574
rect 37996 40404 38052 41580
rect 38556 41076 38612 41086
rect 38556 40982 38612 41020
rect 37996 40338 38052 40348
rect 38444 40516 38500 40526
rect 38444 39172 38500 40460
rect 38556 40404 38612 40414
rect 38556 39730 38612 40348
rect 38556 39678 38558 39730
rect 38610 39678 38612 39730
rect 38556 39666 38612 39678
rect 38444 39116 38612 39172
rect 38332 38722 38388 38734
rect 38332 38670 38334 38722
rect 38386 38670 38388 38722
rect 38332 38668 38388 38670
rect 37772 38546 37828 38556
rect 38108 38612 38388 38668
rect 38108 38052 38164 38612
rect 38444 38610 38500 38622
rect 38444 38558 38446 38610
rect 38498 38558 38500 38610
rect 37996 38050 38164 38052
rect 37996 37998 38110 38050
rect 38162 37998 38164 38050
rect 37996 37996 38164 37998
rect 37884 36484 37940 36494
rect 37884 36390 37940 36428
rect 37548 31724 37716 31780
rect 37772 35364 37828 35374
rect 37324 31668 37380 31678
rect 37324 29764 37380 31612
rect 37436 31556 37492 31566
rect 37436 31462 37492 31500
rect 37548 30772 37604 31724
rect 37772 31668 37828 35308
rect 37996 35026 38052 37996
rect 38108 37986 38164 37996
rect 38332 38052 38388 38062
rect 38108 37828 38164 37838
rect 38108 37378 38164 37772
rect 38332 37492 38388 37996
rect 38444 37604 38500 38558
rect 38444 37538 38500 37548
rect 38332 37426 38388 37436
rect 38108 37326 38110 37378
rect 38162 37326 38164 37378
rect 38108 37314 38164 37326
rect 38332 36258 38388 36270
rect 38332 36206 38334 36258
rect 38386 36206 38388 36258
rect 38332 36036 38388 36206
rect 38332 35924 38388 35980
rect 38556 35924 38612 39116
rect 38780 38724 38836 43262
rect 38892 42980 38948 43652
rect 39116 43426 39172 43438
rect 39116 43374 39118 43426
rect 39170 43374 39172 43426
rect 39116 43314 39172 43374
rect 39116 43262 39118 43314
rect 39170 43262 39172 43314
rect 39116 43250 39172 43262
rect 38892 42924 39060 42980
rect 38892 42754 38948 42766
rect 38892 42702 38894 42754
rect 38946 42702 38948 42754
rect 38892 41972 38948 42702
rect 38892 41188 38948 41916
rect 38892 41122 38948 41132
rect 38892 40404 38948 40414
rect 38892 40310 38948 40348
rect 39004 40292 39060 42924
rect 39116 42754 39172 42766
rect 39116 42702 39118 42754
rect 39170 42702 39172 42754
rect 39116 41860 39172 42702
rect 39116 41794 39172 41804
rect 39228 41636 39284 43652
rect 39340 41858 39396 45724
rect 39452 42868 39508 45948
rect 39564 45668 39620 46622
rect 39676 46114 39732 47292
rect 40012 46786 40068 47404
rect 40348 47348 40404 47358
rect 40348 47254 40404 47292
rect 40572 47348 40628 47358
rect 40572 47254 40628 47292
rect 40012 46734 40014 46786
rect 40066 46734 40068 46786
rect 40012 46722 40068 46734
rect 40460 47124 40516 47134
rect 39676 46062 39678 46114
rect 39730 46062 39732 46114
rect 39676 46050 39732 46062
rect 40236 45780 40292 45790
rect 40236 45686 40292 45724
rect 39564 45574 39620 45612
rect 39788 45218 39844 45230
rect 39788 45166 39790 45218
rect 39842 45166 39844 45218
rect 39676 45106 39732 45118
rect 39676 45054 39678 45106
rect 39730 45054 39732 45106
rect 39676 44436 39732 45054
rect 39676 44370 39732 44380
rect 39676 44212 39732 44222
rect 39788 44212 39844 45166
rect 40012 45106 40068 45118
rect 40012 45054 40014 45106
rect 40066 45054 40068 45106
rect 39900 44436 39956 44446
rect 39900 44342 39956 44380
rect 40012 44324 40068 45054
rect 40348 44996 40404 45006
rect 40348 44902 40404 44940
rect 40236 44436 40292 44446
rect 40236 44342 40292 44380
rect 40012 44258 40068 44268
rect 39732 44156 39844 44212
rect 39676 44118 39732 44156
rect 39564 44100 39620 44110
rect 39564 43708 39620 44044
rect 39564 43652 39732 43708
rect 39676 43558 39732 43596
rect 40348 43652 40404 43662
rect 40348 43558 40404 43596
rect 40460 43428 40516 47068
rect 40572 45668 40628 45678
rect 40572 45574 40628 45612
rect 40572 44660 40628 44670
rect 40572 43708 40628 44604
rect 40572 43652 40740 43708
rect 40572 43540 40628 43550
rect 40572 43446 40628 43484
rect 40460 43362 40516 43372
rect 40460 42868 40516 42878
rect 39452 42812 39956 42868
rect 39788 42644 39844 42654
rect 39340 41806 39342 41858
rect 39394 41806 39396 41858
rect 39340 41794 39396 41806
rect 39676 41860 39732 41870
rect 39228 41580 39620 41636
rect 39564 41298 39620 41580
rect 39564 41246 39566 41298
rect 39618 41246 39620 41298
rect 39564 41234 39620 41246
rect 39452 41188 39508 41198
rect 39452 41094 39508 41132
rect 39676 41186 39732 41804
rect 39788 41858 39844 42588
rect 39788 41806 39790 41858
rect 39842 41806 39844 41858
rect 39788 41794 39844 41806
rect 39676 41134 39678 41186
rect 39730 41134 39732 41186
rect 39676 41122 39732 41134
rect 39788 41524 39844 41534
rect 39004 38668 39060 40236
rect 38780 38658 38836 38668
rect 38892 38612 39060 38668
rect 39228 40852 39284 40862
rect 39228 40402 39284 40796
rect 39228 40350 39230 40402
rect 39282 40350 39284 40402
rect 38668 37604 38724 37614
rect 38668 37378 38724 37548
rect 38780 37492 38836 37502
rect 38780 37398 38836 37436
rect 38668 37326 38670 37378
rect 38722 37326 38724 37378
rect 38668 37314 38724 37326
rect 38780 37044 38836 37054
rect 38332 35922 38612 35924
rect 38332 35870 38558 35922
rect 38610 35870 38612 35922
rect 38332 35868 38612 35870
rect 38556 35858 38612 35868
rect 38668 36932 38724 36942
rect 38108 35586 38164 35598
rect 38108 35534 38110 35586
rect 38162 35534 38164 35586
rect 38108 35140 38164 35534
rect 38108 35074 38164 35084
rect 37996 34974 37998 35026
rect 38050 34974 38052 35026
rect 37996 34962 38052 34974
rect 37884 34916 37940 34926
rect 37884 34132 37940 34860
rect 38220 34914 38276 34926
rect 38220 34862 38222 34914
rect 38274 34862 38276 34914
rect 38220 34244 38276 34862
rect 38220 34178 38276 34188
rect 38556 34580 38612 34590
rect 38108 34132 38164 34142
rect 37884 34130 38164 34132
rect 37884 34078 38110 34130
rect 38162 34078 38164 34130
rect 37884 34076 38164 34078
rect 38108 33684 38164 34076
rect 38332 34132 38388 34142
rect 38332 33908 38388 34076
rect 38108 33618 38164 33628
rect 38220 33852 38388 33908
rect 38220 32562 38276 33852
rect 38556 33460 38612 34524
rect 38556 33394 38612 33404
rect 38444 33346 38500 33358
rect 38444 33294 38446 33346
rect 38498 33294 38500 33346
rect 38444 33012 38500 33294
rect 38668 33124 38724 36876
rect 38780 36594 38836 36988
rect 38780 36542 38782 36594
rect 38834 36542 38836 36594
rect 38780 36530 38836 36542
rect 38892 35028 38948 38612
rect 39228 38274 39284 40350
rect 39228 38222 39230 38274
rect 39282 38222 39284 38274
rect 39228 38210 39284 38222
rect 39340 38722 39396 38734
rect 39340 38670 39342 38722
rect 39394 38670 39396 38722
rect 39004 38052 39060 38062
rect 39004 37958 39060 37996
rect 39228 37826 39284 37838
rect 39228 37774 39230 37826
rect 39282 37774 39284 37826
rect 39004 37604 39060 37614
rect 39004 37490 39060 37548
rect 39004 37438 39006 37490
rect 39058 37438 39060 37490
rect 39004 37426 39060 37438
rect 38892 34916 38948 34972
rect 38780 34860 38948 34916
rect 39004 35588 39060 35598
rect 38780 34802 38836 34860
rect 38780 34750 38782 34802
rect 38834 34750 38836 34802
rect 38780 34738 38836 34750
rect 39004 34802 39060 35532
rect 39116 35586 39172 35598
rect 39116 35534 39118 35586
rect 39170 35534 39172 35586
rect 39116 34916 39172 35534
rect 39228 35588 39284 37774
rect 39340 37492 39396 38670
rect 39788 38668 39844 41468
rect 39676 38612 39844 38668
rect 39900 40964 39956 42812
rect 40012 42866 40516 42868
rect 40012 42814 40462 42866
rect 40514 42814 40516 42866
rect 40012 42812 40516 42814
rect 40012 41186 40068 42812
rect 40460 42802 40516 42812
rect 40348 42644 40404 42654
rect 40348 42550 40404 42588
rect 40572 42530 40628 42542
rect 40572 42478 40574 42530
rect 40626 42478 40628 42530
rect 40124 41972 40180 41982
rect 40124 41970 40516 41972
rect 40124 41918 40126 41970
rect 40178 41918 40516 41970
rect 40124 41916 40516 41918
rect 40124 41906 40180 41916
rect 40012 41134 40014 41186
rect 40066 41134 40068 41186
rect 40012 41122 40068 41134
rect 40460 41186 40516 41916
rect 40572 41524 40628 42478
rect 40684 41748 40740 43652
rect 40796 43428 40852 43438
rect 40796 43334 40852 43372
rect 40796 42532 40852 42542
rect 40796 42438 40852 42476
rect 40908 41972 40964 50372
rect 41020 47460 41076 47470
rect 41020 47366 41076 47404
rect 41132 46452 41188 50372
rect 42028 49810 42084 49822
rect 42028 49758 42030 49810
rect 42082 49758 42084 49810
rect 41916 49698 41972 49710
rect 41916 49646 41918 49698
rect 41970 49646 41972 49698
rect 41804 48916 41860 48926
rect 41916 48916 41972 49646
rect 41860 48860 41972 48916
rect 41804 48822 41860 48860
rect 42028 48804 42084 49758
rect 42140 49252 42196 49262
rect 42252 49252 42308 51438
rect 42924 51380 42980 51390
rect 42588 50820 42644 50830
rect 42588 49698 42644 50764
rect 42924 50818 42980 51324
rect 42924 50766 42926 50818
rect 42978 50766 42980 50818
rect 42924 50596 42980 50766
rect 42924 50530 42980 50540
rect 43036 50036 43092 52894
rect 45276 51492 45332 53340
rect 46060 52274 46116 53676
rect 46172 53666 46228 53676
rect 46844 53638 46900 53676
rect 47292 53506 47348 54460
rect 48076 54450 48132 54460
rect 47516 54292 47572 54302
rect 47516 54198 47572 54236
rect 48188 53842 48244 56364
rect 50204 56308 50260 56590
rect 50204 56242 50260 56252
rect 50316 57538 50372 57550
rect 50316 57486 50318 57538
rect 50370 57486 50372 57538
rect 50204 56084 50260 56094
rect 48300 55970 48356 55982
rect 48300 55918 48302 55970
rect 48354 55918 48356 55970
rect 48300 55300 48356 55918
rect 48300 55234 48356 55244
rect 48524 55972 48580 55982
rect 48412 55188 48468 55226
rect 48412 55122 48468 55132
rect 48524 54964 48580 55916
rect 49532 55972 49588 55982
rect 49532 55878 49588 55916
rect 48300 54908 48580 54964
rect 49084 55074 49140 55086
rect 49084 55022 49086 55074
rect 49138 55022 49140 55074
rect 48300 54738 48356 54908
rect 48300 54686 48302 54738
rect 48354 54686 48356 54738
rect 48300 54292 48356 54686
rect 48412 54740 48468 54750
rect 48412 54646 48468 54684
rect 48524 54628 48580 54666
rect 48524 54562 48580 54572
rect 48748 54516 48804 54526
rect 49084 54516 49140 55022
rect 50204 54628 50260 56028
rect 50316 55970 50372 57486
rect 50540 57540 50596 57550
rect 50540 57446 50596 57484
rect 51324 57426 51380 57438
rect 51324 57374 51326 57426
rect 51378 57374 51380 57426
rect 50652 56868 50708 56878
rect 51212 56868 51268 56878
rect 51324 56868 51380 57374
rect 50652 56866 51156 56868
rect 50652 56814 50654 56866
rect 50706 56814 51156 56866
rect 50652 56812 51156 56814
rect 50652 56802 50708 56812
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 51100 56306 51156 56812
rect 51212 56866 51380 56868
rect 51212 56814 51214 56866
rect 51266 56814 51380 56866
rect 51212 56812 51380 56814
rect 51212 56802 51268 56812
rect 51436 56756 51492 58156
rect 51548 57428 51604 58270
rect 53788 57876 53844 57886
rect 51884 57652 51940 57662
rect 51884 57558 51940 57596
rect 52108 57650 52164 57662
rect 52108 57598 52110 57650
rect 52162 57598 52164 57650
rect 51996 57540 52052 57550
rect 51996 57446 52052 57484
rect 51604 57372 51940 57428
rect 51548 57296 51604 57372
rect 51100 56254 51102 56306
rect 51154 56254 51156 56306
rect 51100 56242 51156 56254
rect 51324 56700 51492 56756
rect 51660 56980 51716 56990
rect 51660 56866 51716 56924
rect 51660 56814 51662 56866
rect 51714 56814 51716 56866
rect 51212 56196 51268 56206
rect 51324 56196 51380 56700
rect 51212 56194 51380 56196
rect 51212 56142 51214 56194
rect 51266 56142 51380 56194
rect 51212 56140 51380 56142
rect 51212 56130 51268 56140
rect 51324 56084 51380 56140
rect 51324 56018 51380 56028
rect 51436 56308 51492 56318
rect 50316 55918 50318 55970
rect 50370 55918 50372 55970
rect 50316 55906 50372 55918
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 51436 54738 51492 56252
rect 51660 56084 51716 56814
rect 51772 56084 51828 56094
rect 51660 56082 51828 56084
rect 51660 56030 51774 56082
rect 51826 56030 51828 56082
rect 51660 56028 51828 56030
rect 51884 56084 51940 57372
rect 51996 57092 52052 57102
rect 51996 56978 52052 57036
rect 51996 56926 51998 56978
rect 52050 56926 52052 56978
rect 51996 56914 52052 56926
rect 52108 56868 52164 57598
rect 52108 56802 52164 56812
rect 52220 57652 52276 57662
rect 52220 56866 52276 57596
rect 52332 57650 52388 57662
rect 52332 57598 52334 57650
rect 52386 57598 52388 57650
rect 52332 56980 52388 57598
rect 53116 57538 53172 57550
rect 53116 57486 53118 57538
rect 53170 57486 53172 57538
rect 53116 57426 53172 57486
rect 53116 57374 53118 57426
rect 53170 57374 53172 57426
rect 53116 57362 53172 57374
rect 53564 57538 53620 57550
rect 53564 57486 53566 57538
rect 53618 57486 53620 57538
rect 52332 56914 52388 56924
rect 53340 56868 53396 56878
rect 52220 56814 52222 56866
rect 52274 56814 52276 56866
rect 52220 56644 52276 56814
rect 52444 56866 53396 56868
rect 52444 56814 53342 56866
rect 53394 56814 53396 56866
rect 52444 56812 53396 56814
rect 52332 56756 52388 56766
rect 52332 56662 52388 56700
rect 52220 56578 52276 56588
rect 52332 56196 52388 56206
rect 52444 56196 52500 56812
rect 53340 56802 53396 56812
rect 52332 56194 52500 56196
rect 52332 56142 52334 56194
rect 52386 56142 52500 56194
rect 52332 56140 52500 56142
rect 52892 56644 52948 56654
rect 52332 56130 52388 56140
rect 51996 56084 52052 56094
rect 51884 56082 52052 56084
rect 51884 56030 51998 56082
rect 52050 56030 52052 56082
rect 51884 56028 52052 56030
rect 51772 55468 51828 56028
rect 51996 56018 52052 56028
rect 52220 56084 52276 56094
rect 52220 55990 52276 56028
rect 52892 55970 52948 56588
rect 53564 56644 53620 57486
rect 53788 56978 53844 57820
rect 54012 57540 54068 57550
rect 53788 56926 53790 56978
rect 53842 56926 53844 56978
rect 53788 56914 53844 56926
rect 53900 57538 54068 57540
rect 53900 57486 54014 57538
rect 54066 57486 54068 57538
rect 53900 57484 54068 57486
rect 53900 57426 53956 57484
rect 54012 57474 54068 57484
rect 53900 57374 53902 57426
rect 53954 57374 53956 57426
rect 53564 56578 53620 56588
rect 53900 56756 53956 57374
rect 52892 55918 52894 55970
rect 52946 55918 52948 55970
rect 52892 55860 52948 55918
rect 53900 55972 53956 56700
rect 54124 56866 54180 56878
rect 54124 56814 54126 56866
rect 54178 56814 54180 56866
rect 53900 55878 53956 55916
rect 54012 56308 54068 56318
rect 54124 56308 54180 56814
rect 54684 56866 54740 56878
rect 54684 56814 54686 56866
rect 54738 56814 54740 56866
rect 54684 56532 54740 56814
rect 55244 56642 55300 56654
rect 55244 56590 55246 56642
rect 55298 56590 55300 56642
rect 55244 56532 55300 56590
rect 54684 56476 55300 56532
rect 54012 56306 54180 56308
rect 54012 56254 54014 56306
rect 54066 56254 54180 56306
rect 54012 56252 54180 56254
rect 52892 55794 52948 55804
rect 54012 55468 54068 56252
rect 54460 55972 54516 55982
rect 54460 55878 54516 55916
rect 55132 55972 55188 55982
rect 51772 55412 52164 55468
rect 53676 55412 53732 55422
rect 51436 54686 51438 54738
rect 51490 54686 51492 54738
rect 51436 54674 51492 54686
rect 51996 55300 52052 55310
rect 50540 54628 50596 54638
rect 50204 54626 50596 54628
rect 50204 54574 50542 54626
rect 50594 54574 50596 54626
rect 50204 54572 50596 54574
rect 50540 54562 50596 54572
rect 49868 54516 49924 54526
rect 48748 54514 49140 54516
rect 48748 54462 48750 54514
rect 48802 54462 49140 54514
rect 48748 54460 49140 54462
rect 49756 54514 49924 54516
rect 49756 54462 49870 54514
rect 49922 54462 49924 54514
rect 49756 54460 49924 54462
rect 48300 54226 48356 54236
rect 48636 54404 48692 54414
rect 48188 53790 48190 53842
rect 48242 53790 48244 53842
rect 48188 53778 48244 53790
rect 48524 53732 48580 53742
rect 48524 53638 48580 53676
rect 48188 53620 48244 53630
rect 48188 53526 48244 53564
rect 47292 53454 47294 53506
rect 47346 53454 47348 53506
rect 47292 53060 47348 53454
rect 47292 52994 47348 53004
rect 47964 53508 48020 53518
rect 47740 52836 47796 52846
rect 47740 52742 47796 52780
rect 46060 52222 46062 52274
rect 46114 52222 46116 52274
rect 46060 52210 46116 52222
rect 45724 52164 45780 52174
rect 45724 51492 45780 52108
rect 46172 52164 46228 52174
rect 46172 52070 46228 52108
rect 46620 52164 46676 52174
rect 46620 52162 46788 52164
rect 46620 52110 46622 52162
rect 46674 52110 46788 52162
rect 46620 52108 46788 52110
rect 46620 52098 46676 52108
rect 45948 52050 46004 52062
rect 45948 51998 45950 52050
rect 46002 51998 46004 52050
rect 45948 51716 46004 51998
rect 45948 51660 46116 51716
rect 45948 51492 46004 51502
rect 45276 51426 45332 51436
rect 45612 51490 46004 51492
rect 45612 51438 45950 51490
rect 46002 51438 46004 51490
rect 45612 51436 46004 51438
rect 43148 51380 43204 51390
rect 43148 51286 43204 51324
rect 44044 51380 44100 51390
rect 44044 51286 44100 51324
rect 44940 51380 44996 51390
rect 44940 51286 44996 51324
rect 43260 51266 43316 51278
rect 43260 51214 43262 51266
rect 43314 51214 43316 51266
rect 43260 50820 43316 51214
rect 43260 50754 43316 50764
rect 44156 51156 44212 51166
rect 43148 50706 43204 50718
rect 43148 50654 43150 50706
rect 43202 50654 43204 50706
rect 43148 50372 43204 50654
rect 43372 50596 43428 50606
rect 43372 50594 43652 50596
rect 43372 50542 43374 50594
rect 43426 50542 43652 50594
rect 43372 50540 43652 50542
rect 43372 50530 43428 50540
rect 43148 50316 43540 50372
rect 43260 50036 43316 50046
rect 43036 50034 43316 50036
rect 43036 49982 43262 50034
rect 43314 49982 43316 50034
rect 43036 49980 43316 49982
rect 43260 49970 43316 49980
rect 42588 49646 42590 49698
rect 42642 49646 42644 49698
rect 42588 49634 42644 49646
rect 42140 49250 42308 49252
rect 42140 49198 42142 49250
rect 42194 49198 42308 49250
rect 42140 49196 42308 49198
rect 43484 49588 43540 50316
rect 43596 49812 43652 50540
rect 43596 49746 43652 49756
rect 43820 49700 43876 49710
rect 43820 49606 43876 49644
rect 43596 49588 43652 49598
rect 43484 49586 43652 49588
rect 43484 49534 43598 49586
rect 43650 49534 43652 49586
rect 43484 49532 43652 49534
rect 42140 49186 42196 49196
rect 42028 48710 42084 48748
rect 43148 49084 43428 49140
rect 43148 48244 43204 49084
rect 42924 48242 43204 48244
rect 42924 48190 43150 48242
rect 43202 48190 43204 48242
rect 42924 48188 43204 48190
rect 42476 47572 42532 47582
rect 42476 47478 42532 47516
rect 41580 47460 41636 47470
rect 41580 47366 41636 47404
rect 41804 47458 41860 47470
rect 41804 47406 41806 47458
rect 41858 47406 41860 47458
rect 41132 45668 41188 46396
rect 41244 47348 41300 47358
rect 41244 46002 41300 47292
rect 41804 47348 41860 47406
rect 41804 47282 41860 47292
rect 41244 45950 41246 46002
rect 41298 45950 41300 46002
rect 41244 45938 41300 45950
rect 41804 46900 41860 46910
rect 41692 45892 41748 45902
rect 41132 45602 41188 45612
rect 41468 45890 41748 45892
rect 41468 45838 41694 45890
rect 41746 45838 41748 45890
rect 41468 45836 41748 45838
rect 41468 45444 41524 45836
rect 41692 45780 41748 45836
rect 41692 45714 41748 45724
rect 41468 45330 41524 45388
rect 41468 45278 41470 45330
rect 41522 45278 41524 45330
rect 41468 45266 41524 45278
rect 41356 45108 41412 45118
rect 41356 44436 41412 45052
rect 41244 44324 41300 44334
rect 41244 44230 41300 44268
rect 41356 44210 41412 44380
rect 41580 44324 41636 44334
rect 41580 44230 41636 44268
rect 41356 44158 41358 44210
rect 41410 44158 41412 44210
rect 41356 44146 41412 44158
rect 41580 43540 41636 43550
rect 41636 43484 41748 43540
rect 41580 43408 41636 43484
rect 41356 42532 41412 42542
rect 41412 42476 41524 42532
rect 41356 42400 41412 42476
rect 40908 41906 40964 41916
rect 41468 41858 41524 42476
rect 41468 41806 41470 41858
rect 41522 41806 41524 41858
rect 40684 41692 40964 41748
rect 40572 41468 40852 41524
rect 40460 41134 40462 41186
rect 40514 41134 40516 41186
rect 40460 41122 40516 41134
rect 40796 41074 40852 41468
rect 40796 41022 40798 41074
rect 40850 41022 40852 41074
rect 39900 40290 39956 40908
rect 40684 40962 40740 40974
rect 40684 40910 40686 40962
rect 40738 40910 40740 40962
rect 40684 40628 40740 40910
rect 40684 40562 40740 40572
rect 40012 40516 40068 40526
rect 40012 40402 40068 40460
rect 40012 40350 40014 40402
rect 40066 40350 40068 40402
rect 40012 40338 40068 40350
rect 39900 40238 39902 40290
rect 39954 40238 39956 40290
rect 39564 38050 39620 38062
rect 39564 37998 39566 38050
rect 39618 37998 39620 38050
rect 39564 37604 39620 37998
rect 39676 37716 39732 38612
rect 39900 38500 39956 40238
rect 40236 40180 40292 40190
rect 40236 40086 40292 40124
rect 40796 40180 40852 41022
rect 40796 40114 40852 40124
rect 40460 39732 40516 39742
rect 40460 39638 40516 39676
rect 40796 38948 40852 38958
rect 40796 38854 40852 38892
rect 40124 38834 40180 38846
rect 40124 38782 40126 38834
rect 40178 38782 40180 38834
rect 40124 38668 40180 38782
rect 40348 38724 40404 38734
rect 39676 37650 39732 37660
rect 39788 38444 39956 38500
rect 40012 38612 40180 38668
rect 40236 38722 40404 38724
rect 40236 38670 40350 38722
rect 40402 38670 40404 38722
rect 40236 38668 40404 38670
rect 39564 37538 39620 37548
rect 39788 37492 39844 38444
rect 40012 37826 40068 38612
rect 40124 38164 40180 38174
rect 40124 38070 40180 38108
rect 40236 38052 40292 38668
rect 40348 38658 40404 38668
rect 40908 38164 40964 41692
rect 41244 40964 41300 40974
rect 41244 40870 41300 40908
rect 41468 40628 41524 41806
rect 41468 40562 41524 40572
rect 41132 40180 41188 40190
rect 41132 39730 41188 40124
rect 41132 39678 41134 39730
rect 41186 39678 41188 39730
rect 41132 39666 41188 39678
rect 41580 39620 41636 39630
rect 41580 39526 41636 39564
rect 41692 39396 41748 43484
rect 41804 43316 41860 46844
rect 42588 46562 42644 46574
rect 42588 46510 42590 46562
rect 42642 46510 42644 46562
rect 42140 45892 42196 45902
rect 41804 43250 41860 43260
rect 41916 45836 42140 45892
rect 41804 42532 41860 42542
rect 41804 42438 41860 42476
rect 41804 40964 41860 40974
rect 41804 40870 41860 40908
rect 41916 40404 41972 45836
rect 42140 45798 42196 45836
rect 42588 45780 42644 46510
rect 42812 45892 42868 45902
rect 42812 45798 42868 45836
rect 42588 45714 42644 45724
rect 42476 45668 42532 45678
rect 42252 45108 42308 45118
rect 42252 45014 42308 45052
rect 42028 44098 42084 44110
rect 42028 44046 42030 44098
rect 42082 44046 42084 44098
rect 42028 43708 42084 44046
rect 42028 43652 42420 43708
rect 42028 41524 42084 43652
rect 42252 43540 42308 43550
rect 42028 41458 42084 41468
rect 42140 42420 42196 42430
rect 42140 41746 42196 42364
rect 42252 42196 42308 43484
rect 42364 43426 42420 43652
rect 42364 43374 42366 43426
rect 42418 43374 42420 43426
rect 42364 43362 42420 43374
rect 42252 42130 42308 42140
rect 42364 42532 42420 42542
rect 42140 41694 42142 41746
rect 42194 41694 42196 41746
rect 42140 40962 42196 41694
rect 42140 40910 42142 40962
rect 42194 40910 42196 40962
rect 42140 40852 42196 40910
rect 42140 40786 42196 40796
rect 42364 42082 42420 42476
rect 42476 42420 42532 45612
rect 42812 45332 42868 45342
rect 42924 45332 42980 48188
rect 43148 48178 43204 48188
rect 43260 48914 43316 48926
rect 43260 48862 43262 48914
rect 43314 48862 43316 48914
rect 43260 48132 43316 48862
rect 43372 48914 43428 49084
rect 43372 48862 43374 48914
rect 43426 48862 43428 48914
rect 43372 48850 43428 48862
rect 43372 48132 43428 48142
rect 43260 48130 43428 48132
rect 43260 48078 43374 48130
rect 43426 48078 43428 48130
rect 43260 48076 43428 48078
rect 43260 47572 43316 48076
rect 43372 48066 43428 48076
rect 43260 47506 43316 47516
rect 43148 46116 43204 46126
rect 43484 46116 43540 49532
rect 43596 49522 43652 49532
rect 43820 48916 43876 48926
rect 43596 48804 43652 48814
rect 43596 48710 43652 48748
rect 43820 48354 43876 48860
rect 43820 48302 43822 48354
rect 43874 48302 43876 48354
rect 43820 48290 43876 48302
rect 43148 46114 43540 46116
rect 43148 46062 43150 46114
rect 43202 46062 43540 46114
rect 43148 46060 43540 46062
rect 44044 47458 44100 47470
rect 44044 47406 44046 47458
rect 44098 47406 44100 47458
rect 44044 47348 44100 47406
rect 43148 46050 43204 46060
rect 43036 45780 43092 45790
rect 43036 45686 43092 45724
rect 42812 45330 42980 45332
rect 42812 45278 42814 45330
rect 42866 45278 42980 45330
rect 42812 45276 42980 45278
rect 42812 45266 42868 45276
rect 43596 45220 43652 45230
rect 42700 45106 42756 45118
rect 42700 45054 42702 45106
rect 42754 45054 42756 45106
rect 42588 44324 42644 44334
rect 42700 44324 42756 45054
rect 42924 45106 42980 45118
rect 42924 45054 42926 45106
rect 42978 45054 42980 45106
rect 42812 44324 42868 44334
rect 42700 44322 42868 44324
rect 42700 44270 42814 44322
rect 42866 44270 42868 44322
rect 42700 44268 42868 44270
rect 42588 44230 42644 44268
rect 42812 43314 42868 44268
rect 42924 44324 42980 45054
rect 42924 44258 42980 44268
rect 43484 44212 43540 44222
rect 43484 44118 43540 44156
rect 43596 43764 43652 45164
rect 43596 43698 43652 43708
rect 43932 43650 43988 43662
rect 43932 43598 43934 43650
rect 43986 43598 43988 43650
rect 43932 43540 43988 43598
rect 43932 43474 43988 43484
rect 44044 43426 44100 47292
rect 44156 45668 44212 51100
rect 45052 51156 45108 51166
rect 45052 51062 45108 51100
rect 44604 50372 44660 50382
rect 44604 49250 44660 50316
rect 44604 49198 44606 49250
rect 44658 49198 44660 49250
rect 44604 49186 44660 49198
rect 45164 49700 45220 49710
rect 44716 49028 44772 49038
rect 44716 48934 44772 48972
rect 44604 48804 44660 48814
rect 44604 48710 44660 48748
rect 44604 47460 44660 47470
rect 44604 47366 44660 47404
rect 44716 47346 44772 47358
rect 44716 47294 44718 47346
rect 44770 47294 44772 47346
rect 44716 46788 44772 47294
rect 44716 46722 44772 46732
rect 44716 46004 44772 46014
rect 44156 45574 44212 45612
rect 44380 46002 44772 46004
rect 44380 45950 44718 46002
rect 44770 45950 44772 46002
rect 44380 45948 44772 45950
rect 44380 45444 44436 45948
rect 44716 45938 44772 45948
rect 45164 45892 45220 49644
rect 45612 47570 45668 51436
rect 45948 51426 46004 51436
rect 45836 51266 45892 51278
rect 45836 51214 45838 51266
rect 45890 51214 45892 51266
rect 45836 50372 45892 51214
rect 46060 50706 46116 51660
rect 46284 51156 46340 51166
rect 46284 50818 46340 51100
rect 46284 50766 46286 50818
rect 46338 50766 46340 50818
rect 46284 50754 46340 50766
rect 46060 50654 46062 50706
rect 46114 50654 46116 50706
rect 46060 50642 46116 50654
rect 46732 50594 46788 52108
rect 47404 51492 47460 51502
rect 47180 51380 47236 51390
rect 47180 51286 47236 51324
rect 46732 50542 46734 50594
rect 46786 50542 46788 50594
rect 46732 50530 46788 50542
rect 47068 51156 47124 51166
rect 47068 50594 47124 51100
rect 47068 50542 47070 50594
rect 47122 50542 47124 50594
rect 47068 50530 47124 50542
rect 47404 50596 47460 51436
rect 47852 51492 47908 51502
rect 47964 51492 48020 53452
rect 47852 51490 48020 51492
rect 47852 51438 47854 51490
rect 47906 51438 48020 51490
rect 47852 51436 48020 51438
rect 48636 52836 48692 54348
rect 48748 53956 48804 54460
rect 49756 54068 49812 54460
rect 49868 54450 49924 54460
rect 51212 54516 51268 54526
rect 51212 54514 51380 54516
rect 51212 54462 51214 54514
rect 51266 54462 51380 54514
rect 51212 54460 51380 54462
rect 51212 54450 51268 54460
rect 48748 53890 48804 53900
rect 49420 54012 49812 54068
rect 50092 54402 50148 54414
rect 50092 54350 50094 54402
rect 50146 54350 50148 54402
rect 49420 53730 49476 54012
rect 49420 53678 49422 53730
rect 49474 53678 49476 53730
rect 49420 53666 49476 53678
rect 50092 53732 50148 54350
rect 50092 53666 50148 53676
rect 51324 53730 51380 54460
rect 51324 53678 51326 53730
rect 51378 53678 51380 53730
rect 47852 51426 47908 51436
rect 45836 50306 45892 50316
rect 46060 50372 46116 50382
rect 46060 50278 46116 50316
rect 46956 50372 47012 50382
rect 46956 50278 47012 50316
rect 45948 50036 46004 50046
rect 45948 50034 46452 50036
rect 45948 49982 45950 50034
rect 46002 49982 46452 50034
rect 45948 49980 46452 49982
rect 45948 49970 46004 49980
rect 45724 49810 45780 49822
rect 45724 49758 45726 49810
rect 45778 49758 45780 49810
rect 45724 49028 45780 49758
rect 45724 48962 45780 48972
rect 46060 49810 46116 49822
rect 46060 49758 46062 49810
rect 46114 49758 46116 49810
rect 46060 48916 46116 49758
rect 46396 49028 46452 49980
rect 47180 49252 47236 49262
rect 47180 49158 47236 49196
rect 46732 49138 46788 49150
rect 46732 49086 46734 49138
rect 46786 49086 46788 49138
rect 46396 49026 46676 49028
rect 46396 48974 46398 49026
rect 46450 48974 46676 49026
rect 46396 48972 46676 48974
rect 46396 48962 46452 48972
rect 46060 48850 46116 48860
rect 46620 48354 46676 48972
rect 46732 48916 46788 49086
rect 46732 48850 46788 48860
rect 46620 48302 46622 48354
rect 46674 48302 46676 48354
rect 46620 48290 46676 48302
rect 46172 48244 46228 48254
rect 46172 48150 46228 48188
rect 46508 48242 46564 48254
rect 46508 48190 46510 48242
rect 46562 48190 46564 48242
rect 45612 47518 45614 47570
rect 45666 47518 45668 47570
rect 45612 47506 45668 47518
rect 46060 47572 46116 47582
rect 45388 47460 45444 47470
rect 44156 45388 44436 45444
rect 44492 45780 44548 45790
rect 44156 45218 44212 45388
rect 44492 45330 44548 45724
rect 44492 45278 44494 45330
rect 44546 45278 44548 45330
rect 44492 45266 44548 45278
rect 45052 45444 45108 45454
rect 45052 45330 45108 45388
rect 45052 45278 45054 45330
rect 45106 45278 45108 45330
rect 45052 45266 45108 45278
rect 45164 45330 45220 45836
rect 45164 45278 45166 45330
rect 45218 45278 45220 45330
rect 45164 45266 45220 45278
rect 45276 47012 45332 47022
rect 44156 45166 44158 45218
rect 44210 45166 44212 45218
rect 44156 44322 44212 45166
rect 44268 45220 44324 45230
rect 44324 45164 44436 45220
rect 44268 45126 44324 45164
rect 44268 44436 44324 44446
rect 44268 44342 44324 44380
rect 44156 44270 44158 44322
rect 44210 44270 44212 44322
rect 44156 43708 44212 44270
rect 44380 44322 44436 45164
rect 45276 45108 45332 46956
rect 45388 46004 45444 47404
rect 46060 47458 46116 47516
rect 46060 47406 46062 47458
rect 46114 47406 46116 47458
rect 46060 47394 46116 47406
rect 45836 47348 45892 47358
rect 46508 47348 46564 48190
rect 46844 48244 46900 48254
rect 46732 47572 46788 47582
rect 46732 47478 46788 47516
rect 46620 47348 46676 47358
rect 46844 47348 46900 48188
rect 45836 47254 45892 47292
rect 46172 47346 46676 47348
rect 46172 47294 46622 47346
rect 46674 47294 46676 47346
rect 46172 47292 46676 47294
rect 46172 47068 46228 47292
rect 46620 47282 46676 47292
rect 46732 47346 46900 47348
rect 46732 47294 46846 47346
rect 46898 47294 46900 47346
rect 46732 47292 46900 47294
rect 45612 47012 46228 47068
rect 45612 46898 45668 47012
rect 45612 46846 45614 46898
rect 45666 46846 45668 46898
rect 45612 46834 45668 46846
rect 45500 46788 45556 46798
rect 45500 46694 45556 46732
rect 46732 46114 46788 47292
rect 46844 47282 46900 47292
rect 47180 47124 47236 47134
rect 47068 46564 47124 46574
rect 47180 46564 47236 47068
rect 47068 46562 47236 46564
rect 47068 46510 47070 46562
rect 47122 46510 47236 46562
rect 47068 46508 47236 46510
rect 47068 46498 47124 46508
rect 46732 46062 46734 46114
rect 46786 46062 46788 46114
rect 46732 46050 46788 46062
rect 45612 46004 45668 46014
rect 45388 46002 45668 46004
rect 45388 45950 45614 46002
rect 45666 45950 45668 46002
rect 45388 45948 45668 45950
rect 45612 45938 45668 45948
rect 45724 45890 45780 45902
rect 45724 45838 45726 45890
rect 45778 45838 45780 45890
rect 45500 45780 45556 45790
rect 45500 45686 45556 45724
rect 44380 44270 44382 44322
rect 44434 44270 44436 44322
rect 44380 43764 44436 44270
rect 45164 45052 45332 45108
rect 45724 45444 45780 45838
rect 45948 45892 46004 45902
rect 45948 45798 46004 45836
rect 44716 44210 44772 44222
rect 44716 44158 44718 44210
rect 44770 44158 44772 44210
rect 44604 44100 44660 44110
rect 44492 43764 44548 43774
rect 44380 43762 44548 43764
rect 44380 43710 44494 43762
rect 44546 43710 44548 43762
rect 44380 43708 44548 43710
rect 44156 43652 44324 43708
rect 44492 43698 44548 43708
rect 44044 43374 44046 43426
rect 44098 43374 44100 43426
rect 44044 43362 44100 43374
rect 42812 43262 42814 43314
rect 42866 43262 42868 43314
rect 42812 43250 42868 43262
rect 43708 43314 43764 43326
rect 43708 43262 43710 43314
rect 43762 43262 43764 43314
rect 42476 42354 42532 42364
rect 42700 42530 42756 42542
rect 43372 42532 43428 42542
rect 43708 42532 43764 43262
rect 44268 43314 44324 43652
rect 44268 43262 44270 43314
rect 44322 43262 44324 43314
rect 44268 43250 44324 43262
rect 44604 42756 44660 44044
rect 44716 43652 44772 44158
rect 44716 43586 44772 43596
rect 44940 43428 44996 43438
rect 44940 43426 45108 43428
rect 44940 43374 44942 43426
rect 44994 43374 45108 43426
rect 44940 43372 45108 43374
rect 44940 43362 44996 43372
rect 45052 43314 45108 43372
rect 45052 43262 45054 43314
rect 45106 43262 45108 43314
rect 44604 42700 44996 42756
rect 42700 42478 42702 42530
rect 42754 42478 42756 42530
rect 42700 42420 42756 42478
rect 42700 42354 42756 42364
rect 43260 42530 43764 42532
rect 43260 42478 43374 42530
rect 43426 42478 43764 42530
rect 43260 42476 43764 42478
rect 44716 42532 44772 42542
rect 42364 42030 42366 42082
rect 42418 42030 42420 42082
rect 42140 40404 42196 40414
rect 42364 40404 42420 42030
rect 43148 41860 43204 41870
rect 43148 41766 43204 41804
rect 42476 41748 42532 41758
rect 43036 41748 43092 41758
rect 42476 41746 43092 41748
rect 42476 41694 42478 41746
rect 42530 41694 43038 41746
rect 43090 41694 43092 41746
rect 42476 41692 43092 41694
rect 42476 41682 42532 41692
rect 43036 41682 43092 41692
rect 43260 41524 43316 42476
rect 43372 42466 43428 42476
rect 44716 42438 44772 42476
rect 44716 42196 44772 42206
rect 43932 42194 44772 42196
rect 43932 42142 44718 42194
rect 44770 42142 44772 42194
rect 43932 42140 44772 42142
rect 43372 41972 43428 42010
rect 43372 41906 43428 41916
rect 43260 41458 43316 41468
rect 43820 41860 43876 41870
rect 43820 41300 43876 41804
rect 43820 41234 43876 41244
rect 43932 41186 43988 42140
rect 44716 42130 44772 42140
rect 44604 41970 44660 41982
rect 44604 41918 44606 41970
rect 44658 41918 44660 41970
rect 44492 41412 44548 41422
rect 44604 41412 44660 41918
rect 44940 41970 44996 42700
rect 44940 41918 44942 41970
rect 44994 41918 44996 41970
rect 44940 41906 44996 41918
rect 44492 41410 44660 41412
rect 44492 41358 44494 41410
rect 44546 41358 44660 41410
rect 44492 41356 44660 41358
rect 44492 41346 44548 41356
rect 43932 41134 43934 41186
rect 43986 41134 43988 41186
rect 43932 41122 43988 41134
rect 43596 41076 43652 41086
rect 44380 41076 44436 41086
rect 43596 40982 43652 41020
rect 44156 41074 44436 41076
rect 44156 41022 44382 41074
rect 44434 41022 44436 41074
rect 44156 41020 44436 41022
rect 42700 40962 42756 40974
rect 42700 40910 42702 40962
rect 42754 40910 42756 40962
rect 42700 40740 42756 40910
rect 42700 40674 42756 40684
rect 43036 40964 43092 40974
rect 41916 40348 42084 40404
rect 42028 39730 42084 40348
rect 42028 39678 42030 39730
rect 42082 39678 42084 39730
rect 42028 39666 42084 39678
rect 42140 40402 42420 40404
rect 42140 40350 42142 40402
rect 42194 40350 42420 40402
rect 42140 40348 42420 40350
rect 42476 40628 42532 40638
rect 42588 40628 42644 40638
rect 42532 40626 42644 40628
rect 42532 40574 42590 40626
rect 42642 40574 42644 40626
rect 42532 40572 42644 40574
rect 42140 39732 42196 40348
rect 42140 39666 42196 39676
rect 40908 38098 40964 38108
rect 41580 39340 41748 39396
rect 40236 37920 40292 37996
rect 40796 37828 40852 37838
rect 40012 37774 40014 37826
rect 40066 37774 40068 37826
rect 39340 37426 39396 37436
rect 39676 37436 39844 37492
rect 39900 37492 39956 37502
rect 39676 37268 39732 37436
rect 39228 35522 39284 35532
rect 39340 37212 39732 37268
rect 39788 37266 39844 37278
rect 39788 37214 39790 37266
rect 39842 37214 39844 37266
rect 39116 34850 39172 34860
rect 39004 34750 39006 34802
rect 39058 34750 39060 34802
rect 38892 34690 38948 34702
rect 38892 34638 38894 34690
rect 38946 34638 38948 34690
rect 38892 34468 38948 34638
rect 39004 34692 39060 34750
rect 39004 34626 39060 34636
rect 38892 34412 39284 34468
rect 39228 34242 39284 34412
rect 39228 34190 39230 34242
rect 39282 34190 39284 34242
rect 39228 34178 39284 34190
rect 39340 34020 39396 37212
rect 39676 37044 39732 37054
rect 39676 36482 39732 36988
rect 39676 36430 39678 36482
rect 39730 36430 39732 36482
rect 39676 36418 39732 36430
rect 39564 36372 39620 36382
rect 39564 35700 39620 36316
rect 39788 36370 39844 37214
rect 39900 37154 39956 37436
rect 39900 37102 39902 37154
rect 39954 37102 39956 37154
rect 39900 37044 39956 37102
rect 39900 36978 39956 36988
rect 40012 36482 40068 37774
rect 40684 37826 40852 37828
rect 40684 37774 40798 37826
rect 40850 37774 40852 37826
rect 40684 37772 40852 37774
rect 40012 36430 40014 36482
rect 40066 36430 40068 36482
rect 40012 36418 40068 36430
rect 40236 37716 40292 37726
rect 39788 36318 39790 36370
rect 39842 36318 39844 36370
rect 39788 36148 39844 36318
rect 39676 36092 39844 36148
rect 39900 36260 39956 36270
rect 39676 35922 39732 36092
rect 39676 35870 39678 35922
rect 39730 35870 39732 35922
rect 39676 35858 39732 35870
rect 39900 35700 39956 36204
rect 39564 35644 39732 35700
rect 39564 35476 39620 35486
rect 39564 35382 39620 35420
rect 39564 34690 39620 34702
rect 39564 34638 39566 34690
rect 39618 34638 39620 34690
rect 39452 34132 39508 34142
rect 39452 34038 39508 34076
rect 39116 33964 39396 34020
rect 39116 33572 39172 33964
rect 39116 33440 39172 33516
rect 39340 33796 39396 33806
rect 39004 33236 39060 33246
rect 38668 33068 38836 33124
rect 38444 32956 38724 33012
rect 38332 32676 38388 32686
rect 38332 32582 38388 32620
rect 38220 32510 38222 32562
rect 38274 32510 38276 32562
rect 37772 31602 37828 31612
rect 38108 32004 38164 32014
rect 37660 31554 37716 31566
rect 37660 31502 37662 31554
rect 37714 31502 37716 31554
rect 37660 31444 37716 31502
rect 38108 31444 38164 31948
rect 37660 31378 37716 31388
rect 37884 31388 38164 31444
rect 37660 30884 37716 30894
rect 37660 30882 37828 30884
rect 37660 30830 37662 30882
rect 37714 30830 37828 30882
rect 37660 30828 37828 30830
rect 37660 30818 37716 30828
rect 37324 29698 37380 29708
rect 37436 30716 37604 30772
rect 37436 29540 37492 30716
rect 36876 26852 37044 26908
rect 36988 26292 37044 26852
rect 36876 26178 36932 26190
rect 36876 26126 36878 26178
rect 36930 26126 36932 26178
rect 36876 26066 36932 26126
rect 36876 26014 36878 26066
rect 36930 26014 36932 26066
rect 36876 26002 36932 26014
rect 36988 25620 37044 26236
rect 36988 25554 37044 25564
rect 37100 26852 37268 26908
rect 37324 28756 37380 28766
rect 36764 24332 36932 24388
rect 36764 23828 36820 23838
rect 36764 23734 36820 23772
rect 36876 23716 36932 24332
rect 36876 23650 36932 23660
rect 36764 23604 36820 23614
rect 36764 23266 36820 23548
rect 37100 23492 37156 26852
rect 36764 23214 36766 23266
rect 36818 23214 36820 23266
rect 36764 23202 36820 23214
rect 36876 23436 37156 23492
rect 37212 26516 37268 26526
rect 36876 23044 36932 23436
rect 36988 23268 37044 23278
rect 36988 23174 37044 23212
rect 37212 23266 37268 26460
rect 37324 26516 37380 28700
rect 37436 28754 37492 29484
rect 37436 28702 37438 28754
rect 37490 28702 37492 28754
rect 37436 28690 37492 28702
rect 37548 30098 37604 30110
rect 37548 30046 37550 30098
rect 37602 30046 37604 30098
rect 37548 29314 37604 30046
rect 37772 29986 37828 30828
rect 37884 30434 37940 31388
rect 38220 31332 38276 32510
rect 38556 32564 38612 32574
rect 38556 32470 38612 32508
rect 38444 32452 38500 32462
rect 38220 31266 38276 31276
rect 38332 31444 38388 31454
rect 38108 31220 38164 31230
rect 38108 31126 38164 31164
rect 37884 30382 37886 30434
rect 37938 30382 37940 30434
rect 37884 30370 37940 30382
rect 38332 30324 38388 31388
rect 38332 30258 38388 30268
rect 37772 29934 37774 29986
rect 37826 29934 37828 29986
rect 37772 29426 37828 29934
rect 37772 29374 37774 29426
rect 37826 29374 37828 29426
rect 37772 29362 37828 29374
rect 37884 29652 37940 29662
rect 37548 29262 37550 29314
rect 37602 29262 37604 29314
rect 37548 28420 37604 29262
rect 37884 28754 37940 29596
rect 38220 29316 38276 29326
rect 38220 28868 38276 29260
rect 38332 29204 38388 29214
rect 38332 29110 38388 29148
rect 38220 28812 38388 28868
rect 37884 28702 37886 28754
rect 37938 28702 37940 28754
rect 37884 28690 37940 28702
rect 38332 28754 38388 28812
rect 38332 28702 38334 28754
rect 38386 28702 38388 28754
rect 38332 28690 38388 28702
rect 38220 28644 38276 28654
rect 37548 28354 37604 28364
rect 38108 28532 38164 28542
rect 38108 28082 38164 28476
rect 38108 28030 38110 28082
rect 38162 28030 38164 28082
rect 37660 27970 37716 27982
rect 37660 27918 37662 27970
rect 37714 27918 37716 27970
rect 37660 27524 37716 27918
rect 37660 27076 37716 27468
rect 37772 27076 37828 27086
rect 37660 27074 37828 27076
rect 37660 27022 37774 27074
rect 37826 27022 37828 27074
rect 37660 27020 37828 27022
rect 37772 26908 37828 27020
rect 37772 26852 38052 26908
rect 37772 26516 37828 26526
rect 37324 26514 37828 26516
rect 37324 26462 37326 26514
rect 37378 26462 37774 26514
rect 37826 26462 37828 26514
rect 37324 26460 37828 26462
rect 37324 26450 37380 26460
rect 37772 26450 37828 26460
rect 37436 25620 37492 25630
rect 37436 25526 37492 25564
rect 37884 25396 37940 25406
rect 37884 25302 37940 25340
rect 37436 24722 37492 24734
rect 37436 24670 37438 24722
rect 37490 24670 37492 24722
rect 37324 24610 37380 24622
rect 37324 24558 37326 24610
rect 37378 24558 37380 24610
rect 37324 23492 37380 24558
rect 37324 23426 37380 23436
rect 37436 23716 37492 24670
rect 37772 24500 37828 24510
rect 37772 24052 37828 24444
rect 37996 24164 38052 26852
rect 38108 26514 38164 28030
rect 38108 26462 38110 26514
rect 38162 26462 38164 26514
rect 38108 26450 38164 26462
rect 37996 24108 38164 24164
rect 37772 23958 37828 23996
rect 37548 23940 37604 23950
rect 37548 23846 37604 23884
rect 37996 23938 38052 23950
rect 37996 23886 37998 23938
rect 38050 23886 38052 23938
rect 37996 23716 38052 23886
rect 37436 23660 38052 23716
rect 37212 23214 37214 23266
rect 37266 23214 37268 23266
rect 37212 23202 37268 23214
rect 37100 23044 37156 23054
rect 37436 23044 37492 23660
rect 36876 22988 37044 23044
rect 36540 22372 36596 22382
rect 36540 22146 36596 22316
rect 36540 22094 36542 22146
rect 36594 22094 36596 22146
rect 36540 21924 36596 22094
rect 36540 21868 36932 21924
rect 36764 21700 36820 21710
rect 36092 20578 36260 20580
rect 36092 20526 36094 20578
rect 36146 20526 36260 20578
rect 36092 20524 36260 20526
rect 36316 21420 36484 21476
rect 36540 21586 36596 21598
rect 36540 21534 36542 21586
rect 36594 21534 36596 21586
rect 35756 19796 35812 19806
rect 35756 19346 35812 19740
rect 36092 19796 36148 20524
rect 36092 19730 36148 19740
rect 35756 19294 35758 19346
rect 35810 19294 35812 19346
rect 35756 19282 35812 19294
rect 36204 19236 36260 19246
rect 36316 19236 36372 21420
rect 36540 20580 36596 21534
rect 36652 21474 36708 21486
rect 36652 21422 36654 21474
rect 36706 21422 36708 21474
rect 36652 20804 36708 21422
rect 36764 21140 36820 21644
rect 36764 20914 36820 21084
rect 36764 20862 36766 20914
rect 36818 20862 36820 20914
rect 36764 20850 36820 20862
rect 36652 20738 36708 20748
rect 36540 20132 36596 20524
rect 36428 20018 36484 20030
rect 36428 19966 36430 20018
rect 36482 19966 36484 20018
rect 36428 19796 36484 19966
rect 36428 19730 36484 19740
rect 36540 19348 36596 20076
rect 36764 20132 36820 20142
rect 36764 20038 36820 20076
rect 36876 20020 36932 21868
rect 36876 19954 36932 19964
rect 36540 19292 36820 19348
rect 36260 19180 36372 19236
rect 36204 19142 36260 19180
rect 36652 19122 36708 19134
rect 36652 19070 36654 19122
rect 36706 19070 36708 19122
rect 35644 18508 36036 18564
rect 35196 18396 35812 18452
rect 35756 18338 35812 18396
rect 35756 18286 35758 18338
rect 35810 18286 35812 18338
rect 35756 18274 35812 18286
rect 34972 18174 34974 18226
rect 35026 18174 35028 18226
rect 34972 18162 35028 18174
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35868 17668 35924 17678
rect 35756 17612 35868 17668
rect 35980 17668 36036 18508
rect 36092 18452 36148 18462
rect 36092 18358 36148 18396
rect 36540 18338 36596 18350
rect 36540 18286 36542 18338
rect 36594 18286 36596 18338
rect 36540 18226 36596 18286
rect 36540 18174 36542 18226
rect 36594 18174 36596 18226
rect 36540 18162 36596 18174
rect 36652 17892 36708 19070
rect 36652 17826 36708 17836
rect 36092 17668 36148 17678
rect 35980 17666 36148 17668
rect 35980 17614 36094 17666
rect 36146 17614 36148 17666
rect 35980 17612 36148 17614
rect 35084 17556 35140 17566
rect 34860 17154 34916 17164
rect 34972 17554 35140 17556
rect 34972 17502 35086 17554
rect 35138 17502 35140 17554
rect 34972 17500 35140 17502
rect 34748 17054 34750 17106
rect 34802 17054 34804 17106
rect 34748 16436 34804 17054
rect 34748 16380 34916 16436
rect 34748 16212 34804 16222
rect 34748 16118 34804 16156
rect 34524 15486 34526 15538
rect 34578 15486 34580 15538
rect 34524 15474 34580 15486
rect 34860 15428 34916 16380
rect 34860 15362 34916 15372
rect 34972 14644 35028 17500
rect 35084 17490 35140 17500
rect 35308 17556 35364 17566
rect 35084 17108 35140 17118
rect 35084 15540 35140 17052
rect 35308 16882 35364 17500
rect 35644 17556 35700 17566
rect 35644 17462 35700 17500
rect 35644 16996 35700 17006
rect 35756 16996 35812 17612
rect 35868 17574 35924 17612
rect 35980 17444 36036 17454
rect 35980 17350 36036 17388
rect 36092 17108 36148 17612
rect 36092 17042 36148 17052
rect 36316 17666 36372 17678
rect 36316 17614 36318 17666
rect 36370 17614 36372 17666
rect 35644 16994 36036 16996
rect 35644 16942 35646 16994
rect 35698 16942 36036 16994
rect 35644 16940 36036 16942
rect 35644 16930 35700 16940
rect 35308 16830 35310 16882
rect 35362 16830 35364 16882
rect 35308 16818 35364 16830
rect 35532 16884 35588 16922
rect 35532 16818 35588 16828
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35420 16212 35476 16222
rect 35420 15986 35476 16156
rect 35756 16100 35812 16110
rect 35420 15934 35422 15986
rect 35474 15934 35476 15986
rect 35196 15540 35252 15550
rect 35084 15538 35252 15540
rect 35084 15486 35198 15538
rect 35250 15486 35252 15538
rect 35084 15484 35252 15486
rect 35196 15474 35252 15484
rect 34860 14588 35028 14644
rect 35084 15316 35140 15326
rect 35084 14754 35140 15260
rect 35420 15092 35476 15934
rect 35644 15986 35700 15998
rect 35644 15934 35646 15986
rect 35698 15934 35700 15986
rect 35644 15876 35700 15934
rect 35644 15810 35700 15820
rect 35756 15148 35812 16044
rect 35980 16098 36036 16940
rect 35980 16046 35982 16098
rect 36034 16046 36036 16098
rect 35980 16034 36036 16046
rect 36092 16658 36148 16670
rect 36092 16606 36094 16658
rect 36146 16606 36148 16658
rect 35868 15874 35924 15886
rect 35868 15822 35870 15874
rect 35922 15822 35924 15874
rect 35868 15428 35924 15822
rect 35868 15314 35924 15372
rect 35868 15262 35870 15314
rect 35922 15262 35924 15314
rect 35868 15250 35924 15262
rect 35980 15540 36036 15550
rect 35980 15314 36036 15484
rect 35980 15262 35982 15314
rect 36034 15262 36036 15314
rect 35980 15250 36036 15262
rect 36092 15316 36148 16606
rect 36204 16660 36260 16670
rect 36204 15540 36260 16604
rect 36316 15652 36372 17614
rect 36764 17556 36820 19292
rect 36764 17462 36820 17500
rect 36540 16996 36596 17006
rect 36540 16902 36596 16940
rect 36428 15988 36484 15998
rect 36428 15894 36484 15932
rect 36316 15596 36484 15652
rect 36204 15474 36260 15484
rect 36204 15316 36260 15326
rect 36092 15260 36204 15316
rect 36204 15184 36260 15260
rect 35756 15092 36036 15148
rect 35420 15026 35476 15036
rect 35756 14980 35812 14990
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35084 14702 35086 14754
rect 35138 14702 35140 14754
rect 34524 14532 34580 14542
rect 34524 14438 34580 14476
rect 34636 13860 34692 13870
rect 34636 13766 34692 13804
rect 33964 12350 33966 12402
rect 34018 12350 34020 12402
rect 33964 12338 34020 12350
rect 34188 13020 34468 13076
rect 34636 13636 34692 13646
rect 33852 11954 33908 11966
rect 33852 11902 33854 11954
rect 33906 11902 33908 11954
rect 33852 11394 33908 11902
rect 33852 11342 33854 11394
rect 33906 11342 33908 11394
rect 33852 11330 33908 11342
rect 34188 11396 34244 13020
rect 34412 12852 34468 12862
rect 34188 11264 34244 11340
rect 34300 12850 34468 12852
rect 34300 12798 34414 12850
rect 34466 12798 34468 12850
rect 34300 12796 34468 12798
rect 33740 10994 33796 11004
rect 33964 11170 34020 11182
rect 33964 11118 33966 11170
rect 34018 11118 34020 11170
rect 33964 10836 34020 11118
rect 33628 10834 34020 10836
rect 33628 10782 33630 10834
rect 33682 10782 34020 10834
rect 33628 10780 34020 10782
rect 34076 11170 34132 11182
rect 34076 11118 34078 11170
rect 34130 11118 34132 11170
rect 33628 10770 33684 10780
rect 34076 10612 34132 11118
rect 33516 10546 33572 10556
rect 33964 10556 34132 10612
rect 34188 11060 34244 11070
rect 33516 9940 33572 9950
rect 33516 9846 33572 9884
rect 33740 9268 33796 9278
rect 33404 9266 33796 9268
rect 33404 9214 33742 9266
rect 33794 9214 33796 9266
rect 33404 9212 33796 9214
rect 33292 8484 33348 8494
rect 33292 8370 33348 8428
rect 33292 8318 33294 8370
rect 33346 8318 33348 8370
rect 33292 8306 33348 8318
rect 33628 8372 33684 8382
rect 33628 7698 33684 8316
rect 33740 8260 33796 9212
rect 33740 8194 33796 8204
rect 33628 7646 33630 7698
rect 33682 7646 33684 7698
rect 33628 7634 33684 7646
rect 32956 6626 33012 6636
rect 32732 6468 32788 6478
rect 32620 6466 32788 6468
rect 32620 6414 32734 6466
rect 32786 6414 32788 6466
rect 32620 6412 32788 6414
rect 32396 5854 32398 5906
rect 32450 5854 32452 5906
rect 32060 5842 32116 5852
rect 32396 5842 32452 5854
rect 32508 5908 32564 5918
rect 32508 5814 32564 5852
rect 31612 5506 31668 5516
rect 31948 5122 32004 5134
rect 31948 5070 31950 5122
rect 32002 5070 32004 5122
rect 30940 4834 30996 4844
rect 31836 4900 31892 4910
rect 30828 4498 30884 4508
rect 31500 4564 31556 4574
rect 29820 4386 29876 4396
rect 29596 4174 29598 4226
rect 29650 4174 29652 4226
rect 29596 4162 29652 4174
rect 29708 4340 29764 4350
rect 29708 3780 29764 4284
rect 31500 4338 31556 4508
rect 31500 4286 31502 4338
rect 31554 4286 31556 4338
rect 31500 4274 31556 4286
rect 31836 4226 31892 4844
rect 31948 4452 32004 5070
rect 32620 4676 32676 6412
rect 32732 6402 32788 6412
rect 32956 6468 33012 6478
rect 33068 6468 33124 6478
rect 32956 6466 33068 6468
rect 32956 6414 32958 6466
rect 33010 6414 33068 6466
rect 32956 6412 33068 6414
rect 32956 6402 33012 6412
rect 31948 4386 32004 4396
rect 32396 4620 32676 4676
rect 32396 4450 32452 4620
rect 32844 4564 32900 4574
rect 32844 4470 32900 4508
rect 32396 4398 32398 4450
rect 32450 4398 32452 4450
rect 31836 4174 31838 4226
rect 31890 4174 31892 4226
rect 31836 4162 31892 4174
rect 32396 3892 32452 4398
rect 32172 3836 32452 3892
rect 29708 3666 29764 3724
rect 29708 3614 29710 3666
rect 29762 3614 29764 3666
rect 29708 3602 29764 3614
rect 30716 3780 30772 3790
rect 29260 3462 29316 3500
rect 27244 3378 27300 3388
rect 30156 3444 30212 3454
rect 14476 3266 14532 3276
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 30156 800 30212 3388
rect 30380 3444 30436 3482
rect 30380 3378 30436 3388
rect 30716 3330 30772 3724
rect 31612 3668 31668 3678
rect 31612 3554 31668 3612
rect 31612 3502 31614 3554
rect 31666 3502 31668 3554
rect 31612 3490 31668 3502
rect 32172 3554 32228 3836
rect 33068 3780 33124 6412
rect 33180 6466 33236 6478
rect 33180 6414 33182 6466
rect 33234 6414 33236 6466
rect 33180 6132 33236 6414
rect 33740 6468 33796 6478
rect 33740 6374 33796 6412
rect 33180 6066 33236 6076
rect 33628 6018 33684 6030
rect 33628 5966 33630 6018
rect 33682 5966 33684 6018
rect 33628 5236 33684 5966
rect 33852 5908 33908 5918
rect 33852 5814 33908 5852
rect 33628 5170 33684 5180
rect 32284 3668 32340 3678
rect 32284 3574 32340 3612
rect 33068 3666 33124 3724
rect 33068 3614 33070 3666
rect 33122 3614 33124 3666
rect 33068 3602 33124 3614
rect 33516 5010 33572 5022
rect 33516 4958 33518 5010
rect 33570 4958 33572 5010
rect 32172 3502 32174 3554
rect 32226 3502 32228 3554
rect 32172 3490 32228 3502
rect 33516 3444 33572 4958
rect 33964 5012 34020 10556
rect 34076 10388 34132 10398
rect 34188 10388 34244 11004
rect 34300 10948 34356 12796
rect 34412 12786 34468 12796
rect 34636 12180 34692 13580
rect 34636 12114 34692 12124
rect 34412 11956 34468 11966
rect 34636 11956 34692 11966
rect 34412 11954 34692 11956
rect 34412 11902 34414 11954
rect 34466 11902 34638 11954
rect 34690 11902 34692 11954
rect 34412 11900 34692 11902
rect 34412 11890 34468 11900
rect 34636 11890 34692 11900
rect 34748 11396 34804 11406
rect 34300 10892 34580 10948
rect 34076 10386 34244 10388
rect 34076 10334 34078 10386
rect 34130 10334 34244 10386
rect 34076 10332 34244 10334
rect 34300 10724 34356 10734
rect 34076 9940 34132 10332
rect 34076 9874 34132 9884
rect 34076 9716 34132 9726
rect 34300 9716 34356 10668
rect 34412 10386 34468 10398
rect 34412 10334 34414 10386
rect 34466 10334 34468 10386
rect 34412 9828 34468 10334
rect 34412 9762 34468 9772
rect 34076 9714 34356 9716
rect 34076 9662 34078 9714
rect 34130 9662 34356 9714
rect 34076 9660 34356 9662
rect 34076 9650 34132 9660
rect 34076 8372 34132 8382
rect 34076 8278 34132 8316
rect 34300 8260 34356 8270
rect 34300 8166 34356 8204
rect 34188 6692 34244 6702
rect 34188 5234 34244 6636
rect 34524 5684 34580 10892
rect 34636 9940 34692 9950
rect 34636 9266 34692 9884
rect 34748 9826 34804 11340
rect 34748 9774 34750 9826
rect 34802 9774 34804 9826
rect 34748 9762 34804 9774
rect 34636 9214 34638 9266
rect 34690 9214 34692 9266
rect 34636 9202 34692 9214
rect 34860 9268 34916 14588
rect 35084 14532 35140 14702
rect 34972 13076 35028 13086
rect 35084 13076 35140 14476
rect 35308 14756 35364 14766
rect 35308 14418 35364 14700
rect 35420 14756 35476 14766
rect 35644 14756 35700 14766
rect 35420 14754 35700 14756
rect 35420 14702 35422 14754
rect 35474 14702 35646 14754
rect 35698 14702 35700 14754
rect 35420 14700 35700 14702
rect 35420 14690 35476 14700
rect 35308 14366 35310 14418
rect 35362 14366 35364 14418
rect 35308 14354 35364 14366
rect 35420 13860 35476 13870
rect 35420 13766 35476 13804
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 34972 13074 35140 13076
rect 34972 13022 34974 13074
rect 35026 13022 35140 13074
rect 34972 13020 35140 13022
rect 34972 13010 35028 13020
rect 35420 12404 35476 12414
rect 34972 12292 35028 12302
rect 34972 12198 35028 12236
rect 35420 12068 35476 12348
rect 35532 12292 35588 14700
rect 35644 14690 35700 14700
rect 35532 12226 35588 12236
rect 35644 12180 35700 12190
rect 35420 12012 35588 12068
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35308 11620 35364 11630
rect 35532 11620 35588 12012
rect 35308 11618 35588 11620
rect 35308 11566 35310 11618
rect 35362 11566 35588 11618
rect 35308 11564 35588 11566
rect 35308 11554 35364 11564
rect 34972 11172 35028 11182
rect 34972 11170 35140 11172
rect 34972 11118 34974 11170
rect 35026 11118 35140 11170
rect 34972 11116 35140 11118
rect 34972 11106 35028 11116
rect 35084 10610 35140 11116
rect 35420 10724 35476 11564
rect 35644 11282 35700 12124
rect 35644 11230 35646 11282
rect 35698 11230 35700 11282
rect 35644 11218 35700 11230
rect 35420 10658 35476 10668
rect 35084 10558 35086 10610
rect 35138 10558 35140 10610
rect 35084 10546 35140 10558
rect 35308 10612 35364 10622
rect 35308 10518 35364 10556
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35084 9940 35140 9950
rect 35084 9826 35140 9884
rect 35084 9774 35086 9826
rect 35138 9774 35140 9826
rect 35084 9762 35140 9774
rect 35308 9828 35364 9838
rect 35308 9734 35364 9772
rect 34972 9716 35028 9726
rect 34972 9622 35028 9660
rect 35756 9604 35812 14924
rect 35980 14642 36036 15092
rect 36316 15090 36372 15102
rect 36316 15038 36318 15090
rect 36370 15038 36372 15090
rect 36316 14980 36372 15038
rect 36316 14914 36372 14924
rect 36428 14754 36484 15596
rect 36764 15540 36820 15550
rect 36764 15314 36820 15484
rect 36764 15262 36766 15314
rect 36818 15262 36820 15314
rect 36764 15250 36820 15262
rect 36428 14702 36430 14754
rect 36482 14702 36484 14754
rect 36428 14690 36484 14702
rect 36764 14756 36820 14766
rect 35980 14590 35982 14642
rect 36034 14590 36036 14642
rect 35980 14578 36036 14590
rect 36764 14642 36820 14700
rect 36764 14590 36766 14642
rect 36818 14590 36820 14642
rect 36764 14578 36820 14590
rect 36316 14420 36372 14430
rect 36316 14326 36372 14364
rect 36988 12516 37044 22988
rect 37100 23042 37492 23044
rect 37100 22990 37102 23042
rect 37154 22990 37492 23042
rect 37100 22988 37492 22990
rect 37548 23266 37604 23278
rect 38108 23268 38164 24108
rect 38220 24052 38276 28588
rect 38444 28196 38500 32396
rect 38668 32452 38724 32956
rect 38332 28140 38500 28196
rect 38556 32340 38612 32350
rect 38332 24164 38388 28140
rect 38556 27860 38612 32284
rect 38668 31220 38724 32396
rect 38780 31668 38836 33068
rect 38780 31602 38836 31612
rect 38892 32900 38948 32910
rect 38892 31666 38948 32844
rect 38892 31614 38894 31666
rect 38946 31614 38948 31666
rect 38892 31602 38948 31614
rect 38668 31164 38948 31220
rect 38892 30772 38948 31164
rect 39004 31108 39060 33180
rect 39116 32900 39172 32910
rect 39116 32786 39172 32844
rect 39116 32734 39118 32786
rect 39170 32734 39172 32786
rect 39116 32722 39172 32734
rect 39340 32788 39396 33740
rect 39564 33236 39620 34638
rect 39564 33170 39620 33180
rect 39676 32900 39732 35644
rect 39900 35606 39956 35644
rect 40124 35476 40180 35486
rect 39900 34692 39956 34702
rect 39900 34598 39956 34636
rect 39900 34244 39956 34254
rect 39676 32834 39732 32844
rect 39788 34188 39900 34244
rect 39228 32564 39284 32574
rect 39116 32338 39172 32350
rect 39116 32286 39118 32338
rect 39170 32286 39172 32338
rect 39116 31444 39172 32286
rect 39228 31778 39284 32508
rect 39228 31726 39230 31778
rect 39282 31726 39284 31778
rect 39228 31714 39284 31726
rect 39116 31378 39172 31388
rect 39116 31108 39172 31118
rect 39004 31052 39116 31108
rect 39116 31014 39172 31052
rect 39228 30884 39284 30894
rect 38892 30770 39060 30772
rect 38892 30718 38894 30770
rect 38946 30718 39060 30770
rect 38892 30716 39060 30718
rect 38892 30706 38948 30716
rect 38780 30660 38836 30670
rect 38780 28754 38836 30604
rect 38892 29988 38948 29998
rect 38892 29764 38948 29932
rect 38892 29650 38948 29708
rect 38892 29598 38894 29650
rect 38946 29598 38948 29650
rect 38892 29586 38948 29598
rect 38780 28702 38782 28754
rect 38834 28702 38836 28754
rect 38780 28420 38836 28702
rect 38780 28354 38836 28364
rect 38556 27794 38612 27804
rect 38668 27636 38724 27646
rect 38668 27188 38724 27580
rect 38668 27076 38724 27132
rect 38444 27020 38724 27076
rect 38892 27186 38948 27198
rect 38892 27134 38894 27186
rect 38946 27134 38948 27186
rect 38444 25618 38500 27020
rect 38780 26740 38836 26750
rect 38556 26516 38612 26526
rect 38556 26422 38612 26460
rect 38780 26516 38836 26684
rect 38444 25566 38446 25618
rect 38498 25566 38500 25618
rect 38444 25554 38500 25566
rect 38780 25618 38836 26460
rect 38780 25566 38782 25618
rect 38834 25566 38836 25618
rect 38780 25554 38836 25566
rect 38892 25956 38948 27134
rect 39004 26852 39060 30716
rect 39228 30098 39284 30828
rect 39228 30046 39230 30098
rect 39282 30046 39284 30098
rect 39228 30034 39284 30046
rect 39340 29988 39396 32732
rect 39788 32452 39844 34188
rect 39900 34150 39956 34188
rect 40012 34130 40068 34142
rect 40012 34078 40014 34130
rect 40066 34078 40068 34130
rect 40012 33796 40068 34078
rect 40012 33730 40068 33740
rect 40124 33572 40180 35420
rect 40236 34018 40292 37660
rect 40572 37156 40628 37166
rect 40572 37062 40628 37100
rect 40460 36258 40516 36270
rect 40460 36206 40462 36258
rect 40514 36206 40516 36258
rect 40460 35476 40516 36206
rect 40460 35382 40516 35420
rect 40684 35810 40740 37772
rect 40796 37762 40852 37772
rect 41244 37828 41300 37838
rect 41244 37826 41412 37828
rect 41244 37774 41246 37826
rect 41298 37774 41412 37826
rect 41244 37772 41412 37774
rect 41244 37762 41300 37772
rect 40684 35758 40686 35810
rect 40738 35758 40740 35810
rect 40236 33966 40238 34018
rect 40290 33966 40292 34018
rect 40236 33954 40292 33966
rect 40460 34690 40516 34702
rect 40460 34638 40462 34690
rect 40514 34638 40516 34690
rect 40460 33796 40516 34638
rect 40460 33730 40516 33740
rect 40012 33516 40180 33572
rect 40012 33234 40068 33516
rect 40012 33182 40014 33234
rect 40066 33182 40068 33234
rect 39900 33124 39956 33134
rect 39900 32562 39956 33068
rect 39900 32510 39902 32562
rect 39954 32510 39956 32562
rect 39900 32498 39956 32510
rect 39676 32396 39844 32452
rect 40012 32452 40068 33182
rect 40236 33460 40292 33470
rect 40124 33124 40180 33134
rect 40124 32562 40180 33068
rect 40236 33122 40292 33404
rect 40236 33070 40238 33122
rect 40290 33070 40292 33122
rect 40236 32788 40292 33070
rect 40236 32722 40292 32732
rect 40124 32510 40126 32562
rect 40178 32510 40180 32562
rect 40124 32498 40180 32510
rect 39452 31444 39508 31454
rect 39452 30210 39508 31388
rect 39452 30158 39454 30210
rect 39506 30158 39508 30210
rect 39452 30146 39508 30158
rect 39340 29932 39620 29988
rect 39452 28530 39508 28542
rect 39452 28478 39454 28530
rect 39506 28478 39508 28530
rect 39116 27748 39172 27758
rect 39452 27748 39508 28478
rect 39564 28196 39620 29932
rect 39676 28532 39732 32396
rect 40012 32386 40068 32396
rect 40684 32340 40740 35758
rect 41132 36482 41188 36494
rect 41132 36430 41134 36482
rect 41186 36430 41188 36482
rect 40796 35700 40852 35710
rect 40796 35586 40852 35644
rect 41132 35700 41188 36430
rect 41356 36484 41412 37772
rect 41468 37492 41524 37502
rect 41468 37398 41524 37436
rect 41356 36390 41412 36428
rect 41580 35812 41636 39340
rect 42028 39060 42084 39070
rect 42028 38966 42084 39004
rect 42140 37826 42196 37838
rect 42140 37774 42142 37826
rect 42194 37774 42196 37826
rect 42140 36932 42196 37774
rect 42140 36866 42196 36876
rect 41692 36596 41748 36606
rect 41692 36502 41748 36540
rect 41132 35634 41188 35644
rect 41356 35756 41636 35812
rect 41804 36484 41860 36494
rect 41804 35812 41860 36428
rect 42252 36260 42308 36270
rect 42252 36166 42308 36204
rect 42476 36036 42532 40572
rect 42588 40562 42644 40572
rect 43036 40514 43092 40908
rect 43148 40962 43204 40974
rect 43148 40910 43150 40962
rect 43202 40910 43204 40962
rect 43148 40740 43204 40910
rect 43148 40674 43204 40684
rect 43708 40962 43764 40974
rect 43708 40910 43710 40962
rect 43762 40910 43764 40962
rect 43708 40852 43764 40910
rect 43036 40462 43038 40514
rect 43090 40462 43092 40514
rect 42812 39844 42868 39854
rect 43036 39844 43092 40462
rect 43708 40404 43764 40796
rect 43708 40338 43764 40348
rect 42812 39842 43092 39844
rect 42812 39790 42814 39842
rect 42866 39790 43092 39842
rect 42812 39788 43092 39790
rect 43820 40292 43876 40302
rect 44156 40292 44212 41020
rect 44380 41010 44436 41020
rect 44604 41076 44660 41086
rect 44492 40962 44548 40974
rect 44492 40910 44494 40962
rect 44546 40910 44548 40962
rect 44268 40404 44324 40414
rect 44268 40310 44324 40348
rect 43820 40290 44212 40292
rect 43820 40238 43822 40290
rect 43874 40238 44212 40290
rect 43820 40236 44212 40238
rect 42588 39732 42644 39742
rect 42588 39058 42644 39676
rect 42588 39006 42590 39058
rect 42642 39006 42644 39058
rect 42588 38994 42644 39006
rect 42812 39060 42868 39788
rect 43148 39730 43204 39742
rect 43148 39678 43150 39730
rect 43202 39678 43204 39730
rect 42812 38994 42868 39004
rect 42924 39620 42980 39630
rect 42924 39058 42980 39564
rect 43148 39620 43204 39678
rect 43820 39730 43876 40236
rect 43820 39678 43822 39730
rect 43874 39678 43876 39730
rect 43820 39666 43876 39678
rect 43148 39554 43204 39564
rect 44268 39620 44324 39630
rect 44492 39620 44548 40910
rect 44604 40290 44660 41020
rect 45052 40404 45108 43262
rect 45052 40338 45108 40348
rect 44604 40238 44606 40290
rect 44658 40238 44660 40290
rect 44604 40226 44660 40238
rect 44268 39618 44548 39620
rect 44268 39566 44270 39618
rect 44322 39566 44548 39618
rect 44268 39564 44548 39566
rect 42924 39006 42926 39058
rect 42978 39006 42980 39058
rect 42924 38724 42980 39006
rect 44268 38948 44324 39564
rect 44716 39508 44772 39518
rect 44716 39414 44772 39452
rect 44268 38882 44324 38892
rect 44492 38836 44548 38846
rect 42924 38658 42980 38668
rect 43708 38724 43764 38734
rect 43596 38052 43652 38062
rect 43484 38050 43652 38052
rect 43484 37998 43598 38050
rect 43650 37998 43652 38050
rect 43484 37996 43652 37998
rect 42588 37266 42644 37278
rect 42588 37214 42590 37266
rect 42642 37214 42644 37266
rect 42588 36932 42644 37214
rect 42700 37156 42756 37166
rect 43372 37156 43428 37166
rect 42756 37100 42980 37156
rect 42700 37062 42756 37100
rect 42588 36372 42644 36876
rect 42924 36706 42980 37100
rect 43372 37062 43428 37100
rect 43484 36820 43540 37996
rect 43596 37986 43652 37996
rect 42924 36654 42926 36706
rect 42978 36654 42980 36706
rect 42924 36642 42980 36654
rect 43260 36764 43540 36820
rect 43260 36706 43316 36764
rect 43260 36654 43262 36706
rect 43314 36654 43316 36706
rect 43260 36642 43316 36654
rect 42700 36372 42756 36382
rect 42588 36370 42756 36372
rect 42588 36318 42702 36370
rect 42754 36318 42756 36370
rect 42588 36316 42756 36318
rect 42476 35970 42532 35980
rect 42700 35924 42756 36316
rect 42700 35858 42756 35868
rect 40796 35534 40798 35586
rect 40850 35534 40852 35586
rect 40796 35522 40852 35534
rect 40796 35028 40852 35038
rect 40796 34934 40852 34972
rect 40796 34244 40852 34254
rect 40796 34150 40852 34188
rect 41244 34244 41300 34254
rect 41244 33346 41300 34188
rect 41244 33294 41246 33346
rect 41298 33294 41300 33346
rect 41244 33282 41300 33294
rect 40908 33236 40964 33246
rect 40908 33142 40964 33180
rect 41020 33124 41076 33134
rect 41020 33030 41076 33068
rect 40684 32274 40740 32284
rect 40796 32450 40852 32462
rect 40796 32398 40798 32450
rect 40850 32398 40852 32450
rect 40012 31892 40068 31902
rect 40012 31798 40068 31836
rect 40236 31892 40292 31902
rect 39788 31444 39844 31454
rect 39788 31106 39844 31388
rect 39788 31054 39790 31106
rect 39842 31054 39844 31106
rect 39788 31042 39844 31054
rect 40012 31106 40068 31118
rect 40012 31054 40014 31106
rect 40066 31054 40068 31106
rect 39900 30882 39956 30894
rect 39900 30830 39902 30882
rect 39954 30830 39956 30882
rect 39788 29428 39844 29438
rect 39900 29428 39956 30830
rect 40012 30884 40068 31054
rect 40012 30818 40068 30828
rect 39788 29426 39956 29428
rect 39788 29374 39790 29426
rect 39842 29374 39956 29426
rect 39788 29372 39956 29374
rect 40012 30100 40068 30110
rect 40012 29428 40068 30044
rect 40012 29426 40180 29428
rect 40012 29374 40014 29426
rect 40066 29374 40180 29426
rect 40012 29372 40180 29374
rect 39788 29362 39844 29372
rect 40012 29362 40068 29372
rect 40012 28868 40068 28878
rect 40012 28774 40068 28812
rect 40124 28644 40180 29372
rect 40236 29426 40292 31836
rect 40572 31332 40628 31342
rect 40572 31218 40628 31276
rect 40572 31166 40574 31218
rect 40626 31166 40628 31218
rect 40572 31154 40628 31166
rect 40796 30884 40852 32398
rect 40796 30818 40852 30828
rect 40236 29374 40238 29426
rect 40290 29374 40292 29426
rect 40236 29362 40292 29374
rect 40348 30324 40404 30334
rect 40348 28754 40404 30268
rect 40572 30100 40628 30110
rect 40572 30006 40628 30044
rect 40460 29986 40516 29998
rect 40460 29934 40462 29986
rect 40514 29934 40516 29986
rect 40460 29428 40516 29934
rect 41244 29986 41300 29998
rect 41244 29934 41246 29986
rect 41298 29934 41300 29986
rect 40460 29334 40516 29372
rect 40684 29426 40740 29438
rect 40684 29374 40686 29426
rect 40738 29374 40740 29426
rect 40572 29314 40628 29326
rect 40572 29262 40574 29314
rect 40626 29262 40628 29314
rect 40572 29092 40628 29262
rect 40572 29026 40628 29036
rect 40684 28868 40740 29374
rect 40684 28802 40740 28812
rect 40348 28702 40350 28754
rect 40402 28702 40404 28754
rect 40348 28690 40404 28702
rect 40796 28756 40852 28766
rect 40796 28662 40852 28700
rect 40124 28588 40292 28644
rect 40236 28532 40292 28588
rect 40908 28532 40964 28542
rect 40236 28476 40404 28532
rect 39676 28400 39732 28476
rect 39900 28418 39956 28430
rect 39900 28366 39902 28418
rect 39954 28366 39956 28418
rect 39900 28196 39956 28366
rect 39564 28140 39732 28196
rect 39116 27746 39508 27748
rect 39116 27694 39118 27746
rect 39170 27694 39508 27746
rect 39116 27692 39508 27694
rect 39564 27858 39620 27870
rect 39564 27806 39566 27858
rect 39618 27806 39620 27858
rect 39116 27300 39172 27692
rect 39116 27234 39172 27244
rect 39452 27300 39508 27310
rect 39228 27188 39284 27198
rect 39228 27074 39284 27132
rect 39228 27022 39230 27074
rect 39282 27022 39284 27074
rect 39228 27010 39284 27022
rect 39004 26786 39060 26796
rect 39340 26964 39396 26974
rect 39340 26740 39396 26908
rect 39452 26962 39508 27244
rect 39564 27076 39620 27806
rect 39564 27010 39620 27020
rect 39452 26910 39454 26962
rect 39506 26910 39508 26962
rect 39452 26898 39508 26910
rect 39676 26908 39732 28140
rect 39900 28130 39956 28140
rect 40236 28196 40292 28206
rect 40012 27746 40068 27758
rect 40012 27694 40014 27746
rect 40066 27694 40068 27746
rect 40012 27636 40068 27694
rect 40012 27570 40068 27580
rect 40236 27412 40292 28140
rect 39676 26852 39844 26908
rect 39340 26684 39620 26740
rect 39228 26402 39284 26414
rect 39228 26350 39230 26402
rect 39282 26350 39284 26402
rect 38780 24724 38836 24734
rect 38780 24630 38836 24668
rect 38332 24108 38724 24164
rect 38220 23986 38276 23996
rect 38332 23940 38388 23950
rect 38332 23846 38388 23884
rect 37548 23214 37550 23266
rect 37602 23214 37604 23266
rect 37100 22978 37156 22988
rect 37436 22484 37492 22494
rect 37548 22484 37604 23214
rect 37436 22482 37604 22484
rect 37436 22430 37438 22482
rect 37490 22430 37604 22482
rect 37436 22428 37604 22430
rect 37660 23212 38164 23268
rect 38220 23828 38276 23838
rect 37436 22418 37492 22428
rect 37324 22148 37380 22158
rect 37212 21812 37268 21822
rect 37100 21588 37156 21598
rect 37100 21494 37156 21532
rect 37100 18452 37156 18462
rect 37212 18452 37268 21756
rect 37324 18676 37380 22092
rect 37436 21586 37492 21598
rect 37436 21534 37438 21586
rect 37490 21534 37492 21586
rect 37436 19906 37492 21534
rect 37548 20804 37604 20814
rect 37548 20710 37604 20748
rect 37548 20132 37604 20142
rect 37548 20038 37604 20076
rect 37436 19854 37438 19906
rect 37490 19854 37492 19906
rect 37436 19842 37492 19854
rect 37324 18610 37380 18620
rect 37436 19010 37492 19022
rect 37436 18958 37438 19010
rect 37490 18958 37492 19010
rect 37436 18674 37492 18958
rect 37436 18622 37438 18674
rect 37490 18622 37492 18674
rect 37436 18564 37492 18622
rect 37436 18498 37492 18508
rect 37100 18450 37268 18452
rect 37100 18398 37102 18450
rect 37154 18398 37268 18450
rect 37100 18396 37268 18398
rect 37100 18386 37156 18396
rect 37660 18116 37716 23212
rect 38220 23154 38276 23772
rect 38220 23102 38222 23154
rect 38274 23102 38276 23154
rect 38220 23090 38276 23102
rect 38444 23716 38500 23726
rect 38668 23716 38724 24108
rect 37996 23044 38052 23054
rect 37884 22148 37940 22158
rect 37996 22148 38052 22988
rect 38444 23042 38500 23660
rect 38444 22990 38446 23042
rect 38498 22990 38500 23042
rect 38444 22978 38500 22990
rect 38556 23660 38724 23716
rect 38332 22148 38388 22158
rect 37772 22146 38388 22148
rect 37772 22094 37886 22146
rect 37938 22094 38334 22146
rect 38386 22094 38388 22146
rect 37772 22092 38388 22094
rect 37772 21810 37828 22092
rect 37884 22082 37940 22092
rect 38332 22082 38388 22092
rect 37772 21758 37774 21810
rect 37826 21758 37828 21810
rect 37772 21746 37828 21758
rect 37884 21924 37940 21934
rect 37884 20802 37940 21868
rect 38220 21812 38276 21822
rect 38220 21718 38276 21756
rect 37884 20750 37886 20802
rect 37938 20750 37940 20802
rect 37884 20738 37940 20750
rect 38108 20916 38164 20926
rect 38108 20802 38164 20860
rect 38108 20750 38110 20802
rect 38162 20750 38164 20802
rect 38108 20738 38164 20750
rect 37996 20578 38052 20590
rect 37996 20526 37998 20578
rect 38050 20526 38052 20578
rect 37996 20244 38052 20526
rect 38556 20580 38612 23660
rect 38780 23044 38836 23054
rect 38780 22950 38836 22988
rect 38780 22146 38836 22158
rect 38780 22094 38782 22146
rect 38834 22094 38836 22146
rect 38780 21812 38836 22094
rect 38780 21746 38836 21756
rect 38892 21588 38948 25900
rect 39004 26292 39060 26302
rect 39004 24050 39060 26236
rect 39228 25732 39284 26350
rect 39564 26290 39620 26684
rect 39564 26238 39566 26290
rect 39618 26238 39620 26290
rect 39284 25676 39396 25732
rect 39228 25666 39284 25676
rect 39228 25284 39284 25294
rect 39228 25190 39284 25228
rect 39004 23998 39006 24050
rect 39058 23998 39060 24050
rect 39004 23828 39060 23998
rect 39004 23762 39060 23772
rect 39340 22708 39396 25676
rect 39452 24498 39508 24510
rect 39452 24446 39454 24498
rect 39506 24446 39508 24498
rect 39452 24164 39508 24446
rect 39452 24098 39508 24108
rect 39564 24050 39620 26238
rect 39564 23998 39566 24050
rect 39618 23998 39620 24050
rect 39564 23986 39620 23998
rect 39676 25844 39732 25854
rect 39676 25618 39732 25788
rect 39676 25566 39678 25618
rect 39730 25566 39732 25618
rect 39676 23380 39732 25566
rect 39564 23324 39732 23380
rect 39340 22652 39508 22708
rect 39340 22484 39396 22494
rect 39340 22390 39396 22428
rect 39228 22036 39284 22046
rect 38780 21532 38948 21588
rect 39116 21924 39172 21934
rect 38556 20486 38612 20524
rect 38668 20916 38724 20926
rect 37996 20178 38052 20188
rect 38668 19460 38724 20860
rect 38780 19572 38836 21532
rect 38892 21364 38948 21374
rect 38892 21270 38948 21308
rect 39116 21026 39172 21868
rect 39228 21588 39284 21980
rect 39228 21522 39284 21532
rect 39116 20974 39118 21026
rect 39170 20974 39172 21026
rect 39004 20578 39060 20590
rect 39004 20526 39006 20578
rect 39058 20526 39060 20578
rect 39004 20356 39060 20526
rect 39004 20290 39060 20300
rect 39116 20130 39172 20974
rect 39116 20078 39118 20130
rect 39170 20078 39172 20130
rect 38780 19516 38948 19572
rect 38668 19404 38836 19460
rect 38444 19348 38500 19358
rect 38444 19346 38724 19348
rect 38444 19294 38446 19346
rect 38498 19294 38724 19346
rect 38444 19292 38724 19294
rect 38444 19282 38500 19292
rect 37884 19236 37940 19246
rect 37884 19142 37940 19180
rect 38668 19234 38724 19292
rect 38668 19182 38670 19234
rect 38722 19182 38724 19234
rect 38668 19170 38724 19182
rect 38780 19346 38836 19404
rect 38780 19294 38782 19346
rect 38834 19294 38836 19346
rect 38780 18564 38836 19294
rect 38668 18562 38836 18564
rect 38668 18510 38782 18562
rect 38834 18510 38836 18562
rect 38668 18508 38836 18510
rect 38556 18452 38612 18462
rect 37996 18450 38612 18452
rect 37996 18398 38558 18450
rect 38610 18398 38612 18450
rect 37996 18396 38612 18398
rect 37884 18340 37940 18350
rect 37548 18060 37716 18116
rect 37772 18338 37940 18340
rect 37772 18286 37886 18338
rect 37938 18286 37940 18338
rect 37772 18284 37940 18286
rect 37436 17892 37492 17902
rect 37436 16882 37492 17836
rect 37436 16830 37438 16882
rect 37490 16830 37492 16882
rect 37436 16818 37492 16830
rect 37548 16772 37604 18060
rect 37660 17892 37716 17902
rect 37660 17798 37716 17836
rect 37772 17556 37828 18284
rect 37884 18274 37940 18284
rect 37996 17890 38052 18396
rect 38556 18386 38612 18396
rect 38668 18116 38724 18508
rect 38780 18498 38836 18508
rect 37996 17838 37998 17890
rect 38050 17838 38052 17890
rect 37996 17826 38052 17838
rect 38556 18060 38724 18116
rect 38892 18116 38948 19516
rect 39116 19458 39172 20078
rect 39116 19406 39118 19458
rect 39170 19406 39172 19458
rect 39116 19394 39172 19406
rect 39228 21362 39284 21374
rect 39228 21310 39230 21362
rect 39282 21310 39284 21362
rect 39228 21252 39284 21310
rect 39004 18564 39060 18574
rect 39004 18470 39060 18508
rect 39116 18450 39172 18462
rect 39116 18398 39118 18450
rect 39170 18398 39172 18450
rect 38892 18060 39060 18116
rect 38556 17892 38612 18060
rect 38556 17836 38724 17892
rect 37772 17490 37828 17500
rect 38332 17780 38388 17790
rect 37884 17444 37940 17454
rect 37884 16882 37940 17388
rect 38332 16994 38388 17724
rect 38668 17668 38724 17836
rect 38892 17780 38948 17790
rect 38892 17686 38948 17724
rect 38780 17668 38836 17678
rect 38668 17666 38836 17668
rect 38668 17614 38782 17666
rect 38834 17614 38836 17666
rect 38668 17612 38836 17614
rect 38780 17108 38836 17612
rect 39004 17444 39060 18060
rect 39116 17780 39172 18398
rect 39116 17714 39172 17724
rect 39004 17388 39172 17444
rect 39004 17220 39060 17230
rect 38892 17108 38948 17118
rect 38780 17106 38948 17108
rect 38780 17054 38894 17106
rect 38946 17054 38948 17106
rect 38780 17052 38948 17054
rect 38892 17042 38948 17052
rect 38332 16942 38334 16994
rect 38386 16942 38388 16994
rect 38332 16930 38388 16942
rect 37884 16830 37886 16882
rect 37938 16830 37940 16882
rect 37884 16818 37940 16830
rect 37548 16706 37604 16716
rect 39004 16324 39060 17164
rect 39116 16436 39172 17388
rect 39116 16370 39172 16380
rect 38892 16268 39060 16324
rect 37436 16212 37492 16222
rect 37436 16118 37492 16156
rect 37884 16212 37940 16222
rect 37884 16118 37940 16156
rect 38444 16212 38500 16222
rect 38444 16118 38500 16156
rect 38108 15540 38164 15550
rect 37436 15428 37492 15438
rect 37436 15334 37492 15372
rect 37996 15428 38052 15438
rect 37996 15334 38052 15372
rect 37212 15316 37268 15326
rect 37212 15222 37268 15260
rect 37324 15202 37380 15214
rect 37324 15150 37326 15202
rect 37378 15150 37380 15202
rect 37324 15148 37380 15150
rect 37324 15092 38052 15148
rect 37772 14980 37828 14990
rect 37772 13858 37828 14924
rect 37772 13806 37774 13858
rect 37826 13806 37828 13858
rect 37772 13794 37828 13806
rect 37996 13858 38052 15092
rect 38108 14418 38164 15484
rect 38892 15538 38948 16268
rect 39116 16212 39172 16222
rect 39004 16100 39060 16110
rect 39004 16006 39060 16044
rect 39116 15986 39172 16156
rect 39116 15934 39118 15986
rect 39170 15934 39172 15986
rect 39116 15922 39172 15934
rect 39228 15652 39284 21196
rect 39452 21028 39508 22652
rect 39564 21924 39620 23324
rect 39676 23156 39732 23166
rect 39676 23062 39732 23100
rect 39788 22932 39844 26852
rect 40124 26292 40180 26302
rect 40124 26198 40180 26236
rect 39900 26180 39956 26190
rect 39900 26086 39956 26124
rect 40236 25844 40292 27356
rect 40348 26404 40404 28476
rect 40460 27746 40516 27758
rect 40460 27694 40462 27746
rect 40514 27694 40516 27746
rect 40460 26852 40516 27694
rect 40572 27076 40628 27086
rect 40572 26982 40628 27020
rect 40908 27074 40964 28476
rect 41132 28308 41188 28318
rect 40908 27022 40910 27074
rect 40962 27022 40964 27074
rect 40908 26964 40964 27022
rect 40908 26898 40964 26908
rect 41020 27636 41076 27646
rect 40460 26786 40516 26796
rect 40796 26852 40852 26862
rect 40796 26758 40852 26796
rect 40348 26338 40404 26348
rect 40460 26516 40516 26526
rect 40236 25778 40292 25788
rect 40124 25732 40180 25742
rect 40012 24948 40068 24958
rect 40124 24948 40180 25676
rect 40012 24946 40180 24948
rect 40012 24894 40014 24946
rect 40066 24894 40180 24946
rect 40012 24892 40180 24894
rect 40460 24946 40516 26460
rect 41020 26292 41076 27580
rect 40684 26068 40740 26078
rect 40684 25508 40740 26012
rect 41020 25618 41076 26236
rect 41020 25566 41022 25618
rect 41074 25566 41076 25618
rect 41020 25554 41076 25566
rect 40460 24894 40462 24946
rect 40514 24894 40516 24946
rect 40012 24882 40068 24892
rect 39900 24500 39956 24510
rect 39900 24050 39956 24444
rect 39900 23998 39902 24050
rect 39954 23998 39956 24050
rect 39900 23986 39956 23998
rect 40012 24498 40068 24510
rect 40012 24446 40014 24498
rect 40066 24446 40068 24498
rect 40012 23828 40068 24446
rect 40460 24498 40516 24894
rect 40460 24446 40462 24498
rect 40514 24446 40516 24498
rect 40460 24434 40516 24446
rect 40572 25506 40740 25508
rect 40572 25454 40686 25506
rect 40738 25454 40740 25506
rect 40572 25452 40740 25454
rect 40460 24052 40516 24062
rect 40572 24052 40628 25452
rect 40684 25442 40740 25452
rect 41132 25172 41188 28252
rect 41244 27748 41300 29934
rect 41244 27682 41300 27692
rect 41356 27636 41412 35756
rect 41804 35698 41860 35756
rect 43484 35812 43540 35822
rect 43484 35718 43540 35756
rect 41804 35646 41806 35698
rect 41858 35646 41860 35698
rect 41804 35634 41860 35646
rect 42028 35700 42084 35710
rect 42028 35606 42084 35644
rect 41580 35586 41636 35598
rect 41580 35534 41582 35586
rect 41634 35534 41636 35586
rect 41580 35140 41636 35534
rect 43036 35586 43092 35598
rect 43036 35534 43038 35586
rect 43090 35534 43092 35586
rect 42476 35476 42532 35486
rect 41692 35140 41748 35150
rect 41580 35084 41692 35140
rect 41692 35008 41748 35084
rect 42028 35026 42084 35038
rect 42028 34974 42030 35026
rect 42082 34974 42084 35026
rect 42028 34916 42084 34974
rect 42028 34850 42084 34860
rect 41916 34690 41972 34702
rect 41916 34638 41918 34690
rect 41970 34638 41972 34690
rect 41468 34132 41524 34142
rect 41468 34038 41524 34076
rect 41916 34020 41972 34638
rect 41916 33954 41972 33964
rect 42028 34692 42084 34702
rect 41468 33684 41524 33694
rect 41468 33124 41524 33628
rect 41692 33572 41748 33582
rect 41580 33124 41636 33134
rect 41468 33122 41636 33124
rect 41468 33070 41582 33122
rect 41634 33070 41636 33122
rect 41468 33068 41636 33070
rect 41468 28308 41524 33068
rect 41580 33058 41636 33068
rect 41692 31778 41748 33516
rect 42028 33124 42084 34636
rect 42364 34020 42420 34030
rect 42364 33926 42420 33964
rect 42476 33570 42532 35420
rect 43036 35476 43092 35534
rect 43036 35410 43092 35420
rect 43708 35364 43764 38668
rect 44156 38052 44212 38062
rect 44156 37958 44212 37996
rect 44044 37826 44100 37838
rect 44044 37774 44046 37826
rect 44098 37774 44100 37826
rect 43932 36708 43988 36718
rect 44044 36708 44100 37774
rect 44268 37826 44324 37838
rect 44268 37774 44270 37826
rect 44322 37774 44324 37826
rect 44156 37156 44212 37166
rect 44268 37156 44324 37774
rect 44212 37100 44324 37156
rect 44380 37266 44436 37278
rect 44380 37214 44382 37266
rect 44434 37214 44436 37266
rect 44156 37062 44212 37100
rect 43932 36706 44100 36708
rect 43932 36654 43934 36706
rect 43986 36654 44100 36706
rect 43932 36652 44100 36654
rect 43932 36642 43988 36652
rect 43820 36596 43876 36606
rect 43820 36502 43876 36540
rect 44380 36596 44436 37214
rect 44380 36530 44436 36540
rect 44156 36260 44212 36270
rect 43708 35298 43764 35308
rect 44044 35586 44100 35598
rect 44044 35534 44046 35586
rect 44098 35534 44100 35586
rect 43932 35140 43988 35150
rect 42588 34916 42644 34926
rect 42588 34822 42644 34860
rect 43260 34916 43316 34926
rect 43596 34916 43652 34926
rect 43260 34914 43652 34916
rect 43260 34862 43262 34914
rect 43314 34862 43598 34914
rect 43650 34862 43652 34914
rect 43260 34860 43652 34862
rect 43260 34850 43316 34860
rect 43596 34850 43652 34860
rect 43932 34914 43988 35084
rect 43932 34862 43934 34914
rect 43986 34862 43988 34914
rect 42700 34804 42756 34814
rect 42700 34710 42756 34748
rect 42812 34690 42868 34702
rect 42812 34638 42814 34690
rect 42866 34638 42868 34690
rect 42588 34244 42644 34254
rect 42588 34150 42644 34188
rect 42812 34244 42868 34638
rect 42812 34178 42868 34188
rect 43820 34692 43876 34702
rect 43820 34020 43876 34636
rect 43932 34130 43988 34862
rect 44044 34692 44100 35534
rect 44044 34626 44100 34636
rect 43932 34078 43934 34130
rect 43986 34078 43988 34130
rect 43932 34066 43988 34078
rect 43820 33954 43876 33964
rect 42476 33518 42478 33570
rect 42530 33518 42532 33570
rect 42476 33458 42532 33518
rect 42476 33406 42478 33458
rect 42530 33406 42532 33458
rect 42476 33394 42532 33406
rect 43372 33570 43428 33582
rect 43372 33518 43374 33570
rect 43426 33518 43428 33570
rect 43372 33458 43428 33518
rect 43372 33406 43374 33458
rect 43426 33406 43428 33458
rect 43372 33394 43428 33406
rect 42028 33122 42308 33124
rect 42028 33070 42030 33122
rect 42082 33070 42308 33122
rect 42028 33068 42308 33070
rect 42028 33058 42084 33068
rect 42252 33012 42308 33068
rect 43036 33122 43092 33134
rect 43036 33070 43038 33122
rect 43090 33070 43092 33122
rect 42252 32956 42420 33012
rect 42140 32900 42196 32910
rect 41916 32564 41972 32574
rect 41916 31892 41972 32508
rect 41916 31826 41972 31836
rect 42028 32338 42084 32350
rect 42028 32286 42030 32338
rect 42082 32286 42084 32338
rect 41692 31726 41694 31778
rect 41746 31726 41748 31778
rect 41692 31668 41748 31726
rect 41692 31602 41748 31612
rect 41804 30994 41860 31006
rect 41804 30942 41806 30994
rect 41858 30942 41860 30994
rect 41804 30212 41860 30942
rect 42028 30434 42084 32286
rect 42140 31556 42196 32844
rect 42252 31780 42308 31790
rect 42252 31686 42308 31724
rect 42140 31500 42308 31556
rect 42140 30884 42196 30894
rect 42140 30790 42196 30828
rect 42028 30382 42030 30434
rect 42082 30382 42084 30434
rect 42028 30370 42084 30382
rect 41804 30146 41860 30156
rect 42252 30210 42308 31500
rect 42252 30158 42254 30210
rect 42306 30158 42308 30210
rect 42252 30146 42308 30158
rect 42028 30100 42084 30110
rect 41692 29988 41748 29998
rect 41692 29894 41748 29932
rect 41692 29428 41748 29438
rect 41692 29334 41748 29372
rect 41916 29426 41972 29438
rect 41916 29374 41918 29426
rect 41970 29374 41972 29426
rect 41580 29204 41636 29214
rect 41580 28530 41636 29148
rect 41916 28868 41972 29374
rect 41916 28802 41972 28812
rect 41580 28478 41582 28530
rect 41634 28478 41636 28530
rect 41580 28466 41636 28478
rect 41916 28532 41972 28542
rect 41916 28438 41972 28476
rect 41692 28418 41748 28430
rect 41692 28366 41694 28418
rect 41746 28366 41748 28418
rect 41692 28308 41748 28366
rect 42028 28308 42084 30044
rect 42364 28644 42420 32956
rect 43036 32676 43092 33070
rect 43036 32610 43092 32620
rect 43820 33122 43876 33134
rect 43820 33070 43822 33122
rect 43874 33070 43876 33122
rect 43820 32788 43876 33070
rect 42924 32564 42980 32574
rect 42924 32470 42980 32508
rect 42700 32450 42756 32462
rect 42700 32398 42702 32450
rect 42754 32398 42756 32450
rect 42588 31780 42644 31790
rect 42588 31108 42644 31724
rect 42588 29988 42644 31052
rect 42700 31220 42756 32398
rect 43596 32450 43652 32462
rect 43596 32398 43598 32450
rect 43650 32398 43652 32450
rect 43596 31780 43652 32398
rect 43820 32340 43876 32732
rect 44044 32900 44100 32910
rect 44044 32786 44100 32844
rect 44044 32734 44046 32786
rect 44098 32734 44100 32786
rect 44044 32722 44100 32734
rect 43820 32274 43876 32284
rect 43596 31714 43652 31724
rect 43820 32004 43876 32014
rect 43820 31778 43876 31948
rect 43820 31726 43822 31778
rect 43874 31726 43876 31778
rect 43820 31714 43876 31726
rect 42700 31106 42756 31164
rect 42700 31054 42702 31106
rect 42754 31054 42756 31106
rect 42700 31042 42756 31054
rect 42812 31666 42868 31678
rect 42812 31614 42814 31666
rect 42866 31614 42868 31666
rect 42812 30884 42868 31614
rect 42812 30818 42868 30828
rect 42924 31554 42980 31566
rect 42924 31502 42926 31554
rect 42978 31502 42980 31554
rect 42924 30212 42980 31502
rect 43148 31554 43204 31566
rect 43148 31502 43150 31554
rect 43202 31502 43204 31554
rect 43148 30994 43204 31502
rect 43820 31220 43876 31230
rect 43820 31126 43876 31164
rect 43148 30942 43150 30994
rect 43202 30942 43204 30994
rect 43148 30930 43204 30942
rect 43596 30994 43652 31006
rect 43596 30942 43598 30994
rect 43650 30942 43652 30994
rect 43596 30434 43652 30942
rect 43708 30884 43764 30894
rect 43708 30790 43764 30828
rect 43596 30382 43598 30434
rect 43650 30382 43652 30434
rect 43596 30370 43652 30382
rect 44044 30770 44100 30782
rect 44044 30718 44046 30770
rect 44098 30718 44100 30770
rect 44044 30322 44100 30718
rect 44044 30270 44046 30322
rect 44098 30270 44100 30322
rect 44044 30258 44100 30270
rect 42924 30146 42980 30156
rect 43484 30100 43540 30110
rect 43484 30006 43540 30044
rect 43036 29988 43092 29998
rect 42588 29986 43092 29988
rect 42588 29934 42590 29986
rect 42642 29934 43038 29986
rect 43090 29934 43092 29986
rect 42588 29932 43092 29934
rect 42588 29922 42644 29932
rect 43036 29922 43092 29932
rect 44156 29764 44212 36204
rect 44380 36258 44436 36270
rect 44380 36206 44382 36258
rect 44434 36206 44436 36258
rect 44380 35924 44436 36206
rect 44380 35858 44436 35868
rect 44492 35922 44548 38780
rect 44940 38836 44996 38846
rect 44940 38742 44996 38780
rect 45164 38668 45220 45052
rect 45724 44994 45780 45388
rect 45724 44942 45726 44994
rect 45778 44942 45780 44994
rect 45276 44882 45332 44894
rect 45276 44830 45278 44882
rect 45330 44830 45332 44882
rect 45276 43652 45332 44830
rect 45724 44548 45780 44942
rect 45500 44492 45724 44548
rect 45500 43762 45556 44492
rect 45724 44482 45780 44492
rect 46620 45778 46676 45790
rect 46620 45726 46622 45778
rect 46674 45726 46676 45778
rect 46620 44994 46676 45726
rect 46732 45666 46788 45678
rect 46732 45614 46734 45666
rect 46786 45614 46788 45666
rect 46732 45108 46788 45614
rect 46732 45042 46788 45052
rect 47068 45108 47124 45118
rect 47068 45014 47124 45052
rect 46620 44942 46622 44994
rect 46674 44942 46676 44994
rect 45836 44436 45892 44446
rect 45836 44342 45892 44380
rect 46172 44436 46228 44446
rect 46172 44322 46228 44380
rect 46172 44270 46174 44322
rect 46226 44270 46228 44322
rect 46172 44258 46228 44270
rect 46620 44322 46676 44942
rect 47180 44660 47236 46508
rect 47180 44594 47236 44604
rect 46620 44270 46622 44322
rect 46674 44270 46676 44322
rect 46620 44258 46676 44270
rect 45500 43710 45502 43762
rect 45554 43710 45556 43762
rect 45500 43698 45556 43710
rect 45276 42980 45332 43596
rect 45836 43428 45892 43438
rect 45500 42980 45556 42990
rect 45276 42978 45556 42980
rect 45276 42926 45502 42978
rect 45554 42926 45556 42978
rect 45276 42924 45556 42926
rect 45500 42914 45556 42924
rect 45836 42978 45892 43372
rect 46060 43426 46116 43438
rect 46060 43374 46062 43426
rect 46114 43374 46116 43426
rect 46060 43316 46116 43374
rect 46060 43250 46116 43260
rect 46620 43426 46676 43438
rect 46620 43374 46622 43426
rect 46674 43374 46676 43426
rect 45836 42926 45838 42978
rect 45890 42926 45892 42978
rect 45836 42532 45892 42926
rect 46060 42756 46116 42766
rect 46620 42756 46676 43374
rect 46956 43428 47012 43438
rect 46956 43334 47012 43372
rect 47404 43426 47460 50540
rect 48524 50706 48580 50718
rect 48524 50654 48526 50706
rect 48578 50654 48580 50706
rect 48412 50484 48468 50494
rect 48412 49924 48468 50428
rect 48412 49858 48468 49868
rect 48188 49812 48244 49822
rect 48188 49718 48244 49756
rect 48524 49700 48580 50654
rect 48412 49588 48468 49598
rect 48524 49588 48580 49644
rect 48412 49586 48580 49588
rect 48412 49534 48414 49586
rect 48466 49534 48580 49586
rect 48412 49532 48580 49534
rect 48412 49252 48468 49532
rect 48412 49186 48468 49196
rect 48636 48804 48692 52780
rect 49084 53620 49140 53630
rect 49084 52836 49140 53564
rect 49196 53508 49252 53518
rect 49196 53414 49252 53452
rect 49868 53508 49924 53518
rect 49868 52946 49924 53452
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 50652 53060 50708 53070
rect 51324 53060 51380 53678
rect 51436 54514 51492 54526
rect 51436 54462 51438 54514
rect 51490 54462 51492 54514
rect 51436 53732 51492 54462
rect 51772 54516 51828 54526
rect 51772 54422 51828 54460
rect 51772 53732 51828 53742
rect 51436 53730 51828 53732
rect 51436 53678 51774 53730
rect 51826 53678 51828 53730
rect 51436 53676 51828 53678
rect 50652 53058 51380 53060
rect 50652 53006 50654 53058
rect 50706 53006 51380 53058
rect 50652 53004 51380 53006
rect 50652 52994 50708 53004
rect 49868 52894 49870 52946
rect 49922 52894 49924 52946
rect 49868 52882 49924 52894
rect 49084 52770 49140 52780
rect 50092 52836 50148 52846
rect 49980 50594 50036 50606
rect 49980 50542 49982 50594
rect 50034 50542 50036 50594
rect 48972 50482 49028 50494
rect 49980 50484 50036 50542
rect 48972 50430 48974 50482
rect 49026 50430 49028 50482
rect 48972 50428 49028 50430
rect 49532 50428 50036 50484
rect 48972 50372 49140 50428
rect 49084 49812 49140 50372
rect 49084 49746 49140 49756
rect 49420 50372 49588 50428
rect 50092 50372 50148 52780
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 51548 51266 51604 51278
rect 51548 51214 51550 51266
rect 51602 51214 51604 51266
rect 51548 50820 51604 51214
rect 51772 51156 51828 53676
rect 50652 50818 51604 50820
rect 50652 50766 51550 50818
rect 51602 50766 51604 50818
rect 50652 50764 51604 50766
rect 50652 50706 50708 50764
rect 51548 50754 51604 50764
rect 51660 51100 51828 51156
rect 51884 51378 51940 51390
rect 51884 51326 51886 51378
rect 51938 51326 51940 51378
rect 50652 50654 50654 50706
rect 50706 50654 50708 50706
rect 50652 50642 50708 50654
rect 51660 50596 51716 51100
rect 48748 49588 48804 49598
rect 48748 49586 49028 49588
rect 48748 49534 48750 49586
rect 48802 49534 49028 49586
rect 48748 49532 49028 49534
rect 48748 49522 48804 49532
rect 48972 49026 49028 49532
rect 48972 48974 48974 49026
rect 49026 48974 49028 49026
rect 48972 48962 49028 48974
rect 49420 49026 49476 50372
rect 49644 50316 50148 50372
rect 51212 50540 51716 50596
rect 51212 50370 51268 50540
rect 51212 50318 51214 50370
rect 51266 50318 51268 50370
rect 49532 49812 49588 49822
rect 49532 49718 49588 49756
rect 49644 49476 49700 50316
rect 51212 50306 51268 50318
rect 51772 50484 51828 50494
rect 51884 50484 51940 51326
rect 51772 50482 51940 50484
rect 51772 50430 51774 50482
rect 51826 50430 51940 50482
rect 51772 50428 51940 50430
rect 51772 50372 51828 50428
rect 51772 50306 51828 50316
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 51996 50148 52052 55244
rect 52108 54740 52164 55412
rect 53452 55410 53732 55412
rect 53452 55358 53678 55410
rect 53730 55358 53732 55410
rect 53452 55356 53732 55358
rect 52220 54740 52276 54750
rect 53452 54740 53508 55356
rect 53676 55346 53732 55356
rect 53788 55412 54068 55468
rect 53788 55186 53844 55412
rect 53788 55134 53790 55186
rect 53842 55134 53844 55186
rect 53788 55122 53844 55134
rect 54012 55186 54068 55198
rect 54012 55134 54014 55186
rect 54066 55134 54068 55186
rect 54012 55076 54068 55134
rect 54012 55010 54068 55020
rect 54460 55076 54516 55086
rect 54460 54982 54516 55020
rect 52108 54738 52276 54740
rect 52108 54686 52222 54738
rect 52274 54686 52276 54738
rect 52108 54684 52276 54686
rect 52220 54674 52276 54684
rect 53340 54738 53508 54740
rect 53340 54686 53454 54738
rect 53506 54686 53508 54738
rect 53340 54684 53508 54686
rect 52444 54628 52500 54638
rect 52444 54534 52500 54572
rect 53228 54628 53284 54638
rect 52556 54514 52612 54526
rect 52556 54462 52558 54514
rect 52610 54462 52612 54514
rect 50556 50138 50820 50148
rect 51772 50092 52052 50148
rect 52108 53956 52164 53966
rect 50204 49812 50260 49822
rect 49756 49700 49812 49710
rect 49756 49606 49812 49644
rect 50092 49588 50148 49598
rect 49532 49420 49700 49476
rect 49868 49586 50148 49588
rect 49868 49534 50094 49586
rect 50146 49534 50148 49586
rect 49868 49532 50148 49534
rect 49532 49138 49588 49420
rect 49532 49086 49534 49138
rect 49586 49086 49588 49138
rect 49532 49074 49588 49086
rect 49420 48974 49422 49026
rect 49474 48974 49476 49026
rect 48188 47346 48244 47358
rect 48188 47294 48190 47346
rect 48242 47294 48244 47346
rect 47852 47124 47908 47134
rect 47852 46674 47908 47068
rect 47852 46622 47854 46674
rect 47906 46622 47908 46674
rect 47852 46610 47908 46622
rect 47964 46564 48020 46574
rect 48188 46564 48244 47294
rect 48300 47234 48356 47246
rect 48300 47182 48302 47234
rect 48354 47182 48356 47234
rect 48300 47124 48356 47182
rect 48300 47058 48356 47068
rect 48524 47234 48580 47246
rect 48524 47182 48526 47234
rect 48578 47182 48580 47234
rect 48524 46900 48580 47182
rect 48636 47012 48692 48748
rect 49420 48468 49476 48974
rect 49644 49028 49700 49038
rect 49868 49028 49924 49532
rect 50092 49522 50148 49532
rect 50204 49364 50260 49756
rect 49644 49026 49924 49028
rect 49644 48974 49646 49026
rect 49698 48974 49924 49026
rect 49644 48972 49924 48974
rect 50092 49308 50260 49364
rect 50876 49698 50932 49710
rect 50876 49646 50878 49698
rect 50930 49646 50932 49698
rect 50876 49364 50932 49646
rect 49644 48962 49700 48972
rect 49532 48468 49588 48478
rect 49420 48466 49588 48468
rect 49420 48414 49534 48466
rect 49586 48414 49588 48466
rect 49420 48412 49588 48414
rect 49532 48402 49588 48412
rect 49644 48130 49700 48142
rect 49644 48078 49646 48130
rect 49698 48078 49700 48130
rect 48860 47234 48916 47246
rect 48860 47182 48862 47234
rect 48914 47182 48916 47234
rect 48860 47124 48916 47182
rect 48860 47058 48916 47068
rect 48636 46946 48692 46956
rect 48524 46834 48580 46844
rect 49644 46898 49700 48078
rect 49644 46846 49646 46898
rect 49698 46846 49700 46898
rect 49644 46834 49700 46846
rect 49980 46900 50036 46910
rect 49980 46806 50036 46844
rect 47964 46562 48244 46564
rect 47964 46510 47966 46562
rect 48018 46510 48244 46562
rect 47964 46508 48244 46510
rect 48748 46676 48804 46686
rect 47964 46340 48020 46508
rect 47628 46284 48020 46340
rect 47516 45220 47572 45230
rect 47628 45220 47684 46284
rect 48748 46002 48804 46620
rect 49532 46676 49588 46686
rect 49532 46582 49588 46620
rect 49756 46674 49812 46686
rect 49756 46622 49758 46674
rect 49810 46622 49812 46674
rect 49756 46004 49812 46622
rect 48748 45950 48750 46002
rect 48802 45950 48804 46002
rect 48748 45938 48804 45950
rect 49532 45948 49812 46004
rect 47516 45218 47684 45220
rect 47516 45166 47518 45218
rect 47570 45166 47684 45218
rect 47516 45164 47684 45166
rect 48972 45892 49028 45902
rect 49532 45892 49588 45948
rect 48972 45890 49588 45892
rect 48972 45838 48974 45890
rect 49026 45838 49588 45890
rect 48972 45836 49588 45838
rect 47516 45154 47572 45164
rect 47740 45108 47796 45118
rect 47404 43374 47406 43426
rect 47458 43374 47460 43426
rect 45836 42466 45892 42476
rect 45948 42754 46676 42756
rect 45948 42702 46062 42754
rect 46114 42702 46676 42754
rect 45948 42700 46676 42702
rect 46732 43316 46788 43326
rect 45724 41972 45780 41982
rect 45724 41878 45780 41916
rect 45276 41858 45332 41870
rect 45276 41806 45278 41858
rect 45330 41806 45332 41858
rect 45276 41748 45332 41806
rect 45276 41682 45332 41692
rect 45612 41748 45668 41758
rect 45500 40962 45556 40974
rect 45500 40910 45502 40962
rect 45554 40910 45556 40962
rect 45500 40180 45556 40910
rect 45500 40114 45556 40124
rect 45612 40402 45668 41692
rect 45612 40350 45614 40402
rect 45666 40350 45668 40402
rect 45500 39732 45556 39742
rect 45612 39732 45668 40350
rect 45500 39730 45668 39732
rect 45500 39678 45502 39730
rect 45554 39678 45668 39730
rect 45500 39676 45668 39678
rect 45724 40290 45780 40302
rect 45724 40238 45726 40290
rect 45778 40238 45780 40290
rect 45724 40180 45780 40238
rect 45500 39058 45556 39676
rect 45500 39006 45502 39058
rect 45554 39006 45556 39058
rect 45500 38994 45556 39006
rect 45724 39618 45780 40124
rect 45724 39566 45726 39618
rect 45778 39566 45780 39618
rect 44492 35870 44494 35922
rect 44546 35870 44548 35922
rect 44492 35812 44548 35870
rect 44492 35746 44548 35756
rect 44604 38612 45220 38668
rect 45724 38724 45780 39566
rect 45724 38658 45780 38668
rect 45948 39396 46004 42700
rect 46060 42690 46116 42700
rect 46508 42532 46564 42542
rect 46508 42530 46676 42532
rect 46508 42478 46510 42530
rect 46562 42478 46676 42530
rect 46508 42476 46676 42478
rect 46508 42466 46564 42476
rect 46396 42084 46452 42094
rect 46172 41972 46228 41982
rect 46172 41186 46228 41916
rect 46396 41970 46452 42028
rect 46396 41918 46398 41970
rect 46450 41918 46452 41970
rect 46396 41906 46452 41918
rect 46620 41748 46676 42476
rect 46732 42084 46788 43260
rect 47404 42756 47460 43374
rect 47404 42690 47460 42700
rect 47628 43428 47684 43438
rect 46732 42018 46788 42028
rect 47404 42530 47460 42542
rect 47404 42478 47406 42530
rect 47458 42478 47460 42530
rect 46620 41746 46788 41748
rect 46620 41694 46622 41746
rect 46674 41694 46788 41746
rect 46620 41692 46788 41694
rect 46620 41682 46676 41692
rect 46172 41134 46174 41186
rect 46226 41134 46228 41186
rect 46172 40516 46228 41134
rect 46172 40450 46228 40460
rect 46060 40404 46116 40414
rect 46060 40178 46116 40348
rect 46060 40126 46062 40178
rect 46114 40126 46116 40178
rect 46060 40114 46116 40126
rect 46732 40292 46788 41692
rect 46844 41746 46900 41758
rect 46844 41694 46846 41746
rect 46898 41694 46900 41746
rect 46844 41076 46900 41694
rect 47292 41746 47348 41758
rect 47292 41694 47294 41746
rect 47346 41694 47348 41746
rect 47292 41636 47348 41694
rect 47404 41636 47460 42478
rect 47628 42530 47684 43372
rect 47740 42866 47796 45052
rect 48748 45108 48804 45118
rect 48748 45014 48804 45052
rect 48524 44996 48580 45006
rect 48524 44902 48580 44940
rect 48188 44882 48244 44894
rect 48188 44830 48190 44882
rect 48242 44830 48244 44882
rect 48188 44324 48244 44830
rect 48188 44258 48244 44268
rect 48300 44434 48356 44446
rect 48300 44382 48302 44434
rect 48354 44382 48356 44434
rect 48300 44212 48356 44382
rect 48300 44146 48356 44156
rect 48412 44322 48468 44334
rect 48412 44270 48414 44322
rect 48466 44270 48468 44322
rect 48412 44100 48468 44270
rect 48412 44034 48468 44044
rect 47852 43428 47908 43438
rect 47852 43334 47908 43372
rect 48412 43426 48468 43438
rect 48412 43374 48414 43426
rect 48466 43374 48468 43426
rect 47740 42814 47742 42866
rect 47794 42814 47796 42866
rect 47740 42802 47796 42814
rect 48188 42756 48244 42766
rect 47628 42478 47630 42530
rect 47682 42478 47684 42530
rect 47628 41860 47684 42478
rect 47852 42530 47908 42542
rect 47852 42478 47854 42530
rect 47906 42478 47908 42530
rect 47852 41972 47908 42478
rect 47852 41906 47908 41916
rect 48188 42532 48244 42700
rect 48300 42532 48356 42542
rect 48188 42530 48356 42532
rect 48188 42478 48302 42530
rect 48354 42478 48356 42530
rect 48188 42476 48356 42478
rect 47628 41794 47684 41804
rect 47292 41580 47572 41636
rect 46956 41300 47012 41310
rect 46956 41206 47012 41244
rect 47516 41188 47572 41580
rect 48076 41188 48132 41198
rect 47516 41186 48132 41188
rect 47516 41134 48078 41186
rect 48130 41134 48132 41186
rect 47516 41132 48132 41134
rect 48076 41122 48132 41132
rect 46844 41010 46900 41020
rect 47404 41076 47460 41086
rect 47460 41020 47908 41076
rect 47404 40944 47460 41020
rect 47852 40964 47908 41020
rect 48188 40964 48244 42476
rect 48300 42466 48356 42476
rect 48412 42532 48468 43374
rect 48860 43426 48916 43438
rect 48860 43374 48862 43426
rect 48914 43374 48916 43426
rect 48412 42466 48468 42476
rect 48748 42754 48804 42766
rect 48748 42702 48750 42754
rect 48802 42702 48804 42754
rect 48748 42082 48804 42702
rect 48860 42196 48916 43374
rect 48972 42978 49028 45836
rect 49644 45780 49700 45790
rect 49644 45778 49812 45780
rect 49644 45726 49646 45778
rect 49698 45726 49812 45778
rect 49644 45724 49812 45726
rect 49644 45714 49700 45724
rect 49756 45108 49812 45724
rect 49868 45108 49924 45118
rect 49756 45052 49868 45108
rect 49868 45014 49924 45052
rect 49084 44996 49140 45006
rect 49084 44434 49140 44940
rect 49644 44996 49700 45006
rect 49644 44902 49700 44940
rect 50092 44884 50148 49308
rect 50876 49298 50932 49308
rect 51436 49698 51492 49710
rect 51436 49646 51438 49698
rect 51490 49646 51492 49698
rect 51436 49588 51492 49646
rect 51100 48804 51156 48814
rect 51100 48710 51156 48748
rect 51436 48804 51492 49532
rect 51772 49138 51828 50092
rect 52108 50036 52164 53900
rect 52220 53842 52276 53854
rect 52220 53790 52222 53842
rect 52274 53790 52276 53842
rect 52220 53732 52276 53790
rect 52220 53666 52276 53676
rect 52556 53732 52612 54462
rect 52556 53666 52612 53676
rect 53004 54516 53060 54526
rect 52668 52276 52724 52286
rect 52444 52164 52500 52174
rect 52444 52050 52500 52108
rect 52444 51998 52446 52050
rect 52498 51998 52500 52050
rect 52332 51492 52388 51502
rect 52444 51492 52500 51998
rect 52556 51940 52612 51950
rect 52668 51940 52724 52220
rect 52780 52164 52836 52174
rect 53004 52164 53060 54460
rect 53228 52946 53284 54572
rect 53228 52894 53230 52946
rect 53282 52894 53284 52946
rect 52780 52162 53060 52164
rect 52780 52110 52782 52162
rect 52834 52110 53060 52162
rect 52780 52108 53060 52110
rect 53116 52834 53172 52846
rect 53116 52782 53118 52834
rect 53170 52782 53172 52834
rect 52780 52098 52836 52108
rect 52556 51938 52724 51940
rect 52556 51886 52558 51938
rect 52610 51886 52724 51938
rect 52556 51884 52724 51886
rect 52556 51874 52612 51884
rect 52332 51490 52500 51492
rect 52332 51438 52334 51490
rect 52386 51438 52500 51490
rect 52332 51436 52500 51438
rect 52332 51426 52388 51436
rect 51996 49980 52108 50036
rect 51884 49588 51940 49598
rect 51884 49494 51940 49532
rect 51772 49086 51774 49138
rect 51826 49086 51828 49138
rect 51772 49074 51828 49086
rect 51660 49026 51716 49038
rect 51660 48974 51662 49026
rect 51714 48974 51716 49026
rect 51660 48916 51716 48974
rect 51996 49026 52052 49980
rect 52108 49970 52164 49980
rect 52556 50260 52612 50270
rect 52556 50034 52612 50204
rect 52668 50148 52724 51884
rect 53116 50260 53172 52782
rect 53228 52836 53284 52894
rect 53340 52948 53396 54684
rect 53452 54674 53508 54684
rect 54348 54628 54404 54638
rect 54348 54534 54404 54572
rect 53676 54516 53732 54526
rect 53676 54422 53732 54460
rect 54236 54516 54292 54526
rect 54236 54422 54292 54460
rect 53564 54402 53620 54414
rect 53564 54350 53566 54402
rect 53618 54350 53620 54402
rect 53452 53956 53508 53966
rect 53452 53730 53508 53900
rect 53452 53678 53454 53730
rect 53506 53678 53508 53730
rect 53452 53666 53508 53678
rect 53564 53730 53620 54350
rect 53564 53678 53566 53730
rect 53618 53678 53620 53730
rect 53564 53666 53620 53678
rect 53900 53732 53956 53742
rect 53900 53638 53956 53676
rect 53564 52948 53620 52958
rect 53340 52946 53620 52948
rect 53340 52894 53566 52946
rect 53618 52894 53620 52946
rect 53340 52892 53620 52894
rect 53564 52882 53620 52892
rect 53228 52780 53508 52836
rect 53452 52274 53508 52780
rect 53452 52222 53454 52274
rect 53506 52222 53508 52274
rect 53452 52210 53508 52222
rect 53900 52276 53956 52286
rect 53564 52164 53620 52174
rect 53564 52070 53620 52108
rect 53900 52162 53956 52220
rect 53900 52110 53902 52162
rect 53954 52110 53956 52162
rect 53900 52098 53956 52110
rect 55132 51602 55188 55916
rect 55244 55076 55300 56476
rect 57148 55860 57204 55870
rect 55244 55010 55300 55020
rect 57036 55076 57092 55086
rect 55132 51550 55134 51602
rect 55186 51550 55188 51602
rect 55132 51538 55188 51550
rect 55692 51268 55748 51278
rect 56252 51268 56308 51278
rect 55580 51266 55972 51268
rect 55580 51214 55694 51266
rect 55746 51214 55972 51266
rect 55580 51212 55972 51214
rect 55468 51154 55524 51166
rect 55468 51102 55470 51154
rect 55522 51102 55524 51154
rect 53788 50596 53844 50606
rect 53788 50484 53844 50540
rect 54236 50596 54292 50606
rect 54236 50502 54292 50540
rect 54460 50594 54516 50606
rect 54460 50542 54462 50594
rect 54514 50542 54516 50594
rect 53564 50428 53844 50484
rect 53900 50484 53956 50494
rect 53116 50194 53172 50204
rect 53452 50372 53508 50382
rect 52668 50092 52836 50148
rect 52556 49982 52558 50034
rect 52610 49982 52612 50034
rect 52556 49970 52612 49982
rect 51996 48974 51998 49026
rect 52050 48974 52052 49026
rect 51996 48962 52052 48974
rect 52220 49810 52276 49822
rect 52220 49758 52222 49810
rect 52274 49758 52276 49810
rect 51660 48850 51716 48860
rect 51436 48738 51492 48748
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 51660 48242 51716 48254
rect 51996 48244 52052 48254
rect 51660 48190 51662 48242
rect 51714 48190 51716 48242
rect 49084 44382 49086 44434
rect 49138 44382 49140 44434
rect 49084 44370 49140 44382
rect 49756 44828 50148 44884
rect 50204 48132 50260 48142
rect 50652 48132 50708 48142
rect 50204 48130 50708 48132
rect 50204 48078 50206 48130
rect 50258 48078 50654 48130
rect 50706 48078 50708 48130
rect 50204 48076 50708 48078
rect 50204 47236 50260 48076
rect 50652 48066 50708 48076
rect 51212 48132 51268 48142
rect 51660 48132 51716 48190
rect 51212 48130 51716 48132
rect 51212 48078 51214 48130
rect 51266 48078 51716 48130
rect 51212 48076 51716 48078
rect 51772 48242 52052 48244
rect 51772 48190 51998 48242
rect 52050 48190 52052 48242
rect 51772 48188 52052 48190
rect 52220 48244 52276 49758
rect 52332 49810 52388 49822
rect 52332 49758 52334 49810
rect 52386 49758 52388 49810
rect 52332 49364 52388 49758
rect 52332 49298 52388 49308
rect 52444 49698 52500 49710
rect 52444 49646 52446 49698
rect 52498 49646 52500 49698
rect 52444 49252 52500 49646
rect 52668 49252 52724 49262
rect 52444 49250 52724 49252
rect 52444 49198 52670 49250
rect 52722 49198 52724 49250
rect 52444 49196 52724 49198
rect 52668 49186 52724 49196
rect 52556 49026 52612 49038
rect 52556 48974 52558 49026
rect 52610 48974 52612 49026
rect 52332 48916 52388 48926
rect 52332 48822 52388 48860
rect 52556 48466 52612 48974
rect 52556 48414 52558 48466
rect 52610 48414 52612 48466
rect 52556 48402 52612 48414
rect 52668 48468 52724 48478
rect 52668 48354 52724 48412
rect 52668 48302 52670 48354
rect 52722 48302 52724 48354
rect 52668 48290 52724 48302
rect 52444 48244 52500 48254
rect 52220 48188 52444 48244
rect 51212 48066 51268 48076
rect 50876 48018 50932 48030
rect 50876 47966 50878 48018
rect 50930 47966 50932 48018
rect 50876 47460 50932 47966
rect 50876 47394 50932 47404
rect 51660 47458 51716 47470
rect 51660 47406 51662 47458
rect 51714 47406 51716 47458
rect 49756 44434 49812 44828
rect 49756 44382 49758 44434
rect 49810 44382 49812 44434
rect 49756 44370 49812 44382
rect 49868 44322 49924 44334
rect 49868 44270 49870 44322
rect 49922 44270 49924 44322
rect 49644 44212 49700 44222
rect 49644 44118 49700 44156
rect 49868 44100 49924 44270
rect 50092 44324 50148 44334
rect 50092 44230 50148 44268
rect 49868 44034 49924 44044
rect 50204 43708 50260 47180
rect 51100 47236 51156 47246
rect 51100 47142 51156 47180
rect 51660 47236 51716 47406
rect 51660 47170 51716 47180
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 51324 45890 51380 45902
rect 51324 45838 51326 45890
rect 51378 45838 51380 45890
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 50540 44996 50596 45006
rect 50540 44902 50596 44940
rect 51100 44996 51156 45006
rect 50876 44884 50932 44894
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 50204 43652 50372 43708
rect 48972 42926 48974 42978
rect 49026 42926 49028 42978
rect 48972 42914 49028 42926
rect 49084 42532 49140 42542
rect 49084 42438 49140 42476
rect 49308 42530 49364 42542
rect 49308 42478 49310 42530
rect 49362 42478 49364 42530
rect 49308 42196 49364 42478
rect 48860 42140 49364 42196
rect 49532 42532 49588 42542
rect 48748 42030 48750 42082
rect 48802 42030 48804 42082
rect 48748 42018 48804 42030
rect 48300 41970 48356 41982
rect 48300 41918 48302 41970
rect 48354 41918 48356 41970
rect 48300 41860 48356 41918
rect 48300 41794 48356 41804
rect 48636 41972 48692 41982
rect 48636 41410 48692 41916
rect 48636 41358 48638 41410
rect 48690 41358 48692 41410
rect 48636 41346 48692 41358
rect 47852 40908 48244 40964
rect 49084 41300 49140 42140
rect 49084 40964 49140 41244
rect 49196 41188 49252 41198
rect 49420 41188 49476 41198
rect 49196 41186 49364 41188
rect 49196 41134 49198 41186
rect 49250 41134 49364 41186
rect 49196 41132 49364 41134
rect 49196 41122 49252 41132
rect 49196 40964 49252 40974
rect 49084 40908 49196 40964
rect 46844 40516 46900 40526
rect 46844 40422 46900 40460
rect 47180 40516 47236 40526
rect 46732 39620 46788 40236
rect 46060 39396 46116 39406
rect 45948 39394 46116 39396
rect 45948 39342 46062 39394
rect 46114 39342 46116 39394
rect 45948 39340 46116 39342
rect 44380 34692 44436 34702
rect 44380 34598 44436 34636
rect 44492 34020 44548 34030
rect 44492 33926 44548 33964
rect 44380 33122 44436 33134
rect 44380 33070 44382 33122
rect 44434 33070 44436 33122
rect 44380 33012 44436 33070
rect 44380 31890 44436 32956
rect 44380 31838 44382 31890
rect 44434 31838 44436 31890
rect 44268 31668 44324 31678
rect 44268 31218 44324 31612
rect 44268 31166 44270 31218
rect 44322 31166 44324 31218
rect 44268 31154 44324 31166
rect 44380 30770 44436 31838
rect 44380 30718 44382 30770
rect 44434 30718 44436 30770
rect 44380 30706 44436 30718
rect 44492 32676 44548 32686
rect 44156 29698 44212 29708
rect 44380 29540 44436 29550
rect 43484 29538 44436 29540
rect 43484 29486 44382 29538
rect 44434 29486 44436 29538
rect 43484 29484 44436 29486
rect 43484 29428 43540 29484
rect 44380 29474 44436 29484
rect 43036 29426 43540 29428
rect 43036 29374 43486 29426
rect 43538 29374 43540 29426
rect 43036 29372 43540 29374
rect 42364 28578 42420 28588
rect 42588 29314 42644 29326
rect 42588 29262 42590 29314
rect 42642 29262 42644 29314
rect 41468 28252 41636 28308
rect 41356 27412 41412 27580
rect 41468 27746 41524 27758
rect 41468 27694 41470 27746
rect 41522 27694 41524 27746
rect 41468 27524 41524 27694
rect 41468 27458 41524 27468
rect 41356 27346 41412 27356
rect 41356 27188 41412 27198
rect 41356 27094 41412 27132
rect 41580 26908 41636 28252
rect 41692 28242 41748 28252
rect 41916 28252 42084 28308
rect 42364 28418 42420 28430
rect 42364 28366 42366 28418
rect 42418 28366 42420 28418
rect 41916 28082 41972 28252
rect 41916 28030 41918 28082
rect 41970 28030 41972 28082
rect 41916 28018 41972 28030
rect 42364 28084 42420 28366
rect 42588 28420 42644 29262
rect 42924 28644 42980 28654
rect 42924 28550 42980 28588
rect 42588 28354 42644 28364
rect 41804 27524 41860 27534
rect 41804 27186 41860 27468
rect 41804 27134 41806 27186
rect 41858 27134 41860 27186
rect 41804 27122 41860 27134
rect 41132 25106 41188 25116
rect 41244 26852 41300 26862
rect 41132 24164 41188 24174
rect 41132 24070 41188 24108
rect 40460 24050 40628 24052
rect 40460 23998 40462 24050
rect 40514 23998 40628 24050
rect 40460 23996 40628 23998
rect 40460 23986 40516 23996
rect 40908 23940 40964 23950
rect 40908 23846 40964 23884
rect 39788 22866 39844 22876
rect 39900 23772 40068 23828
rect 40572 23828 40628 23838
rect 39900 23378 39956 23772
rect 39900 23326 39902 23378
rect 39954 23326 39956 23378
rect 39900 22484 39956 23326
rect 40012 23380 40068 23390
rect 40012 23286 40068 23324
rect 40124 23154 40180 23166
rect 40124 23102 40126 23154
rect 40178 23102 40180 23154
rect 40124 22932 40180 23102
rect 40124 22866 40180 22876
rect 40236 23154 40292 23166
rect 40236 23102 40238 23154
rect 40290 23102 40292 23154
rect 39900 22418 39956 22428
rect 40124 22258 40180 22270
rect 40124 22206 40126 22258
rect 40178 22206 40180 22258
rect 39564 21868 39732 21924
rect 39452 20972 39620 21028
rect 39452 20580 39508 20590
rect 39452 20486 39508 20524
rect 39452 19906 39508 19918
rect 39452 19854 39454 19906
rect 39506 19854 39508 19906
rect 39452 19460 39508 19854
rect 39452 19394 39508 19404
rect 39340 19348 39396 19358
rect 39340 19254 39396 19292
rect 39452 19012 39508 19022
rect 39452 16324 39508 18956
rect 39452 16258 39508 16268
rect 39564 17108 39620 20972
rect 39676 19572 39732 21868
rect 40124 21812 40180 22206
rect 40124 21746 40180 21756
rect 39788 21586 39844 21598
rect 39788 21534 39790 21586
rect 39842 21534 39844 21586
rect 39788 21476 39844 21534
rect 39788 21028 39844 21420
rect 39788 20962 39844 20972
rect 39900 21026 39956 21038
rect 39900 20974 39902 21026
rect 39954 20974 39956 21026
rect 39900 20914 39956 20974
rect 39900 20862 39902 20914
rect 39954 20862 39956 20914
rect 39900 20850 39956 20862
rect 40012 21028 40068 21038
rect 40012 20242 40068 20972
rect 40236 21028 40292 23102
rect 40348 23156 40404 23166
rect 40348 22148 40404 23100
rect 40572 22372 40628 23772
rect 40796 23042 40852 23054
rect 40796 22990 40798 23042
rect 40850 22990 40852 23042
rect 40796 22932 40852 22990
rect 40796 22866 40852 22876
rect 41132 22594 41188 22606
rect 41132 22542 41134 22594
rect 41186 22542 41188 22594
rect 41132 22372 41188 22542
rect 40572 22316 41188 22372
rect 40572 22258 40628 22316
rect 40572 22206 40574 22258
rect 40626 22206 40628 22258
rect 40572 22194 40628 22206
rect 40460 22148 40516 22158
rect 40348 22146 40460 22148
rect 40348 22094 40350 22146
rect 40402 22094 40460 22146
rect 40348 22092 40460 22094
rect 40348 22082 40404 22092
rect 40236 20962 40292 20972
rect 40348 21364 40404 21374
rect 40012 20190 40014 20242
rect 40066 20190 40068 20242
rect 40012 20178 40068 20190
rect 40124 20132 40180 20142
rect 39676 19516 39844 19572
rect 39676 19348 39732 19358
rect 39676 18674 39732 19292
rect 39676 18622 39678 18674
rect 39730 18622 39732 18674
rect 39676 18610 39732 18622
rect 39788 18452 39844 19516
rect 40124 19012 40180 20076
rect 40348 19908 40404 21308
rect 40460 20690 40516 22092
rect 40684 22146 40740 22158
rect 41020 22148 41076 22158
rect 40684 22094 40686 22146
rect 40738 22094 40740 22146
rect 40460 20638 40462 20690
rect 40514 20638 40516 20690
rect 40460 20132 40516 20638
rect 40572 21812 40628 21822
rect 40572 20356 40628 21756
rect 40684 21364 40740 22094
rect 40684 21298 40740 21308
rect 40908 22146 41076 22148
rect 40908 22094 41022 22146
rect 41074 22094 41076 22146
rect 40908 22092 41076 22094
rect 40684 21028 40740 21038
rect 40908 21028 40964 22092
rect 41020 22082 41076 22092
rect 40740 20972 40964 21028
rect 40684 20934 40740 20972
rect 40572 20290 40628 20300
rect 40796 20356 40852 20366
rect 40460 20066 40516 20076
rect 40348 19906 40516 19908
rect 40348 19854 40350 19906
rect 40402 19854 40516 19906
rect 40348 19852 40516 19854
rect 40348 19842 40404 19852
rect 40348 19236 40404 19246
rect 40236 19012 40292 19022
rect 40124 18956 40236 19012
rect 40236 18918 40292 18956
rect 39788 18386 39844 18396
rect 40236 18452 40292 18462
rect 40236 18358 40292 18396
rect 40236 17668 40292 17678
rect 40348 17668 40404 19180
rect 40460 18228 40516 19852
rect 40796 19572 40852 20300
rect 40908 20242 40964 20972
rect 41020 20804 41076 20814
rect 41020 20710 41076 20748
rect 40908 20190 40910 20242
rect 40962 20190 40964 20242
rect 40908 20178 40964 20190
rect 40796 19516 40964 19572
rect 40908 19346 40964 19516
rect 40908 19294 40910 19346
rect 40962 19294 40964 19346
rect 40908 19236 40964 19294
rect 40908 19170 40964 19180
rect 41020 19348 41076 19358
rect 40908 18900 40964 18910
rect 40460 18162 40516 18172
rect 40796 18788 40852 18798
rect 40236 17666 40404 17668
rect 40236 17614 40238 17666
rect 40290 17614 40404 17666
rect 40236 17612 40404 17614
rect 39676 17556 39732 17566
rect 39676 17554 40068 17556
rect 39676 17502 39678 17554
rect 39730 17502 40068 17554
rect 39676 17500 40068 17502
rect 39676 17490 39732 17500
rect 39564 16212 39620 17052
rect 39564 16146 39620 16156
rect 39788 15986 39844 15998
rect 39788 15934 39790 15986
rect 39842 15934 39844 15986
rect 38892 15486 38894 15538
rect 38946 15486 38948 15538
rect 38892 15474 38948 15486
rect 39004 15596 39284 15652
rect 39340 15874 39396 15886
rect 39340 15822 39342 15874
rect 39394 15822 39396 15874
rect 38332 15316 38388 15354
rect 38332 15250 38388 15260
rect 38332 15090 38388 15102
rect 38332 15038 38334 15090
rect 38386 15038 38388 15090
rect 38332 14530 38388 15038
rect 38332 14478 38334 14530
rect 38386 14478 38388 14530
rect 38332 14466 38388 14478
rect 38108 14366 38110 14418
rect 38162 14366 38164 14418
rect 38108 14354 38164 14366
rect 37996 13806 37998 13858
rect 38050 13806 38052 13858
rect 37996 13794 38052 13806
rect 38332 13860 38388 13870
rect 38332 13766 38388 13804
rect 38220 13636 38276 13646
rect 38220 13542 38276 13580
rect 37772 13412 37828 13422
rect 37660 13074 37716 13086
rect 37660 13022 37662 13074
rect 37714 13022 37716 13074
rect 37548 12850 37604 12862
rect 37548 12798 37550 12850
rect 37602 12798 37604 12850
rect 37324 12740 37380 12750
rect 36988 12460 37156 12516
rect 35868 12292 35924 12302
rect 35868 11282 35924 12236
rect 36876 12290 36932 12302
rect 36876 12238 36878 12290
rect 36930 12238 36932 12290
rect 36652 12180 36708 12190
rect 36652 12086 36708 12124
rect 36876 11956 36932 12238
rect 36988 12292 37044 12302
rect 36988 12198 37044 12236
rect 36876 11890 36932 11900
rect 35868 11230 35870 11282
rect 35922 11230 35924 11282
rect 35868 11218 35924 11230
rect 36540 10612 36596 10622
rect 36540 10518 36596 10556
rect 35308 9548 35812 9604
rect 35980 10498 36036 10510
rect 35980 10446 35982 10498
rect 36034 10446 36036 10498
rect 35308 9492 35364 9548
rect 34860 9202 34916 9212
rect 34972 9436 35364 9492
rect 34972 9266 35028 9436
rect 34972 9214 34974 9266
rect 35026 9214 35028 9266
rect 34972 8372 35028 9214
rect 35644 9380 35700 9390
rect 35644 9266 35700 9324
rect 35644 9214 35646 9266
rect 35698 9214 35700 9266
rect 35644 9202 35700 9214
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35980 8484 36036 10446
rect 36316 10164 36372 10174
rect 36204 9380 36260 9390
rect 36204 9154 36260 9324
rect 36204 9102 36206 9154
rect 36258 9102 36260 9154
rect 36204 9090 36260 9102
rect 36316 9266 36372 10108
rect 37100 10164 37156 12460
rect 37324 12178 37380 12684
rect 37324 12126 37326 12178
rect 37378 12126 37380 12178
rect 37324 12114 37380 12126
rect 37548 12180 37604 12798
rect 37548 12114 37604 12124
rect 37436 12066 37492 12078
rect 37436 12014 37438 12066
rect 37490 12014 37492 12066
rect 37436 10612 37492 12014
rect 37548 10612 37604 10622
rect 37436 10610 37604 10612
rect 37436 10558 37550 10610
rect 37602 10558 37604 10610
rect 37436 10556 37604 10558
rect 37660 10612 37716 13022
rect 37772 12962 37828 13356
rect 38892 13412 38948 13422
rect 38892 13074 38948 13356
rect 38892 13022 38894 13074
rect 38946 13022 38948 13074
rect 38892 13010 38948 13022
rect 37772 12910 37774 12962
rect 37826 12910 37828 12962
rect 37772 12898 37828 12910
rect 37996 12740 38052 12750
rect 38444 12740 38500 12750
rect 37884 12738 38052 12740
rect 37884 12686 37998 12738
rect 38050 12686 38052 12738
rect 37884 12684 38052 12686
rect 37884 12066 37940 12684
rect 37996 12674 38052 12684
rect 38332 12738 38500 12740
rect 38332 12686 38446 12738
rect 38498 12686 38500 12738
rect 38332 12684 38500 12686
rect 37884 12014 37886 12066
rect 37938 12014 37940 12066
rect 37884 11956 37940 12014
rect 37884 11890 37940 11900
rect 38332 12066 38388 12684
rect 38444 12674 38500 12684
rect 38556 12740 38612 12750
rect 38332 12014 38334 12066
rect 38386 12014 38388 12066
rect 38332 11956 38388 12014
rect 38332 11890 38388 11900
rect 38108 11284 38164 11294
rect 38108 11282 38276 11284
rect 38108 11230 38110 11282
rect 38162 11230 38276 11282
rect 38108 11228 38276 11230
rect 38108 11218 38164 11228
rect 37772 10612 37828 10622
rect 37660 10610 37828 10612
rect 37660 10558 37774 10610
rect 37826 10558 37828 10610
rect 37660 10556 37828 10558
rect 37548 10546 37604 10556
rect 37772 10546 37828 10556
rect 37100 10098 37156 10108
rect 38108 10386 38164 10398
rect 38108 10334 38110 10386
rect 38162 10334 38164 10386
rect 38108 10052 38164 10334
rect 38108 9986 38164 9996
rect 36316 9214 36318 9266
rect 36370 9214 36372 9266
rect 35980 8418 36036 8428
rect 34972 8306 35028 8316
rect 35196 8370 35252 8382
rect 35196 8318 35198 8370
rect 35250 8318 35252 8370
rect 34636 8036 34692 8046
rect 34636 8034 34804 8036
rect 34636 7982 34638 8034
rect 34690 7982 34804 8034
rect 34636 7980 34804 7982
rect 34636 7970 34692 7980
rect 34748 7586 34804 7980
rect 34748 7534 34750 7586
rect 34802 7534 34804 7586
rect 34636 7250 34692 7262
rect 34636 7198 34638 7250
rect 34690 7198 34692 7250
rect 34636 6802 34692 7198
rect 34636 6750 34638 6802
rect 34690 6750 34692 6802
rect 34636 6738 34692 6750
rect 34748 5908 34804 7534
rect 34972 7588 35028 7598
rect 35196 7588 35252 8318
rect 35308 8372 35364 8382
rect 35308 8146 35364 8316
rect 35532 8260 35588 8270
rect 35532 8166 35588 8204
rect 35980 8260 36036 8270
rect 35980 8166 36036 8204
rect 35308 8094 35310 8146
rect 35362 8094 35364 8146
rect 35308 8082 35364 8094
rect 36316 8148 36372 9214
rect 37436 9940 37492 9950
rect 37436 9042 37492 9884
rect 37884 9940 37940 9950
rect 37884 9826 37940 9884
rect 37884 9774 37886 9826
rect 37938 9774 37940 9826
rect 37884 9762 37940 9774
rect 37996 9828 38052 9838
rect 37996 9734 38052 9772
rect 37436 8990 37438 9042
rect 37490 8990 37492 9042
rect 37436 8978 37492 8990
rect 37548 9716 37604 9726
rect 37548 8930 37604 9660
rect 37548 8878 37550 8930
rect 37602 8878 37604 8930
rect 37548 8866 37604 8878
rect 37772 9602 37828 9614
rect 37772 9550 37774 9602
rect 37826 9550 37828 9602
rect 36316 8082 36372 8092
rect 37324 8484 37380 8494
rect 34972 7586 35252 7588
rect 34972 7534 34974 7586
rect 35026 7534 35252 7586
rect 34972 7532 35252 7534
rect 37324 7586 37380 8428
rect 37772 8260 37828 9550
rect 37884 9044 37940 9054
rect 37884 8950 37940 8988
rect 38108 8484 38164 8494
rect 38108 8370 38164 8428
rect 38108 8318 38110 8370
rect 38162 8318 38164 8370
rect 38108 8306 38164 8318
rect 37884 8260 37940 8270
rect 37324 7534 37326 7586
rect 37378 7534 37380 7586
rect 34860 6692 34916 6702
rect 34860 6598 34916 6636
rect 34748 5842 34804 5852
rect 34860 5908 34916 5918
rect 34972 5908 35028 7532
rect 37324 7522 37380 7534
rect 37660 8258 37940 8260
rect 37660 8206 37886 8258
rect 37938 8206 37940 8258
rect 37660 8204 37940 8206
rect 37660 7474 37716 8204
rect 37884 8194 37940 8204
rect 37660 7422 37662 7474
rect 37714 7422 37716 7474
rect 37660 7410 37716 7422
rect 37660 7250 37716 7262
rect 37660 7198 37662 7250
rect 37714 7198 37716 7250
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 34860 5906 35028 5908
rect 34860 5854 34862 5906
rect 34914 5854 35028 5906
rect 34860 5852 35028 5854
rect 35084 6692 35140 6702
rect 35084 5906 35140 6636
rect 35980 6692 36036 6702
rect 35980 6598 36036 6636
rect 35532 6578 35588 6590
rect 35532 6526 35534 6578
rect 35586 6526 35588 6578
rect 35532 6244 35588 6526
rect 35532 6188 35812 6244
rect 35532 6020 35588 6030
rect 35532 5926 35588 5964
rect 35084 5854 35086 5906
rect 35138 5854 35140 5906
rect 34860 5842 34916 5852
rect 35084 5842 35140 5854
rect 35308 5908 35364 5918
rect 35308 5814 35364 5852
rect 35756 5908 35812 6188
rect 36988 6020 37044 6030
rect 36540 5908 36596 5918
rect 35756 5906 36596 5908
rect 35756 5854 35758 5906
rect 35810 5854 36542 5906
rect 36594 5854 36596 5906
rect 35756 5852 36596 5854
rect 35756 5842 35812 5852
rect 36540 5842 36596 5852
rect 36988 5906 37044 5964
rect 36988 5854 36990 5906
rect 37042 5854 37044 5906
rect 36988 5842 37044 5854
rect 37660 5908 37716 7198
rect 37660 5842 37716 5852
rect 35644 5796 35700 5806
rect 35644 5702 35700 5740
rect 37436 5794 37492 5806
rect 37436 5742 37438 5794
rect 37490 5742 37492 5794
rect 34524 5628 34804 5684
rect 34188 5182 34190 5234
rect 34242 5182 34244 5234
rect 34188 5170 34244 5182
rect 34748 5236 34804 5628
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 36652 5236 36708 5246
rect 34748 5234 34916 5236
rect 34748 5182 34750 5234
rect 34802 5182 34916 5234
rect 34748 5180 34916 5182
rect 34748 5170 34804 5180
rect 33964 4946 34020 4956
rect 34412 4788 34468 4798
rect 33516 3378 33572 3388
rect 33628 4450 33684 4462
rect 33628 4398 33630 4450
rect 33682 4398 33684 4450
rect 30716 3278 30718 3330
rect 30770 3278 30772 3330
rect 30716 3266 30772 3278
rect 33628 3332 33684 4398
rect 34076 4452 34132 4462
rect 33852 4338 33908 4350
rect 33852 4286 33854 4338
rect 33906 4286 33908 4338
rect 33852 3668 33908 4286
rect 33852 3602 33908 3612
rect 34076 3666 34132 4396
rect 34412 4226 34468 4732
rect 34860 4452 34916 5180
rect 34972 5122 35028 5134
rect 34972 5070 34974 5122
rect 35026 5070 35028 5122
rect 34972 5012 35028 5070
rect 35644 5124 35700 5134
rect 35644 5030 35700 5068
rect 36428 5124 36484 5134
rect 36428 5030 36484 5068
rect 34972 4946 35028 4956
rect 35308 5012 35364 5022
rect 35196 4452 35252 4462
rect 34412 4174 34414 4226
rect 34466 4174 34468 4226
rect 34412 3780 34468 4174
rect 34412 3714 34468 3724
rect 34524 4450 35252 4452
rect 34524 4398 35198 4450
rect 35250 4398 35252 4450
rect 34524 4396 35252 4398
rect 34076 3614 34078 3666
rect 34130 3614 34132 3666
rect 34076 3602 34132 3614
rect 34524 3668 34580 4396
rect 35196 4386 35252 4396
rect 35308 4116 35364 4956
rect 36652 5010 36708 5180
rect 36652 4958 36654 5010
rect 36706 4958 36708 5010
rect 36652 4946 36708 4958
rect 36540 4898 36596 4910
rect 36540 4846 36542 4898
rect 36594 4846 36596 4898
rect 35532 4340 35588 4350
rect 36092 4340 36148 4350
rect 35532 4338 36148 4340
rect 35532 4286 35534 4338
rect 35586 4286 36094 4338
rect 36146 4286 36148 4338
rect 35532 4284 36148 4286
rect 35532 4274 35588 4284
rect 36092 4274 36148 4284
rect 36540 4340 36596 4846
rect 36540 4274 36596 4284
rect 37212 4340 37268 4350
rect 35420 4228 35476 4238
rect 35420 4134 35476 4172
rect 36204 4226 36260 4238
rect 36204 4174 36206 4226
rect 36258 4174 36260 4226
rect 35308 4050 35364 4060
rect 35532 4116 35588 4126
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 34524 3536 34580 3612
rect 35420 3668 35476 3678
rect 35532 3668 35588 4060
rect 36204 4116 36260 4174
rect 36988 4228 37044 4238
rect 36988 4134 37044 4172
rect 35420 3666 35588 3668
rect 35420 3614 35422 3666
rect 35474 3614 35588 3666
rect 35420 3612 35588 3614
rect 35756 3668 35812 3678
rect 35420 3602 35476 3612
rect 35756 3574 35812 3612
rect 36204 3666 36260 4060
rect 36204 3614 36206 3666
rect 36258 3614 36260 3666
rect 36204 3602 36260 3614
rect 37100 3556 37156 3566
rect 37212 3556 37268 4284
rect 37436 4340 37492 5742
rect 38220 5236 38276 11228
rect 38556 9940 38612 12684
rect 38892 12292 38948 12302
rect 39004 12292 39060 15596
rect 39228 15428 39284 15438
rect 39228 15334 39284 15372
rect 39340 15316 39396 15822
rect 39340 15250 39396 15260
rect 39788 15148 39844 15934
rect 39564 15092 39844 15148
rect 39900 15316 39956 15326
rect 39564 14418 39620 15092
rect 39564 14366 39566 14418
rect 39618 14366 39620 14418
rect 39564 13860 39620 14366
rect 39564 13794 39620 13804
rect 39676 14306 39732 14318
rect 39676 14254 39678 14306
rect 39730 14254 39732 14306
rect 39676 13076 39732 14254
rect 39788 13972 39844 13982
rect 39788 13878 39844 13916
rect 39900 13076 39956 15260
rect 40012 14084 40068 17500
rect 40124 16996 40180 17006
rect 40236 16996 40292 17612
rect 40348 17444 40404 17482
rect 40572 17444 40628 17454
rect 40348 17378 40404 17388
rect 40460 17442 40628 17444
rect 40460 17390 40574 17442
rect 40626 17390 40628 17442
rect 40460 17388 40628 17390
rect 40124 16994 40292 16996
rect 40124 16942 40126 16994
rect 40178 16942 40292 16994
rect 40124 16940 40292 16942
rect 40348 17220 40404 17230
rect 40348 17106 40404 17164
rect 40348 17054 40350 17106
rect 40402 17054 40404 17106
rect 40124 16100 40180 16940
rect 40124 16034 40180 16044
rect 40236 16436 40292 16446
rect 40236 16098 40292 16380
rect 40236 16046 40238 16098
rect 40290 16046 40292 16098
rect 40236 15428 40292 16046
rect 40236 15362 40292 15372
rect 40348 15314 40404 17054
rect 40348 15262 40350 15314
rect 40402 15262 40404 15314
rect 40348 15250 40404 15262
rect 40460 14980 40516 17388
rect 40572 17378 40628 17388
rect 40572 17108 40628 17118
rect 40572 17014 40628 17052
rect 40684 16660 40740 16670
rect 40684 16566 40740 16604
rect 40796 16436 40852 18732
rect 40908 18674 40964 18844
rect 40908 18622 40910 18674
rect 40962 18622 40964 18674
rect 40908 18610 40964 18622
rect 40908 17780 40964 17790
rect 41020 17780 41076 19292
rect 40908 17778 41076 17780
rect 40908 17726 40910 17778
rect 40962 17726 41076 17778
rect 40908 17724 41076 17726
rect 40908 17444 40964 17724
rect 40908 17378 40964 17388
rect 40460 14914 40516 14924
rect 40572 16380 40852 16436
rect 40012 14018 40068 14028
rect 39676 13010 39732 13020
rect 39788 13020 39956 13076
rect 40124 13972 40180 13982
rect 39788 12964 39844 13020
rect 39564 12852 39620 12862
rect 39788 12852 39844 12908
rect 39564 12850 39844 12852
rect 39564 12798 39566 12850
rect 39618 12798 39844 12850
rect 39564 12796 39844 12798
rect 40124 12962 40180 13916
rect 40124 12910 40126 12962
rect 40178 12910 40180 12962
rect 39564 12786 39620 12796
rect 39452 12740 39508 12750
rect 39452 12646 39508 12684
rect 39452 12292 39508 12302
rect 38892 12290 39172 12292
rect 38892 12238 38894 12290
rect 38946 12238 39172 12290
rect 38892 12236 39172 12238
rect 38892 12226 38948 12236
rect 39004 12066 39060 12078
rect 39004 12014 39006 12066
rect 39058 12014 39060 12066
rect 38780 11732 38836 11742
rect 38780 11394 38836 11676
rect 39004 11506 39060 12014
rect 39004 11454 39006 11506
rect 39058 11454 39060 11506
rect 39004 11442 39060 11454
rect 38780 11342 38782 11394
rect 38834 11342 38836 11394
rect 38780 11330 38836 11342
rect 39116 10388 39172 12236
rect 39452 12198 39508 12236
rect 39228 12178 39284 12190
rect 39228 12126 39230 12178
rect 39282 12126 39284 12178
rect 39228 11956 39284 12126
rect 39228 11890 39284 11900
rect 40012 11954 40068 11966
rect 40012 11902 40014 11954
rect 40066 11902 40068 11954
rect 39340 11732 39396 11742
rect 39340 10836 39396 11676
rect 40012 11732 40068 11902
rect 40012 11666 40068 11676
rect 40124 11282 40180 12910
rect 40236 12738 40292 12750
rect 40236 12686 40238 12738
rect 40290 12686 40292 12738
rect 40236 12292 40292 12686
rect 40236 12178 40292 12236
rect 40236 12126 40238 12178
rect 40290 12126 40292 12178
rect 40236 12114 40292 12126
rect 40348 12738 40404 12750
rect 40348 12686 40350 12738
rect 40402 12686 40404 12738
rect 40348 11956 40404 12686
rect 40460 12404 40516 12414
rect 40572 12404 40628 16380
rect 40684 16098 40740 16110
rect 40684 16046 40686 16098
rect 40738 16046 40740 16098
rect 40684 15428 40740 16046
rect 40796 15428 40852 15438
rect 40684 15426 40852 15428
rect 40684 15374 40798 15426
rect 40850 15374 40852 15426
rect 40684 15372 40852 15374
rect 40796 15316 40852 15372
rect 40796 15250 40852 15260
rect 41132 13972 41188 22316
rect 41244 19348 41300 26796
rect 41356 26852 41636 26908
rect 41916 27076 41972 27086
rect 41356 22148 41412 26852
rect 41804 26516 41860 26526
rect 41916 26516 41972 27020
rect 42252 26964 42308 27002
rect 42252 26898 42308 26908
rect 41804 26514 41972 26516
rect 41804 26462 41806 26514
rect 41858 26462 41972 26514
rect 41804 26460 41972 26462
rect 41804 26450 41860 26460
rect 42364 26404 42420 28028
rect 43036 28308 43092 29372
rect 43484 29362 43540 29372
rect 44044 29316 44100 29326
rect 43036 27860 43092 28252
rect 42700 27858 43092 27860
rect 42700 27806 43038 27858
rect 43090 27806 43092 27858
rect 42700 27804 43092 27806
rect 42700 27188 42756 27804
rect 43036 27794 43092 27804
rect 43148 29204 43204 29214
rect 43148 27746 43204 29148
rect 43148 27694 43150 27746
rect 43202 27694 43204 27746
rect 43148 27682 43204 27694
rect 43372 29204 43428 29214
rect 42700 27056 42756 27132
rect 42924 27636 42980 27646
rect 42252 26348 42420 26404
rect 41692 26290 41748 26302
rect 41692 26238 41694 26290
rect 41746 26238 41748 26290
rect 41692 26068 41748 26238
rect 41916 26292 41972 26302
rect 41916 26198 41972 26236
rect 41580 26012 41692 26068
rect 41468 25620 41524 25630
rect 41468 25526 41524 25564
rect 41468 24948 41524 24958
rect 41580 24948 41636 26012
rect 41692 26002 41748 26012
rect 42140 26178 42196 26190
rect 42140 26126 42142 26178
rect 42194 26126 42196 26178
rect 42140 25284 42196 26126
rect 42140 25218 42196 25228
rect 42252 25060 42308 26348
rect 42364 26180 42420 26190
rect 42364 26086 42420 26124
rect 42588 26068 42644 26078
rect 42476 26066 42644 26068
rect 42476 26014 42590 26066
rect 42642 26014 42644 26066
rect 42476 26012 42644 26014
rect 42364 25620 42420 25630
rect 42476 25620 42532 26012
rect 42588 26002 42644 26012
rect 42420 25564 42532 25620
rect 42364 25526 42420 25564
rect 42812 25508 42868 25518
rect 42812 25414 42868 25452
rect 42252 24994 42308 25004
rect 42364 25284 42420 25294
rect 41468 24946 41636 24948
rect 41468 24894 41470 24946
rect 41522 24894 41636 24946
rect 41468 24892 41636 24894
rect 41468 24882 41524 24892
rect 42364 24612 42420 25228
rect 42252 24610 42420 24612
rect 42252 24558 42366 24610
rect 42418 24558 42420 24610
rect 42252 24556 42420 24558
rect 41692 24164 41748 24174
rect 41468 23828 41524 23838
rect 41468 23734 41524 23772
rect 41692 23154 41748 24108
rect 41692 23102 41694 23154
rect 41746 23102 41748 23154
rect 41692 23090 41748 23102
rect 42028 23940 42084 23950
rect 42028 23154 42084 23884
rect 42028 23102 42030 23154
rect 42082 23102 42084 23154
rect 42028 23090 42084 23102
rect 41692 22932 41748 22942
rect 41468 22148 41524 22158
rect 41356 22092 41468 22148
rect 41468 22054 41524 22092
rect 41468 21588 41524 21598
rect 41468 21494 41524 21532
rect 41244 19282 41300 19292
rect 41468 19236 41524 19246
rect 41356 18676 41412 18686
rect 41356 17780 41412 18620
rect 41356 17648 41412 17724
rect 41468 17556 41524 19180
rect 41580 19124 41636 19134
rect 41692 19124 41748 22876
rect 41916 22594 41972 22606
rect 41916 22542 41918 22594
rect 41970 22542 41972 22594
rect 41916 22482 41972 22542
rect 41916 22430 41918 22482
rect 41970 22430 41972 22482
rect 41916 22418 41972 22430
rect 41916 21474 41972 21486
rect 41916 21422 41918 21474
rect 41970 21422 41972 21474
rect 41916 21252 41972 21422
rect 41916 21186 41972 21196
rect 42028 21364 42084 21374
rect 42028 20802 42084 21308
rect 42028 20750 42030 20802
rect 42082 20750 42084 20802
rect 42028 20738 42084 20750
rect 42252 20356 42308 24556
rect 42364 24546 42420 24556
rect 42924 24164 42980 27580
rect 43148 26964 43204 27002
rect 43148 26898 43204 26908
rect 43148 26290 43204 26302
rect 43148 26238 43150 26290
rect 43202 26238 43204 26290
rect 43036 26180 43092 26190
rect 43036 24722 43092 26124
rect 43148 25956 43204 26238
rect 43148 25890 43204 25900
rect 43036 24670 43038 24722
rect 43090 24670 43092 24722
rect 43036 24658 43092 24670
rect 43148 25618 43204 25630
rect 43148 25566 43150 25618
rect 43202 25566 43204 25618
rect 42812 24108 42980 24164
rect 42476 23828 42532 23838
rect 42700 23828 42756 23838
rect 42476 23734 42532 23772
rect 42588 23826 42756 23828
rect 42588 23774 42702 23826
rect 42754 23774 42756 23826
rect 42588 23772 42756 23774
rect 42588 23156 42644 23772
rect 42700 23762 42756 23772
rect 42588 23062 42644 23100
rect 42812 22482 42868 24108
rect 42924 23940 42980 23950
rect 42924 23846 42980 23884
rect 43148 23938 43204 25566
rect 43260 25284 43316 25294
rect 43260 24722 43316 25228
rect 43260 24670 43262 24722
rect 43314 24670 43316 24722
rect 43260 24658 43316 24670
rect 43148 23886 43150 23938
rect 43202 23886 43204 23938
rect 43148 23156 43204 23886
rect 43260 23156 43316 23166
rect 43148 23154 43316 23156
rect 43148 23102 43262 23154
rect 43314 23102 43316 23154
rect 43148 23100 43316 23102
rect 43260 23090 43316 23100
rect 42812 22430 42814 22482
rect 42866 22430 42868 22482
rect 42364 22148 42420 22158
rect 42364 22054 42420 22092
rect 42812 21812 42868 22430
rect 43260 22484 43316 22494
rect 43372 22484 43428 29148
rect 43484 29202 43540 29214
rect 44044 29204 44100 29260
rect 44492 29204 44548 32620
rect 43484 29150 43486 29202
rect 43538 29150 43540 29202
rect 43484 28642 43540 29150
rect 43820 29148 44100 29204
rect 44268 29148 44548 29204
rect 43820 28756 43876 29148
rect 43484 28590 43486 28642
rect 43538 28590 43540 28642
rect 43484 28578 43540 28590
rect 43596 28700 43876 28756
rect 43932 28980 43988 28990
rect 43932 28754 43988 28924
rect 43932 28702 43934 28754
rect 43986 28702 43988 28754
rect 43596 28084 43652 28700
rect 43932 28690 43988 28702
rect 43708 28532 43764 28542
rect 43708 28438 43764 28476
rect 44044 28530 44100 28542
rect 44044 28478 44046 28530
rect 44098 28478 44100 28530
rect 43596 28018 43652 28028
rect 44044 28420 44100 28478
rect 44044 27860 44100 28364
rect 44156 27860 44212 27870
rect 44044 27858 44212 27860
rect 44044 27806 44158 27858
rect 44210 27806 44212 27858
rect 44044 27804 44212 27806
rect 44156 27794 44212 27804
rect 43596 27636 43652 27646
rect 43596 27186 43652 27580
rect 43596 27134 43598 27186
rect 43650 27134 43652 27186
rect 43596 27122 43652 27134
rect 44044 26964 44100 27002
rect 44044 26898 44100 26908
rect 44268 26964 44324 29148
rect 44604 29092 44660 38612
rect 45724 37828 45780 37838
rect 45724 37734 45780 37772
rect 45052 37380 45108 37390
rect 45052 37286 45108 37324
rect 45052 36596 45108 36606
rect 44940 35812 44996 35822
rect 44940 35718 44996 35756
rect 44940 34692 44996 34702
rect 44940 34354 44996 34636
rect 44940 34302 44942 34354
rect 44994 34302 44996 34354
rect 44940 34290 44996 34302
rect 44828 33012 44884 33022
rect 44828 32674 44884 32956
rect 44828 32622 44830 32674
rect 44882 32622 44884 32674
rect 44828 32610 44884 32622
rect 44940 32674 44996 32686
rect 44940 32622 44942 32674
rect 44994 32622 44996 32674
rect 44940 32452 44996 32622
rect 44828 32004 44884 32014
rect 44940 32004 44996 32396
rect 44884 31948 44996 32004
rect 44716 31668 44772 31678
rect 44716 31574 44772 31612
rect 44716 31220 44772 31230
rect 44828 31220 44884 31948
rect 44716 31218 44884 31220
rect 44716 31166 44718 31218
rect 44770 31166 44884 31218
rect 44716 31164 44884 31166
rect 44716 31154 44772 31164
rect 44268 26898 44324 26908
rect 44380 29036 44660 29092
rect 43708 26516 43764 26526
rect 43708 26422 43764 26460
rect 43596 26404 43652 26414
rect 43596 26310 43652 26348
rect 43820 26292 43876 26302
rect 43708 26290 44100 26292
rect 43708 26238 43822 26290
rect 43874 26238 44100 26290
rect 43708 26236 44100 26238
rect 43484 23156 43540 23166
rect 43484 23062 43540 23100
rect 43260 22482 43428 22484
rect 43260 22430 43262 22482
rect 43314 22430 43428 22482
rect 43260 22428 43428 22430
rect 43260 22418 43316 22428
rect 43372 21812 43428 22428
rect 42812 21746 42868 21756
rect 43036 21810 43428 21812
rect 43036 21758 43374 21810
rect 43426 21758 43428 21810
rect 43036 21756 43428 21758
rect 42588 21474 42644 21486
rect 42588 21422 42590 21474
rect 42642 21422 42644 21474
rect 42588 21252 42644 21422
rect 42364 20804 42420 20814
rect 42364 20710 42420 20748
rect 42588 20802 42644 21196
rect 42588 20750 42590 20802
rect 42642 20750 42644 20802
rect 42588 20738 42644 20750
rect 43036 20914 43092 21756
rect 43372 21746 43428 21756
rect 43484 21698 43540 21710
rect 43484 21646 43486 21698
rect 43538 21646 43540 21698
rect 43148 21586 43204 21598
rect 43148 21534 43150 21586
rect 43202 21534 43204 21586
rect 43148 21252 43204 21534
rect 43484 21364 43540 21646
rect 43484 21298 43540 21308
rect 43148 21186 43204 21196
rect 43708 21140 43764 26236
rect 43820 26226 43876 26236
rect 43820 26068 43876 26078
rect 43820 25730 43876 26012
rect 44044 26066 44100 26236
rect 44044 26014 44046 26066
rect 44098 26014 44100 26066
rect 44044 26002 44100 26014
rect 44268 26178 44324 26190
rect 44268 26126 44270 26178
rect 44322 26126 44324 26178
rect 44268 25956 44324 26126
rect 44268 25890 44324 25900
rect 43820 25678 43822 25730
rect 43874 25678 43876 25730
rect 43820 25666 43876 25678
rect 43932 25508 43988 25518
rect 44380 25508 44436 29036
rect 44716 28644 44772 28654
rect 44604 28418 44660 28430
rect 44604 28366 44606 28418
rect 44658 28366 44660 28418
rect 44604 28196 44660 28366
rect 44604 28130 44660 28140
rect 44492 27188 44548 27198
rect 44492 26850 44548 27132
rect 44492 26798 44494 26850
rect 44546 26798 44548 26850
rect 44492 26786 44548 26798
rect 44716 26178 44772 28588
rect 44716 26126 44718 26178
rect 44770 26126 44772 26178
rect 44716 26066 44772 26126
rect 44716 26014 44718 26066
rect 44770 26014 44772 26066
rect 44716 26002 44772 26014
rect 44940 27746 44996 27758
rect 44940 27694 44942 27746
rect 44994 27694 44996 27746
rect 43932 25414 43988 25452
rect 44268 25452 44436 25508
rect 44044 25284 44100 25294
rect 44044 25190 44100 25228
rect 43932 24612 43988 24622
rect 43932 24610 44212 24612
rect 43932 24558 43934 24610
rect 43986 24558 44212 24610
rect 43932 24556 44212 24558
rect 43932 24546 43988 24556
rect 44156 24498 44212 24556
rect 44156 24446 44158 24498
rect 44210 24446 44212 24498
rect 44156 24434 44212 24446
rect 43932 24052 43988 24062
rect 43820 23492 43876 23502
rect 43820 21586 43876 23436
rect 43932 22482 43988 23996
rect 43932 22430 43934 22482
rect 43986 22430 43988 22482
rect 43932 22418 43988 22430
rect 44156 23042 44212 23054
rect 44156 22990 44158 23042
rect 44210 22990 44212 23042
rect 44156 21812 44212 22990
rect 44156 21746 44212 21756
rect 43820 21534 43822 21586
rect 43874 21534 43876 21586
rect 43820 21522 43876 21534
rect 43932 21476 43988 21486
rect 43932 21382 43988 21420
rect 43708 21074 43764 21084
rect 43036 20862 43038 20914
rect 43090 20862 43092 20914
rect 43036 20804 43092 20862
rect 42476 20578 42532 20590
rect 42476 20526 42478 20578
rect 42530 20526 42532 20578
rect 42252 20300 42420 20356
rect 42252 20018 42308 20030
rect 42252 19966 42254 20018
rect 42306 19966 42308 20018
rect 41804 19236 41860 19246
rect 42252 19236 42308 19966
rect 41804 19234 42308 19236
rect 41804 19182 41806 19234
rect 41858 19182 42308 19234
rect 41804 19180 42308 19182
rect 41804 19170 41860 19180
rect 41580 19122 41748 19124
rect 41580 19070 41582 19122
rect 41634 19070 41748 19122
rect 41580 19068 41748 19070
rect 41580 18900 41636 19068
rect 41580 18834 41636 18844
rect 41580 18676 41636 18686
rect 41580 18562 41636 18620
rect 42252 18676 42308 19180
rect 42252 18610 42308 18620
rect 41580 18510 41582 18562
rect 41634 18510 41636 18562
rect 41580 18498 41636 18510
rect 41804 18228 41860 18238
rect 42140 18228 42196 18238
rect 42364 18228 42420 20300
rect 42476 19906 42532 20526
rect 42476 19854 42478 19906
rect 42530 19854 42532 19906
rect 42476 19842 42532 19854
rect 42588 20020 42644 20030
rect 42588 19236 42644 19964
rect 42924 19906 42980 19918
rect 42924 19854 42926 19906
rect 42978 19854 42980 19906
rect 42924 19346 42980 19854
rect 42924 19294 42926 19346
rect 42978 19294 42980 19346
rect 42924 19236 42980 19294
rect 42588 19234 42868 19236
rect 42588 19182 42590 19234
rect 42642 19182 42868 19234
rect 42588 19180 42868 19182
rect 42588 19170 42644 19180
rect 42812 19124 42868 19180
rect 42924 19170 42980 19180
rect 42812 18676 42868 19068
rect 42924 18676 42980 18686
rect 42812 18674 42980 18676
rect 42812 18622 42926 18674
rect 42978 18622 42980 18674
rect 42812 18620 42980 18622
rect 42924 18610 42980 18620
rect 43036 18452 43092 20748
rect 44044 19236 44100 19246
rect 44044 19142 44100 19180
rect 43484 19122 43540 19134
rect 43484 19070 43486 19122
rect 43538 19070 43540 19122
rect 43484 18674 43540 19070
rect 44156 19124 44212 19134
rect 44156 19030 44212 19068
rect 44268 18788 44324 25452
rect 44940 25396 44996 27694
rect 44940 25330 44996 25340
rect 44380 25284 44436 25294
rect 44380 24946 44436 25228
rect 44604 25284 44660 25294
rect 44604 25190 44660 25228
rect 45052 25172 45108 36540
rect 45500 36260 45556 36270
rect 45500 36258 45668 36260
rect 45500 36206 45502 36258
rect 45554 36206 45668 36258
rect 45500 36204 45668 36206
rect 45500 36194 45556 36204
rect 45500 35924 45556 35934
rect 45500 35830 45556 35868
rect 45388 35812 45444 35822
rect 45388 35476 45444 35756
rect 45612 35700 45668 36204
rect 45948 35812 46004 39340
rect 46060 39330 46116 39340
rect 46508 39396 46564 39406
rect 45948 35746 46004 35756
rect 46060 38724 46116 38734
rect 45724 35700 45780 35710
rect 45612 35698 45892 35700
rect 45612 35646 45726 35698
rect 45778 35646 45892 35698
rect 45612 35644 45892 35646
rect 45724 35634 45780 35644
rect 45836 35588 45892 35644
rect 45948 35588 46004 35598
rect 45836 35532 45948 35588
rect 45724 35476 45780 35486
rect 45388 35420 45668 35476
rect 45612 35026 45668 35420
rect 45612 34974 45614 35026
rect 45666 34974 45668 35026
rect 45612 34962 45668 34974
rect 45500 33908 45556 33918
rect 45500 33458 45556 33852
rect 45500 33406 45502 33458
rect 45554 33406 45556 33458
rect 45500 33394 45556 33406
rect 45164 32564 45220 32574
rect 45164 32562 45332 32564
rect 45164 32510 45166 32562
rect 45218 32510 45332 32562
rect 45164 32508 45332 32510
rect 45164 32498 45220 32508
rect 45164 32340 45220 32350
rect 45164 31556 45220 32284
rect 45276 31780 45332 32508
rect 45500 32452 45556 32462
rect 45500 32358 45556 32396
rect 45724 32004 45780 35420
rect 45836 34914 45892 35532
rect 45948 35522 46004 35532
rect 45836 34862 45838 34914
rect 45890 34862 45892 34914
rect 45836 34468 45892 34862
rect 45836 34402 45892 34412
rect 46060 34356 46116 38668
rect 46284 38724 46340 38734
rect 46508 38724 46564 39340
rect 46732 39058 46788 39564
rect 46732 39006 46734 39058
rect 46786 39006 46788 39058
rect 46732 38994 46788 39006
rect 46956 40404 47012 40414
rect 46340 38668 46564 38724
rect 46732 38836 46788 38846
rect 46284 38630 46340 38668
rect 46172 38612 46228 38622
rect 46172 35812 46228 38556
rect 46732 38162 46788 38780
rect 46732 38110 46734 38162
rect 46786 38110 46788 38162
rect 46732 38098 46788 38110
rect 46284 37828 46340 37838
rect 46620 37828 46676 37838
rect 46284 37044 46340 37772
rect 46508 37826 46676 37828
rect 46508 37774 46622 37826
rect 46674 37774 46676 37826
rect 46508 37772 46676 37774
rect 46284 36706 46340 36988
rect 46284 36654 46286 36706
rect 46338 36654 46340 36706
rect 46284 36642 46340 36654
rect 46396 37266 46452 37278
rect 46396 37214 46398 37266
rect 46450 37214 46452 37266
rect 46396 36260 46452 37214
rect 46508 36594 46564 37772
rect 46620 37762 46676 37772
rect 46844 37826 46900 37838
rect 46844 37774 46846 37826
rect 46898 37774 46900 37826
rect 46844 37380 46900 37774
rect 46844 37266 46900 37324
rect 46844 37214 46846 37266
rect 46898 37214 46900 37266
rect 46844 37202 46900 37214
rect 46508 36542 46510 36594
rect 46562 36542 46564 36594
rect 46508 36530 46564 36542
rect 46732 37044 46788 37054
rect 46508 36260 46564 36270
rect 46396 36258 46564 36260
rect 46396 36206 46510 36258
rect 46562 36206 46564 36258
rect 46396 36204 46564 36206
rect 46508 35924 46564 36204
rect 46508 35858 46564 35868
rect 46620 36148 46676 36158
rect 46172 35756 46452 35812
rect 46172 35588 46228 35626
rect 46172 35522 46228 35532
rect 45612 31948 45780 32004
rect 45948 34300 46116 34356
rect 45388 31780 45444 31790
rect 45276 31778 45444 31780
rect 45276 31726 45390 31778
rect 45442 31726 45444 31778
rect 45276 31724 45444 31726
rect 45388 31714 45444 31724
rect 45164 31500 45556 31556
rect 45388 30660 45444 30670
rect 45164 29764 45220 29774
rect 45164 29650 45220 29708
rect 45164 29598 45166 29650
rect 45218 29598 45220 29650
rect 45164 29586 45220 29598
rect 45388 28756 45444 30604
rect 45388 28624 45444 28700
rect 45500 28196 45556 31500
rect 45612 30100 45668 31948
rect 45948 31892 46004 34300
rect 46060 34130 46116 34142
rect 46060 34078 46062 34130
rect 46114 34078 46116 34130
rect 46060 33908 46116 34078
rect 46060 33124 46116 33852
rect 46396 33572 46452 35756
rect 46060 33058 46116 33068
rect 46284 33516 46452 33572
rect 46508 34802 46564 34814
rect 46508 34750 46510 34802
rect 46562 34750 46564 34802
rect 46508 34018 46564 34750
rect 46508 33966 46510 34018
rect 46562 33966 46564 34018
rect 45612 30034 45668 30044
rect 45724 31836 46004 31892
rect 45724 29540 45780 31836
rect 46060 31780 46116 31790
rect 45836 31668 45892 31678
rect 45836 30994 45892 31612
rect 45948 31556 46004 31566
rect 45948 31462 46004 31500
rect 45836 30942 45838 30994
rect 45890 30942 45892 30994
rect 45836 30930 45892 30942
rect 46060 30882 46116 31724
rect 46060 30830 46062 30882
rect 46114 30830 46116 30882
rect 46060 30818 46116 30830
rect 46060 29988 46116 29998
rect 45724 29484 45892 29540
rect 45388 28140 45556 28196
rect 45724 29316 45780 29326
rect 45388 26908 45444 28140
rect 45612 27972 45668 27982
rect 45612 27878 45668 27916
rect 45500 27860 45556 27870
rect 45500 27300 45556 27804
rect 45612 27300 45668 27310
rect 45500 27244 45612 27300
rect 45612 27168 45668 27244
rect 45724 26908 45780 29260
rect 45836 28754 45892 29484
rect 46060 29204 46116 29932
rect 46284 29876 46340 33516
rect 46396 33348 46452 33358
rect 46508 33348 46564 33966
rect 46396 33346 46564 33348
rect 46396 33294 46398 33346
rect 46450 33294 46564 33346
rect 46396 33292 46564 33294
rect 46396 33282 46452 33292
rect 46508 33124 46564 33134
rect 46508 33030 46564 33068
rect 46396 30772 46452 30782
rect 46396 30678 46452 30716
rect 46620 30660 46676 36092
rect 46732 35922 46788 36988
rect 46732 35870 46734 35922
rect 46786 35870 46788 35922
rect 46732 35858 46788 35870
rect 46956 35140 47012 40348
rect 47068 40178 47124 40190
rect 47068 40126 47070 40178
rect 47122 40126 47124 40178
rect 47068 39506 47124 40126
rect 47068 39454 47070 39506
rect 47122 39454 47124 39506
rect 47068 39396 47124 39454
rect 47068 39330 47124 39340
rect 47180 39058 47236 40460
rect 47852 40404 47908 40908
rect 48300 40514 48356 40526
rect 48300 40462 48302 40514
rect 48354 40462 48356 40514
rect 47404 40178 47460 40190
rect 47404 40126 47406 40178
rect 47458 40126 47460 40178
rect 47292 39620 47348 39630
rect 47292 39526 47348 39564
rect 47180 39006 47182 39058
rect 47234 39006 47236 39058
rect 47180 38994 47236 39006
rect 47404 38668 47460 40126
rect 47404 38612 47684 38668
rect 47068 37826 47124 37838
rect 47068 37774 47070 37826
rect 47122 37774 47124 37826
rect 47068 36482 47124 37774
rect 47516 37268 47572 37278
rect 47068 36430 47070 36482
rect 47122 36430 47124 36482
rect 47068 36418 47124 36430
rect 47404 37266 47572 37268
rect 47404 37214 47518 37266
rect 47570 37214 47572 37266
rect 47404 37212 47572 37214
rect 47404 37044 47460 37212
rect 47516 37202 47572 37212
rect 47404 36482 47460 36988
rect 47404 36430 47406 36482
rect 47458 36430 47460 36482
rect 47404 36418 47460 36430
rect 47292 36258 47348 36270
rect 47292 36206 47294 36258
rect 47346 36206 47348 36258
rect 47180 36036 47236 36046
rect 46956 35084 47124 35140
rect 46956 34916 47012 34926
rect 46732 34914 47012 34916
rect 46732 34862 46958 34914
rect 47010 34862 47012 34914
rect 46732 34860 47012 34862
rect 46732 33346 46788 34860
rect 46956 34850 47012 34860
rect 47068 34692 47124 35084
rect 46732 33294 46734 33346
rect 46786 33294 46788 33346
rect 46732 33282 46788 33294
rect 46844 34636 47124 34692
rect 46620 30594 46676 30604
rect 46396 30212 46452 30222
rect 46844 30212 46900 34636
rect 46956 34244 47012 34254
rect 46956 34150 47012 34188
rect 47068 33124 47124 33134
rect 47068 33030 47124 33068
rect 47068 31892 47124 31902
rect 47180 31892 47236 35980
rect 47292 35924 47348 36206
rect 47292 35858 47348 35868
rect 47516 35252 47572 35262
rect 47516 35026 47572 35196
rect 47516 34974 47518 35026
rect 47570 34974 47572 35026
rect 47516 34962 47572 34974
rect 47628 35028 47684 38612
rect 47852 37268 47908 40348
rect 48188 40402 48244 40414
rect 48188 40350 48190 40402
rect 48242 40350 48244 40402
rect 48188 39844 48244 40350
rect 47964 39788 48244 39844
rect 47964 39508 48020 39788
rect 47964 38722 48020 39452
rect 48076 38836 48132 38846
rect 48300 38836 48356 40462
rect 48524 40516 48580 40526
rect 48524 40422 48580 40460
rect 48636 39396 48692 39406
rect 48636 39302 48692 39340
rect 48132 38780 48356 38836
rect 48076 38742 48132 38780
rect 47964 38670 47966 38722
rect 48018 38670 48020 38722
rect 47964 38658 48020 38670
rect 48748 38724 48804 38734
rect 48748 38630 48804 38668
rect 47852 37212 48020 37268
rect 47852 37044 47908 37054
rect 47852 36594 47908 36988
rect 47852 36542 47854 36594
rect 47906 36542 47908 36594
rect 47852 36530 47908 36542
rect 47740 35588 47796 35598
rect 47740 35494 47796 35532
rect 47628 34962 47684 34972
rect 47740 35364 47796 35374
rect 47404 34690 47460 34702
rect 47404 34638 47406 34690
rect 47458 34638 47460 34690
rect 47404 34244 47460 34638
rect 47404 34178 47460 34188
rect 47628 34690 47684 34702
rect 47628 34638 47630 34690
rect 47682 34638 47684 34690
rect 47628 34020 47684 34638
rect 47628 33926 47684 33964
rect 47068 31890 47236 31892
rect 47068 31838 47070 31890
rect 47122 31838 47236 31890
rect 47068 31836 47236 31838
rect 47068 31826 47124 31836
rect 47180 31780 47236 31836
rect 47180 31714 47236 31724
rect 47516 31554 47572 31566
rect 47516 31502 47518 31554
rect 47570 31502 47572 31554
rect 47516 31332 47572 31502
rect 47180 31276 47572 31332
rect 47180 31218 47236 31276
rect 47180 31166 47182 31218
rect 47234 31166 47236 31218
rect 47180 31154 47236 31166
rect 47404 31108 47460 31118
rect 47404 30322 47460 31052
rect 47404 30270 47406 30322
rect 47458 30270 47460 30322
rect 47404 30258 47460 30270
rect 46396 30210 46900 30212
rect 46396 30158 46398 30210
rect 46450 30158 46846 30210
rect 46898 30158 46900 30210
rect 46396 30156 46900 30158
rect 46396 30146 46452 30156
rect 46284 29810 46340 29820
rect 46396 29764 46452 29774
rect 46284 29652 46340 29662
rect 46284 29558 46340 29596
rect 46396 29650 46452 29708
rect 46396 29598 46398 29650
rect 46450 29598 46452 29650
rect 46060 29138 46116 29148
rect 46172 29316 46228 29326
rect 45836 28702 45838 28754
rect 45890 28702 45892 28754
rect 45836 28196 45892 28702
rect 45836 28130 45892 28140
rect 45948 28756 46004 28766
rect 46172 28756 46228 29260
rect 46284 28756 46340 28766
rect 46172 28700 46284 28756
rect 45948 27860 46004 28700
rect 46284 28624 46340 28700
rect 46396 28420 46452 29598
rect 45948 27794 46004 27804
rect 46060 28364 46452 28420
rect 46620 28644 46676 28654
rect 45948 27634 46004 27646
rect 45948 27582 45950 27634
rect 46002 27582 46004 27634
rect 45836 27074 45892 27086
rect 45836 27022 45838 27074
rect 45890 27022 45892 27074
rect 45836 26908 45892 27022
rect 45388 26852 45556 26908
rect 45724 26852 45892 26908
rect 44380 24894 44382 24946
rect 44434 24894 44436 24946
rect 44380 24882 44436 24894
rect 44940 25116 45108 25172
rect 45388 26628 45444 26638
rect 45388 26514 45444 26572
rect 45388 26462 45390 26514
rect 45442 26462 45444 26514
rect 44828 24498 44884 24510
rect 44828 24446 44830 24498
rect 44882 24446 44884 24498
rect 44380 24052 44436 24062
rect 44380 22148 44436 23996
rect 44828 23156 44884 24446
rect 44940 23268 44996 25116
rect 45052 24948 45108 24958
rect 45388 24948 45444 26462
rect 45500 26404 45556 26852
rect 45500 26338 45556 26348
rect 45612 26292 45668 26302
rect 45612 26198 45668 26236
rect 45500 26178 45556 26190
rect 45500 26126 45502 26178
rect 45554 26126 45556 26178
rect 45500 25620 45556 26126
rect 45836 26066 45892 26852
rect 45948 26852 46004 27582
rect 46060 27412 46116 28364
rect 46060 27074 46116 27356
rect 46508 28196 46564 28206
rect 46508 27858 46564 28140
rect 46508 27806 46510 27858
rect 46562 27806 46564 27858
rect 46172 27188 46228 27198
rect 46172 27094 46228 27132
rect 46060 27022 46062 27074
rect 46114 27022 46116 27074
rect 46060 26908 46116 27022
rect 46508 26964 46564 27806
rect 46060 26852 46228 26908
rect 45948 26786 46004 26796
rect 46060 26404 46116 26414
rect 46060 26310 46116 26348
rect 45836 26014 45838 26066
rect 45890 26014 45892 26066
rect 45836 26002 45892 26014
rect 45948 26292 46004 26302
rect 45500 25564 45780 25620
rect 45052 24946 45444 24948
rect 45052 24894 45054 24946
rect 45106 24894 45444 24946
rect 45052 24892 45444 24894
rect 45500 25396 45556 25406
rect 45052 24882 45108 24892
rect 45388 24724 45444 24734
rect 44940 23202 44996 23212
rect 45052 24052 45108 24062
rect 44492 23154 44884 23156
rect 44492 23102 44830 23154
rect 44882 23102 44884 23154
rect 44492 23100 44884 23102
rect 44492 22370 44548 23100
rect 44828 23090 44884 23100
rect 45052 23154 45108 23996
rect 45052 23102 45054 23154
rect 45106 23102 45108 23154
rect 45052 23090 45108 23102
rect 45388 22932 45444 24668
rect 45500 24052 45556 25340
rect 45612 25284 45668 25294
rect 45612 25190 45668 25228
rect 45612 24052 45668 24062
rect 45500 24050 45668 24052
rect 45500 23998 45614 24050
rect 45666 23998 45668 24050
rect 45500 23996 45668 23998
rect 45612 23986 45668 23996
rect 45724 23492 45780 25564
rect 45836 25506 45892 25518
rect 45836 25454 45838 25506
rect 45890 25454 45892 25506
rect 45836 23940 45892 25454
rect 45836 23846 45892 23884
rect 45948 23492 46004 26236
rect 46060 24500 46116 24510
rect 46060 24406 46116 24444
rect 45724 23426 45780 23436
rect 45836 23436 46004 23492
rect 45388 22866 45444 22876
rect 45612 23044 45668 23054
rect 44492 22318 44494 22370
rect 44546 22318 44548 22370
rect 44492 22306 44548 22318
rect 44828 22372 44884 22382
rect 44828 22278 44884 22316
rect 45500 22372 45556 22382
rect 45500 22278 45556 22316
rect 44604 22148 44660 22158
rect 44380 22146 44660 22148
rect 44380 22094 44606 22146
rect 44658 22094 44660 22146
rect 44380 22092 44660 22094
rect 44604 22082 44660 22092
rect 45052 21700 45108 21710
rect 45052 21606 45108 21644
rect 44492 21474 44548 21486
rect 44492 21422 44494 21474
rect 44546 21422 44548 21474
rect 44492 21364 44548 21422
rect 44716 21476 44772 21486
rect 44716 21382 44772 21420
rect 44492 21298 44548 21308
rect 45612 20916 45668 22988
rect 45724 23042 45780 23054
rect 45724 22990 45726 23042
rect 45778 22990 45780 23042
rect 45724 22260 45780 22990
rect 45724 21586 45780 22204
rect 45724 21534 45726 21586
rect 45778 21534 45780 21586
rect 45724 21522 45780 21534
rect 45836 21028 45892 23436
rect 46060 22372 46116 22382
rect 46172 22372 46228 26852
rect 46284 26852 46564 26908
rect 46284 26850 46340 26852
rect 46284 26798 46286 26850
rect 46338 26798 46340 26850
rect 46284 26786 46340 26798
rect 46620 26628 46676 28588
rect 46508 26178 46564 26190
rect 46508 26126 46510 26178
rect 46562 26126 46564 26178
rect 46508 26066 46564 26126
rect 46508 26014 46510 26066
rect 46562 26014 46564 26066
rect 46508 26002 46564 26014
rect 46620 25396 46676 26572
rect 46732 27972 46788 27982
rect 46732 26292 46788 27916
rect 46732 26226 46788 26236
rect 46844 25508 46900 30156
rect 47516 30212 47572 31276
rect 47628 31220 47684 31230
rect 47740 31220 47796 35308
rect 47852 34244 47908 34254
rect 47852 34130 47908 34188
rect 47852 34078 47854 34130
rect 47906 34078 47908 34130
rect 47852 34066 47908 34078
rect 47628 31218 47740 31220
rect 47628 31166 47630 31218
rect 47682 31166 47740 31218
rect 47628 31164 47740 31166
rect 47628 31154 47684 31164
rect 47740 31088 47796 31164
rect 47516 30146 47572 30156
rect 47292 29988 47348 29998
rect 47292 29894 47348 29932
rect 47516 29986 47572 29998
rect 47516 29934 47518 29986
rect 47570 29934 47572 29986
rect 46956 29876 47012 29886
rect 46956 29652 47012 29820
rect 47516 29652 47572 29934
rect 46956 29650 47236 29652
rect 46956 29598 46958 29650
rect 47010 29598 47236 29650
rect 46956 29596 47236 29598
rect 46956 29586 47012 29596
rect 47068 28756 47124 28766
rect 47068 28662 47124 28700
rect 47180 28644 47236 29596
rect 47516 29586 47572 29596
rect 47740 29988 47796 29998
rect 47740 29650 47796 29932
rect 47740 29598 47742 29650
rect 47794 29598 47796 29650
rect 47740 29586 47796 29598
rect 47180 28512 47236 28588
rect 47404 27972 47460 27982
rect 47404 27878 47460 27916
rect 47964 27972 48020 37212
rect 48300 37154 48356 37166
rect 48300 37102 48302 37154
rect 48354 37102 48356 37154
rect 48300 35700 48356 37102
rect 48300 35634 48356 35644
rect 48188 35586 48244 35598
rect 48188 35534 48190 35586
rect 48242 35534 48244 35586
rect 48188 35028 48244 35534
rect 49084 35140 49140 35150
rect 48188 34962 48244 34972
rect 48972 35028 49028 35038
rect 48972 34802 49028 34972
rect 48972 34750 48974 34802
rect 49026 34750 49028 34802
rect 48972 34132 49028 34750
rect 48972 34066 49028 34076
rect 49084 34914 49140 35084
rect 49084 34862 49086 34914
rect 49138 34862 49140 34914
rect 48524 34018 48580 34030
rect 48524 33966 48526 34018
rect 48578 33966 48580 34018
rect 48300 31890 48356 31902
rect 48300 31838 48302 31890
rect 48354 31838 48356 31890
rect 48188 31220 48244 31230
rect 48188 31106 48244 31164
rect 48188 31054 48190 31106
rect 48242 31054 48244 31106
rect 48188 30660 48244 31054
rect 48300 30772 48356 31838
rect 48524 31892 48580 33966
rect 48972 33570 49028 33582
rect 48972 33518 48974 33570
rect 49026 33518 49028 33570
rect 48972 33124 49028 33518
rect 48524 31826 48580 31836
rect 48636 33122 49028 33124
rect 48636 33070 48974 33122
rect 49026 33070 49028 33122
rect 48636 33068 49028 33070
rect 48412 31780 48468 31790
rect 48412 31220 48468 31724
rect 48412 31154 48468 31164
rect 48412 30772 48468 30782
rect 48300 30770 48580 30772
rect 48300 30718 48414 30770
rect 48466 30718 48580 30770
rect 48300 30716 48580 30718
rect 48412 30706 48468 30716
rect 48188 30594 48244 30604
rect 48412 30324 48468 30334
rect 48412 30230 48468 30268
rect 48524 30212 48580 30716
rect 48524 30146 48580 30156
rect 48076 30098 48132 30110
rect 48076 30046 48078 30098
rect 48130 30046 48132 30098
rect 48076 29652 48132 30046
rect 48300 29988 48356 29998
rect 48300 29894 48356 29932
rect 48076 29586 48132 29596
rect 48076 28868 48132 28878
rect 48636 28868 48692 33068
rect 48972 33058 49028 33068
rect 49084 32900 49140 34862
rect 48860 32844 49140 32900
rect 48748 31220 48804 31230
rect 48860 31220 48916 32844
rect 49196 32788 49252 40908
rect 49196 32722 49252 32732
rect 49308 39396 49364 41132
rect 49420 41094 49476 41132
rect 49084 31668 49140 31678
rect 49084 31574 49140 31612
rect 49308 31556 49364 39340
rect 49532 40404 49588 42476
rect 49756 42530 49812 42542
rect 49756 42478 49758 42530
rect 49810 42478 49812 42530
rect 49756 41860 49812 42478
rect 50092 41970 50148 41982
rect 50092 41918 50094 41970
rect 50146 41918 50148 41970
rect 49980 41860 50036 41870
rect 49812 41858 50036 41860
rect 49812 41806 49982 41858
rect 50034 41806 50036 41858
rect 49812 41804 50036 41806
rect 49756 41728 49812 41804
rect 49980 41412 50036 41804
rect 50092 41412 50148 41918
rect 50204 41412 50260 41422
rect 50092 41410 50260 41412
rect 50092 41358 50206 41410
rect 50258 41358 50260 41410
rect 50092 41356 50260 41358
rect 49980 41346 50036 41356
rect 50204 41346 50260 41356
rect 50092 41074 50148 41086
rect 50092 41022 50094 41074
rect 50146 41022 50148 41074
rect 50092 40740 50148 41022
rect 50204 40964 50260 40974
rect 50204 40870 50260 40908
rect 49756 40684 50148 40740
rect 49756 40404 49812 40684
rect 50316 40516 50372 43652
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 50764 40964 50820 41002
rect 50764 40898 50820 40908
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 50204 40460 50372 40516
rect 50764 40516 50820 40526
rect 49980 40404 50036 40414
rect 49532 40402 49812 40404
rect 49532 40350 49534 40402
rect 49586 40350 49812 40402
rect 49532 40348 49812 40350
rect 49868 40402 50036 40404
rect 49868 40350 49982 40402
rect 50034 40350 50036 40402
rect 49868 40348 50036 40350
rect 49532 38668 49588 40348
rect 49868 39396 49924 40348
rect 49980 40338 50036 40348
rect 49868 39330 49924 39340
rect 49980 39506 50036 39518
rect 49980 39454 49982 39506
rect 50034 39454 50036 39506
rect 49868 38948 49924 38958
rect 49868 38834 49924 38892
rect 49868 38782 49870 38834
rect 49922 38782 49924 38834
rect 49868 38770 49924 38782
rect 49420 38612 49588 38668
rect 49980 38724 50036 39454
rect 50092 39394 50148 39406
rect 50092 39342 50094 39394
rect 50146 39342 50148 39394
rect 50092 38836 50148 39342
rect 50092 38770 50148 38780
rect 49980 38658 50036 38668
rect 49420 35588 49476 38612
rect 50204 36596 50260 40460
rect 50764 40422 50820 40460
rect 50652 40404 50708 40414
rect 50316 40402 50708 40404
rect 50316 40350 50654 40402
rect 50706 40350 50708 40402
rect 50316 40348 50708 40350
rect 50316 39618 50372 40348
rect 50652 40338 50708 40348
rect 50876 39730 50932 44828
rect 51100 44434 51156 44940
rect 51100 44382 51102 44434
rect 51154 44382 51156 44434
rect 51100 44370 51156 44382
rect 51324 44322 51380 45838
rect 51548 45890 51604 45902
rect 51548 45838 51550 45890
rect 51602 45838 51604 45890
rect 51548 44996 51604 45838
rect 51548 44930 51604 44940
rect 51324 44270 51326 44322
rect 51378 44270 51380 44322
rect 51324 43708 51380 44270
rect 50988 43652 51380 43708
rect 50988 40626 51044 43652
rect 51772 42868 51828 48188
rect 51996 48178 52052 48188
rect 52444 48150 52500 48188
rect 52220 48018 52276 48030
rect 52220 47966 52222 48018
rect 52274 47966 52276 48018
rect 52220 47682 52276 47966
rect 52220 47630 52222 47682
rect 52274 47630 52276 47682
rect 52220 47618 52276 47630
rect 51884 47460 51940 47470
rect 51884 47366 51940 47404
rect 52780 46564 52836 50092
rect 53116 50036 53172 50046
rect 53116 49942 53172 49980
rect 53340 48916 53396 48926
rect 53340 48822 53396 48860
rect 53452 48580 53508 50316
rect 53564 50370 53620 50428
rect 53564 50318 53566 50370
rect 53618 50318 53620 50370
rect 53564 50306 53620 50318
rect 53676 50260 53732 50270
rect 53564 49364 53620 49374
rect 53564 48914 53620 49308
rect 53676 49026 53732 50204
rect 53676 48974 53678 49026
rect 53730 48974 53732 49026
rect 53676 48962 53732 48974
rect 53788 49700 53844 49710
rect 53564 48862 53566 48914
rect 53618 48862 53620 48914
rect 53564 48850 53620 48862
rect 53452 48524 53620 48580
rect 53116 48468 53172 48478
rect 53116 48374 53172 48412
rect 53228 46786 53284 46798
rect 53228 46734 53230 46786
rect 53282 46734 53284 46786
rect 53116 46564 53172 46574
rect 52780 46562 53172 46564
rect 52780 46510 53118 46562
rect 53170 46510 53172 46562
rect 52780 46508 53172 46510
rect 53116 46498 53172 46508
rect 52892 45892 52948 45902
rect 51884 45666 51940 45678
rect 51884 45614 51886 45666
rect 51938 45614 51940 45666
rect 51884 45220 51940 45614
rect 51884 45154 51940 45164
rect 52892 45218 52948 45836
rect 53228 45892 53284 46734
rect 53452 46452 53508 46462
rect 53452 46358 53508 46396
rect 53228 45826 53284 45836
rect 53564 45330 53620 48524
rect 53788 47068 53844 49644
rect 53564 45278 53566 45330
rect 53618 45278 53620 45330
rect 53564 45266 53620 45278
rect 53676 47012 53844 47068
rect 52892 45166 52894 45218
rect 52946 45166 52948 45218
rect 52892 45154 52948 45166
rect 51996 45106 52052 45118
rect 51996 45054 51998 45106
rect 52050 45054 52052 45106
rect 51996 44884 52052 45054
rect 51996 44818 52052 44828
rect 52108 45108 52164 45118
rect 52108 44994 52164 45052
rect 53340 45108 53396 45118
rect 53340 45014 53396 45052
rect 52108 44942 52110 44994
rect 52162 44942 52164 44994
rect 51996 44436 52052 44446
rect 52108 44436 52164 44942
rect 51996 44434 52164 44436
rect 51996 44382 51998 44434
rect 52050 44382 52164 44434
rect 51996 44380 52164 44382
rect 51996 44370 52052 44380
rect 51772 42802 51828 42812
rect 52108 44212 52164 44222
rect 51100 41972 51156 41982
rect 51100 41878 51156 41916
rect 51772 41746 51828 41758
rect 51772 41694 51774 41746
rect 51826 41694 51828 41746
rect 50988 40574 50990 40626
rect 51042 40574 51044 40626
rect 50988 40562 51044 40574
rect 51212 41188 51268 41198
rect 51212 40962 51268 41132
rect 51212 40910 51214 40962
rect 51266 40910 51268 40962
rect 50876 39678 50878 39730
rect 50930 39678 50932 39730
rect 50876 39666 50932 39678
rect 50316 39566 50318 39618
rect 50370 39566 50372 39618
rect 50316 39554 50372 39566
rect 50764 39396 50820 39406
rect 50988 39396 51044 39406
rect 50428 39394 50820 39396
rect 50428 39342 50766 39394
rect 50818 39342 50820 39394
rect 50428 39340 50820 39342
rect 50428 38836 50484 39340
rect 50764 39330 50820 39340
rect 50876 39394 51044 39396
rect 50876 39342 50990 39394
rect 51042 39342 51044 39394
rect 50876 39340 51044 39342
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 50876 38948 50932 39340
rect 50988 39330 51044 39340
rect 50316 38834 50484 38836
rect 50316 38782 50430 38834
rect 50482 38782 50484 38834
rect 50316 38780 50484 38782
rect 50316 38274 50372 38780
rect 50428 38770 50484 38780
rect 50540 38836 50596 38846
rect 50540 38742 50596 38780
rect 50316 38222 50318 38274
rect 50370 38222 50372 38274
rect 50316 38210 50372 38222
rect 50764 38164 50820 38174
rect 50764 38070 50820 38108
rect 50428 38052 50484 38062
rect 50428 37958 50484 37996
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 50876 37492 50932 38892
rect 50204 36530 50260 36540
rect 50652 37436 50932 37492
rect 50652 36594 50708 37436
rect 50652 36542 50654 36594
rect 50706 36542 50708 36594
rect 50652 36530 50708 36542
rect 50876 36482 50932 36494
rect 50876 36430 50878 36482
rect 50930 36430 50932 36482
rect 50204 36372 50260 36382
rect 49756 36370 50260 36372
rect 49756 36318 50206 36370
rect 50258 36318 50260 36370
rect 49756 36316 50260 36318
rect 49756 35922 49812 36316
rect 50204 36306 50260 36316
rect 50428 36370 50484 36382
rect 50428 36318 50430 36370
rect 50482 36318 50484 36370
rect 49756 35870 49758 35922
rect 49810 35870 49812 35922
rect 49756 35858 49812 35870
rect 50428 35924 50484 36318
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 50876 35924 50932 36430
rect 51212 36260 51268 40910
rect 51660 40964 51716 40974
rect 51436 39620 51492 39630
rect 51436 39618 51604 39620
rect 51436 39566 51438 39618
rect 51490 39566 51604 39618
rect 51436 39564 51604 39566
rect 51436 39554 51492 39564
rect 51324 38836 51380 38846
rect 51324 38742 51380 38780
rect 51436 38724 51492 38734
rect 51436 38630 51492 38668
rect 51548 38050 51604 39564
rect 51548 37998 51550 38050
rect 51602 37998 51604 38050
rect 51548 37986 51604 37998
rect 51660 37828 51716 40908
rect 51772 39284 51828 41694
rect 52108 41188 52164 44156
rect 53676 43708 53732 47012
rect 53788 45892 53844 45902
rect 53788 45798 53844 45836
rect 53788 45106 53844 45118
rect 53788 45054 53790 45106
rect 53842 45054 53844 45106
rect 53788 44884 53844 45054
rect 53788 44818 53844 44828
rect 53900 44212 53956 50428
rect 54124 50484 54180 50494
rect 54124 50390 54180 50428
rect 54460 49700 54516 50542
rect 55468 50036 55524 51102
rect 54460 49634 54516 49644
rect 55356 49980 55524 50036
rect 54124 49364 54180 49374
rect 54124 49138 54180 49308
rect 55356 49364 55412 49980
rect 55356 49298 55412 49308
rect 55468 49812 55524 49822
rect 55580 49812 55636 51212
rect 55692 51202 55748 51212
rect 55916 50818 55972 51212
rect 56252 51266 56420 51268
rect 56252 51214 56254 51266
rect 56306 51214 56420 51266
rect 56252 51212 56420 51214
rect 56252 51202 56308 51212
rect 55916 50766 55918 50818
rect 55970 50766 55972 50818
rect 55916 50754 55972 50766
rect 56140 50596 56196 50606
rect 55468 49810 55636 49812
rect 55468 49758 55470 49810
rect 55522 49758 55636 49810
rect 55468 49756 55636 49758
rect 55692 50594 56196 50596
rect 55692 50542 56142 50594
rect 56194 50542 56196 50594
rect 55692 50540 56196 50542
rect 55692 49810 55748 50540
rect 55692 49758 55694 49810
rect 55746 49758 55748 49810
rect 55468 49250 55524 49756
rect 55692 49746 55748 49758
rect 55916 49700 55972 49710
rect 55916 49606 55972 49644
rect 55468 49198 55470 49250
rect 55522 49198 55524 49250
rect 55468 49186 55524 49198
rect 55580 49252 55636 49262
rect 54124 49086 54126 49138
rect 54178 49086 54180 49138
rect 54124 49074 54180 49086
rect 55356 48916 55412 48926
rect 55244 48914 55412 48916
rect 55244 48862 55358 48914
rect 55410 48862 55412 48914
rect 55244 48860 55412 48862
rect 54796 48244 54852 48254
rect 54796 48150 54852 48188
rect 54460 47796 54516 47806
rect 54012 46562 54068 46574
rect 54012 46510 54014 46562
rect 54066 46510 54068 46562
rect 54012 46452 54068 46510
rect 54012 45892 54068 46396
rect 54460 46002 54516 47740
rect 54572 47460 54628 47470
rect 54572 47366 54628 47404
rect 55244 47458 55300 48860
rect 55356 48850 55412 48860
rect 55468 48804 55524 48814
rect 55468 48692 55524 48748
rect 55356 48636 55524 48692
rect 55356 48242 55412 48636
rect 55356 48190 55358 48242
rect 55410 48190 55412 48242
rect 55356 48178 55412 48190
rect 55244 47406 55246 47458
rect 55298 47406 55300 47458
rect 55244 47348 55300 47406
rect 55356 47570 55412 47582
rect 55356 47518 55358 47570
rect 55410 47518 55412 47570
rect 55356 47460 55412 47518
rect 55356 47394 55412 47404
rect 55244 47282 55300 47292
rect 55468 46788 55524 46798
rect 55244 46676 55300 46686
rect 55244 46582 55300 46620
rect 55468 46674 55524 46732
rect 55468 46622 55470 46674
rect 55522 46622 55524 46674
rect 55468 46610 55524 46622
rect 55580 46452 55636 49196
rect 55692 48130 55748 48142
rect 55692 48078 55694 48130
rect 55746 48078 55748 48130
rect 55692 47572 55748 48078
rect 55692 47506 55748 47516
rect 55692 47348 55748 47358
rect 55692 46786 55748 47292
rect 56140 47124 56196 50540
rect 56252 50596 56308 50606
rect 56252 50370 56308 50540
rect 56252 50318 56254 50370
rect 56306 50318 56308 50370
rect 56252 50306 56308 50318
rect 56364 50594 56420 51212
rect 56364 50542 56366 50594
rect 56418 50542 56420 50594
rect 56364 49812 56420 50542
rect 56812 50596 56868 50606
rect 56812 50502 56868 50540
rect 56364 49746 56420 49756
rect 56700 49700 56756 49710
rect 56756 49644 56980 49700
rect 56364 49588 56420 49598
rect 56364 49586 56532 49588
rect 56364 49534 56366 49586
rect 56418 49534 56532 49586
rect 56700 49568 56756 49644
rect 56364 49532 56532 49534
rect 56364 49522 56420 49532
rect 56476 49138 56532 49532
rect 56476 49086 56478 49138
rect 56530 49086 56532 49138
rect 56476 49074 56532 49086
rect 56700 49028 56756 49038
rect 56588 48972 56700 49028
rect 56364 47572 56420 47582
rect 56588 47572 56644 48972
rect 56700 48934 56756 48972
rect 56812 48244 56868 48254
rect 56700 48132 56756 48142
rect 56812 48132 56868 48188
rect 56700 48130 56868 48132
rect 56700 48078 56702 48130
rect 56754 48078 56868 48130
rect 56700 48076 56868 48078
rect 56700 48066 56756 48076
rect 56812 47684 56868 48076
rect 56364 47478 56420 47516
rect 56476 47516 56644 47572
rect 56700 47628 56868 47684
rect 56252 47348 56308 47358
rect 56252 47254 56308 47292
rect 56140 47068 56308 47124
rect 55692 46734 55694 46786
rect 55746 46734 55748 46786
rect 55692 46722 55748 46734
rect 55916 46676 55972 46686
rect 55916 46674 56196 46676
rect 55916 46622 55918 46674
rect 55970 46622 56196 46674
rect 55916 46620 56196 46622
rect 55916 46610 55972 46620
rect 55580 46114 55636 46396
rect 56028 46452 56084 46462
rect 56028 46358 56084 46396
rect 55580 46062 55582 46114
rect 55634 46062 55636 46114
rect 55580 46050 55636 46062
rect 55804 46228 55860 46238
rect 54460 45950 54462 46002
rect 54514 45950 54516 46002
rect 54460 45938 54516 45950
rect 54236 45892 54292 45902
rect 54012 45890 54292 45892
rect 54012 45838 54238 45890
rect 54290 45838 54292 45890
rect 54012 45836 54292 45838
rect 54236 45668 54292 45836
rect 54012 45220 54068 45230
rect 54012 45126 54068 45164
rect 53900 44146 53956 44156
rect 53564 43652 53732 43708
rect 53340 42754 53396 42766
rect 53340 42702 53342 42754
rect 53394 42702 53396 42754
rect 52220 42530 52276 42542
rect 52220 42478 52222 42530
rect 52274 42478 52276 42530
rect 52220 41972 52276 42478
rect 53340 42194 53396 42702
rect 53340 42142 53342 42194
rect 53394 42142 53396 42194
rect 53340 42130 53396 42142
rect 53564 42084 53620 43652
rect 54124 43538 54180 43550
rect 54124 43486 54126 43538
rect 54178 43486 54180 43538
rect 53900 42868 53956 42878
rect 53900 42774 53956 42812
rect 54012 42756 54068 42766
rect 54124 42756 54180 43486
rect 54012 42754 54180 42756
rect 54012 42702 54014 42754
rect 54066 42702 54180 42754
rect 54012 42700 54180 42702
rect 54012 42690 54068 42700
rect 53788 42530 53844 42542
rect 53788 42478 53790 42530
rect 53842 42478 53844 42530
rect 53788 42084 53844 42478
rect 53900 42084 53956 42094
rect 53788 42082 53956 42084
rect 53788 42030 53902 42082
rect 53954 42030 53956 42082
rect 53788 42028 53956 42030
rect 52220 41906 52276 41916
rect 52668 41972 52724 41982
rect 52668 41878 52724 41916
rect 53452 41972 53508 41982
rect 52108 41122 52164 41132
rect 52444 41746 52500 41758
rect 52444 41694 52446 41746
rect 52498 41694 52500 41746
rect 52444 41636 52500 41694
rect 51884 40964 51940 40974
rect 51884 40870 51940 40908
rect 52444 40964 52500 41580
rect 53004 41746 53060 41758
rect 53004 41694 53006 41746
rect 53058 41694 53060 41746
rect 53004 41300 53060 41694
rect 53228 41748 53284 41758
rect 53228 41654 53284 41692
rect 53004 41234 53060 41244
rect 53452 41524 53508 41916
rect 53340 41188 53396 41198
rect 52444 40898 52500 40908
rect 52668 40964 52724 40974
rect 52668 40870 52724 40908
rect 53228 40404 53284 40414
rect 51772 39228 51940 39284
rect 51884 38164 51940 39228
rect 52220 38948 52276 38958
rect 52220 38854 52276 38892
rect 51772 38052 51828 38062
rect 51772 37938 51828 37996
rect 51884 38050 51940 38108
rect 51884 37998 51886 38050
rect 51938 37998 51940 38050
rect 51884 37986 51940 37998
rect 51772 37886 51774 37938
rect 51826 37886 51828 37938
rect 51772 37874 51828 37886
rect 50428 35858 50484 35868
rect 50764 35868 50932 35924
rect 51100 36258 51268 36260
rect 51100 36206 51214 36258
rect 51266 36206 51268 36258
rect 51100 36204 51268 36206
rect 51100 35924 51156 36204
rect 51212 36194 51268 36204
rect 51436 37772 51716 37828
rect 49420 35522 49476 35532
rect 49532 35698 49588 35710
rect 49532 35646 49534 35698
rect 49586 35646 49588 35698
rect 49532 35140 49588 35646
rect 49980 35588 50036 35598
rect 50764 35588 50820 35868
rect 51100 35698 51156 35868
rect 51100 35646 51102 35698
rect 51154 35646 51156 35698
rect 51100 35634 51156 35646
rect 49868 35476 49924 35486
rect 49532 35074 49588 35084
rect 49644 35474 49924 35476
rect 49644 35422 49870 35474
rect 49922 35422 49924 35474
rect 49644 35420 49924 35422
rect 49532 34244 49588 34254
rect 49644 34244 49700 35420
rect 49868 35410 49924 35420
rect 49532 34242 49700 34244
rect 49532 34190 49534 34242
rect 49586 34190 49700 34242
rect 49532 34188 49700 34190
rect 49868 34916 49924 34926
rect 49980 34916 50036 35532
rect 50540 35586 50820 35588
rect 50540 35534 50766 35586
rect 50818 35534 50820 35586
rect 50540 35532 50820 35534
rect 50540 35026 50596 35532
rect 50764 35522 50820 35532
rect 50540 34974 50542 35026
rect 50594 34974 50596 35026
rect 50540 34962 50596 34974
rect 49868 34914 50036 34916
rect 49868 34862 49870 34914
rect 49922 34862 50036 34914
rect 49868 34860 50036 34862
rect 51212 34916 51268 34926
rect 49532 34178 49588 34188
rect 49196 31500 49364 31556
rect 49420 34132 49476 34142
rect 49420 33122 49476 34076
rect 49756 34132 49812 34142
rect 49868 34132 49924 34860
rect 50876 34804 50932 34814
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 49756 34130 49924 34132
rect 49756 34078 49758 34130
rect 49810 34078 49924 34130
rect 49756 34076 49924 34078
rect 49980 34132 50036 34142
rect 49532 33572 49588 33582
rect 49756 33572 49812 34076
rect 49980 34038 50036 34076
rect 49532 33570 49812 33572
rect 49532 33518 49534 33570
rect 49586 33518 49812 33570
rect 49532 33516 49812 33518
rect 49532 33506 49588 33516
rect 49420 33070 49422 33122
rect 49474 33070 49476 33122
rect 49196 31444 49252 31500
rect 48748 31218 48916 31220
rect 48748 31166 48750 31218
rect 48802 31166 48916 31218
rect 48748 31164 48916 31166
rect 49084 31388 49252 31444
rect 48748 31154 48804 31164
rect 49084 31108 49140 31388
rect 49084 31052 49364 31108
rect 48076 28866 48692 28868
rect 48076 28814 48078 28866
rect 48130 28814 48692 28866
rect 48076 28812 48692 28814
rect 49084 30212 49140 30222
rect 48076 28802 48132 28812
rect 48300 28644 48356 28654
rect 48300 28642 48580 28644
rect 48300 28590 48302 28642
rect 48354 28590 48580 28642
rect 48300 28588 48580 28590
rect 48300 28578 48356 28588
rect 47964 27906 48020 27916
rect 48524 28420 48580 28588
rect 48636 28420 48692 28430
rect 48524 28418 48692 28420
rect 48524 28366 48638 28418
rect 48690 28366 48692 28418
rect 48524 28364 48692 28366
rect 47740 27860 47796 27870
rect 47404 27412 47460 27422
rect 46956 27300 47012 27310
rect 46956 26514 47012 27244
rect 47180 26962 47236 26974
rect 47180 26910 47182 26962
rect 47234 26910 47236 26962
rect 47180 26908 47236 26910
rect 46956 26462 46958 26514
rect 47010 26462 47012 26514
rect 46956 26450 47012 26462
rect 47068 26852 47236 26908
rect 46620 25330 46676 25340
rect 46732 25506 46900 25508
rect 46732 25454 46846 25506
rect 46898 25454 46900 25506
rect 46732 25452 46900 25454
rect 46396 24500 46452 24510
rect 46284 24498 46452 24500
rect 46284 24446 46398 24498
rect 46450 24446 46452 24498
rect 46284 24444 46452 24446
rect 46284 23492 46340 24444
rect 46396 24434 46452 24444
rect 46732 24164 46788 25452
rect 46844 25442 46900 25452
rect 46844 25282 46900 25294
rect 46844 25230 46846 25282
rect 46898 25230 46900 25282
rect 46844 24500 46900 25230
rect 46844 24276 46900 24444
rect 47068 24722 47124 26852
rect 47404 26514 47460 27356
rect 47404 26462 47406 26514
rect 47458 26462 47460 26514
rect 47404 26450 47460 26462
rect 47516 27074 47572 27086
rect 47516 27022 47518 27074
rect 47570 27022 47572 27074
rect 47516 26964 47572 27022
rect 47740 27074 47796 27804
rect 47740 27022 47742 27074
rect 47794 27022 47796 27074
rect 47740 27010 47796 27022
rect 48188 27746 48244 27758
rect 48188 27694 48190 27746
rect 48242 27694 48244 27746
rect 47516 26066 47572 26908
rect 48188 26964 48244 27694
rect 48412 27300 48468 27310
rect 48412 27206 48468 27244
rect 48188 26898 48244 26908
rect 48300 26962 48356 26974
rect 48300 26910 48302 26962
rect 48354 26910 48356 26962
rect 47516 26014 47518 26066
rect 47570 26014 47572 26066
rect 47180 25396 47236 25406
rect 47180 24834 47236 25340
rect 47180 24782 47182 24834
rect 47234 24782 47236 24834
rect 47180 24770 47236 24782
rect 47068 24670 47070 24722
rect 47122 24670 47124 24722
rect 47068 24388 47124 24670
rect 47068 24332 47236 24388
rect 46844 24220 47124 24276
rect 46732 24108 47012 24164
rect 46956 24050 47012 24108
rect 46956 23998 46958 24050
rect 47010 23998 47012 24050
rect 46508 23828 46564 23838
rect 46508 23734 46564 23772
rect 46284 23426 46340 23436
rect 46396 23604 46452 23614
rect 46396 23378 46452 23548
rect 46396 23326 46398 23378
rect 46450 23326 46452 23378
rect 46396 23314 46452 23326
rect 46956 23604 47012 23998
rect 46732 23044 46788 23054
rect 46732 22594 46788 22988
rect 46956 22820 47012 23548
rect 47068 23042 47124 24220
rect 47180 23716 47236 24332
rect 47516 24276 47572 26014
rect 47628 26852 47684 26862
rect 47628 25506 47684 26796
rect 48300 26516 48356 26910
rect 48524 26908 48580 28364
rect 48636 28354 48692 28364
rect 48636 27972 48692 27982
rect 48636 27878 48692 27916
rect 48972 27860 49028 27870
rect 48972 27186 49028 27804
rect 48972 27134 48974 27186
rect 49026 27134 49028 27186
rect 48972 27122 49028 27134
rect 48412 26852 48468 26862
rect 48524 26852 48804 26908
rect 48412 26758 48468 26796
rect 48300 26450 48356 26460
rect 48300 26292 48356 26302
rect 48300 26198 48356 26236
rect 47852 26178 47908 26190
rect 47852 26126 47854 26178
rect 47906 26126 47908 26178
rect 47852 26066 47908 26126
rect 47852 26014 47854 26066
rect 47906 26014 47908 26066
rect 47852 26002 47908 26014
rect 48748 26178 48804 26852
rect 48748 26126 48750 26178
rect 48802 26126 48804 26178
rect 47628 25454 47630 25506
rect 47682 25454 47684 25506
rect 47628 25442 47684 25454
rect 47740 25396 47796 25406
rect 47740 24946 47796 25340
rect 47964 25394 48020 25406
rect 47964 25342 47966 25394
rect 48018 25342 48020 25394
rect 47740 24894 47742 24946
rect 47794 24894 47796 24946
rect 47740 24882 47796 24894
rect 47852 25282 47908 25294
rect 47852 25230 47854 25282
rect 47906 25230 47908 25282
rect 47852 24948 47908 25230
rect 47852 24882 47908 24892
rect 47964 24724 48020 25342
rect 48412 25396 48468 25406
rect 48748 25396 48804 26126
rect 48860 26516 48916 26526
rect 48860 25618 48916 26460
rect 49084 25844 49140 30156
rect 49196 30100 49252 30110
rect 49196 30006 49252 30044
rect 49308 28754 49364 31052
rect 49308 28702 49310 28754
rect 49362 28702 49364 28754
rect 49308 26180 49364 28702
rect 49420 26908 49476 33070
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 49868 32788 49924 32798
rect 49868 32694 49924 32732
rect 50876 32786 50932 34748
rect 51212 34354 51268 34860
rect 51436 34692 51492 37772
rect 53228 37492 53284 40348
rect 53340 37940 53396 41132
rect 53340 37874 53396 37884
rect 53452 40404 53508 41468
rect 53564 41188 53620 42028
rect 53900 42018 53956 42028
rect 54236 41972 54292 45612
rect 54908 45668 54964 45678
rect 54908 45574 54964 45612
rect 55020 44548 55076 44558
rect 55020 43538 55076 44492
rect 55020 43486 55022 43538
rect 55074 43486 55076 43538
rect 55020 43474 55076 43486
rect 54908 43426 54964 43438
rect 54908 43374 54910 43426
rect 54962 43374 54964 43426
rect 54908 42868 54964 43374
rect 55804 42980 55860 46172
rect 56140 46002 56196 46620
rect 56140 45950 56142 46002
rect 56194 45950 56196 46002
rect 55916 45890 55972 45902
rect 55916 45838 55918 45890
rect 55970 45838 55972 45890
rect 55916 43708 55972 45838
rect 56140 44996 56196 45950
rect 56252 45220 56308 47068
rect 56476 46788 56532 47516
rect 56588 47346 56644 47358
rect 56588 47294 56590 47346
rect 56642 47294 56644 47346
rect 56588 47236 56644 47294
rect 56588 47170 56644 47180
rect 56532 46732 56644 46788
rect 56476 46722 56532 46732
rect 56476 46564 56532 46574
rect 56476 46470 56532 46508
rect 56588 46004 56644 46732
rect 56700 46228 56756 47628
rect 56812 47460 56868 47470
rect 56812 47366 56868 47404
rect 56700 46162 56756 46172
rect 56924 46564 56980 49644
rect 57036 49138 57092 55020
rect 57148 50370 57204 55804
rect 58044 51268 58100 51278
rect 58380 51268 58436 51278
rect 58044 51266 58324 51268
rect 58044 51214 58046 51266
rect 58098 51214 58324 51266
rect 58044 51212 58324 51214
rect 58044 51202 58100 51212
rect 57708 51156 57764 51166
rect 57260 51154 57764 51156
rect 57260 51102 57710 51154
rect 57762 51102 57764 51154
rect 57260 51100 57764 51102
rect 57260 50594 57316 51100
rect 57708 51090 57764 51100
rect 58156 50820 58212 50830
rect 57260 50542 57262 50594
rect 57314 50542 57316 50594
rect 57260 50530 57316 50542
rect 57484 50818 58212 50820
rect 57484 50766 58158 50818
rect 58210 50766 58212 50818
rect 57484 50764 58212 50766
rect 57484 50594 57540 50764
rect 58156 50754 58212 50764
rect 57484 50542 57486 50594
rect 57538 50542 57540 50594
rect 57484 50530 57540 50542
rect 58044 50484 58100 50494
rect 57148 50318 57150 50370
rect 57202 50318 57204 50370
rect 57148 50306 57204 50318
rect 57820 50482 58100 50484
rect 57820 50430 58046 50482
rect 58098 50430 58100 50482
rect 57820 50428 58100 50430
rect 57596 50036 57652 50046
rect 57036 49086 57038 49138
rect 57090 49086 57092 49138
rect 57036 49074 57092 49086
rect 57260 50034 57652 50036
rect 57260 49982 57598 50034
rect 57650 49982 57652 50034
rect 57260 49980 57652 49982
rect 57260 47796 57316 49980
rect 57596 49924 57652 49980
rect 57596 49858 57652 49868
rect 57820 50034 57876 50428
rect 58044 50418 58100 50428
rect 57820 49982 57822 50034
rect 57874 49982 57876 50034
rect 57484 49812 57540 49822
rect 57260 47730 57316 47740
rect 57372 49810 57540 49812
rect 57372 49758 57486 49810
rect 57538 49758 57540 49810
rect 57372 49756 57540 49758
rect 56588 45872 56644 45948
rect 56252 45154 56308 45164
rect 56364 45220 56420 45230
rect 56700 45220 56756 45230
rect 56364 45218 56532 45220
rect 56364 45166 56366 45218
rect 56418 45166 56532 45218
rect 56364 45164 56532 45166
rect 56364 45154 56420 45164
rect 56252 44996 56308 45006
rect 56140 44994 56308 44996
rect 56140 44942 56254 44994
rect 56306 44942 56308 44994
rect 56140 44940 56308 44942
rect 56252 44930 56308 44940
rect 55916 43652 56420 43708
rect 56364 43650 56420 43652
rect 56364 43598 56366 43650
rect 56418 43598 56420 43650
rect 56364 43586 56420 43598
rect 55804 42914 55860 42924
rect 56028 43538 56084 43550
rect 56252 43540 56308 43550
rect 56028 43486 56030 43538
rect 56082 43486 56084 43538
rect 55020 42868 55076 42878
rect 54908 42866 55076 42868
rect 54908 42814 55022 42866
rect 55074 42814 55076 42866
rect 54908 42812 55076 42814
rect 55020 42802 55076 42812
rect 55580 42756 55636 42766
rect 55916 42756 55972 42766
rect 55580 42754 55972 42756
rect 55580 42702 55582 42754
rect 55634 42702 55918 42754
rect 55970 42702 55972 42754
rect 55580 42700 55972 42702
rect 55580 42690 55636 42700
rect 55916 42690 55972 42700
rect 54908 42644 54964 42654
rect 54124 41916 54292 41972
rect 54684 42588 54908 42644
rect 54684 42084 54740 42588
rect 54908 42550 54964 42588
rect 55132 42532 55188 42542
rect 53788 41860 53844 41870
rect 53788 41412 53844 41804
rect 54012 41746 54068 41758
rect 54012 41694 54014 41746
rect 54066 41694 54068 41746
rect 53900 41636 53956 41646
rect 54012 41636 54068 41694
rect 53956 41580 54068 41636
rect 53900 41570 53956 41580
rect 54124 41524 54180 41916
rect 54012 41468 54180 41524
rect 54236 41746 54292 41758
rect 54236 41694 54238 41746
rect 54290 41694 54292 41746
rect 54236 41524 54292 41694
rect 53788 41410 53956 41412
rect 53788 41358 53790 41410
rect 53842 41358 53956 41410
rect 53788 41356 53956 41358
rect 53788 41346 53844 41356
rect 53676 41300 53732 41310
rect 53676 41206 53732 41244
rect 53564 41122 53620 41132
rect 53900 41186 53956 41356
rect 53900 41134 53902 41186
rect 53954 41134 53956 41186
rect 53900 41122 53956 41134
rect 53564 40964 53620 40974
rect 53564 40870 53620 40908
rect 53564 40404 53620 40414
rect 53452 40402 53620 40404
rect 53452 40350 53566 40402
rect 53618 40350 53620 40402
rect 53452 40348 53620 40350
rect 53228 37426 53284 37436
rect 53340 36484 53396 36494
rect 52332 36482 53396 36484
rect 52332 36430 53342 36482
rect 53394 36430 53396 36482
rect 52332 36428 53396 36430
rect 51996 35924 52052 35934
rect 51996 35830 52052 35868
rect 51548 35588 51604 35598
rect 51548 35586 51828 35588
rect 51548 35534 51550 35586
rect 51602 35534 51828 35586
rect 51548 35532 51828 35534
rect 51548 35522 51604 35532
rect 51772 35026 51828 35532
rect 51772 34974 51774 35026
rect 51826 34974 51828 35026
rect 51660 34916 51716 34926
rect 51660 34822 51716 34860
rect 51772 34804 51828 34974
rect 52108 34916 52164 34926
rect 51772 34748 52052 34804
rect 51436 34636 51940 34692
rect 51212 34302 51214 34354
rect 51266 34302 51268 34354
rect 51212 34290 51268 34302
rect 50876 32734 50878 32786
rect 50930 32734 50932 32786
rect 50876 32722 50932 32734
rect 49980 32564 50036 32574
rect 49980 32004 50036 32508
rect 50428 32564 50484 32574
rect 50428 32470 50484 32508
rect 50764 32564 50820 32574
rect 50764 32470 50820 32508
rect 50988 32562 51044 32574
rect 50988 32510 50990 32562
rect 51042 32510 51044 32562
rect 49868 31948 50036 32004
rect 49756 31778 49812 31790
rect 49756 31726 49758 31778
rect 49810 31726 49812 31778
rect 49756 31668 49812 31726
rect 49756 31444 49812 31612
rect 49644 31388 49812 31444
rect 49532 31108 49588 31118
rect 49644 31108 49700 31388
rect 49532 31106 49700 31108
rect 49532 31054 49534 31106
rect 49586 31054 49700 31106
rect 49532 31052 49700 31054
rect 49756 31108 49812 31118
rect 49532 31042 49588 31052
rect 49756 31014 49812 31052
rect 49868 30882 49924 31948
rect 49980 31778 50036 31790
rect 49980 31726 49982 31778
rect 50034 31726 50036 31778
rect 49980 31108 50036 31726
rect 50652 31668 50708 31678
rect 50988 31668 51044 32510
rect 50652 31666 51044 31668
rect 50652 31614 50654 31666
rect 50706 31614 51044 31666
rect 50652 31612 51044 31614
rect 50652 31602 50708 31612
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 49980 31042 50036 31052
rect 49868 30830 49870 30882
rect 49922 30830 49924 30882
rect 49868 30818 49924 30830
rect 50876 30994 50932 31006
rect 50876 30942 50878 30994
rect 50930 30942 50932 30994
rect 49868 30324 49924 30334
rect 49868 30230 49924 30268
rect 50092 30210 50148 30222
rect 50092 30158 50094 30210
rect 50146 30158 50148 30210
rect 50092 30100 50148 30158
rect 50764 30100 50820 30110
rect 50148 30044 50372 30100
rect 50092 30034 50148 30044
rect 49868 28642 49924 28654
rect 49868 28590 49870 28642
rect 49922 28590 49924 28642
rect 49868 27970 49924 28590
rect 49868 27918 49870 27970
rect 49922 27918 49924 27970
rect 49644 27748 49700 27758
rect 49532 27692 49644 27748
rect 49532 27188 49588 27692
rect 49644 27616 49700 27692
rect 49532 27094 49588 27132
rect 49756 27188 49812 27198
rect 49756 27094 49812 27132
rect 49420 26852 49588 26908
rect 49420 26180 49476 26190
rect 49308 26124 49420 26180
rect 49084 25788 49364 25844
rect 48860 25566 48862 25618
rect 48914 25566 48916 25618
rect 48860 25554 48916 25566
rect 49084 25508 49140 25518
rect 48972 25506 49140 25508
rect 48972 25454 49086 25506
rect 49138 25454 49140 25506
rect 48972 25452 49140 25454
rect 48972 25396 49028 25452
rect 49084 25442 49140 25452
rect 49196 25508 49252 25518
rect 48748 25340 49028 25396
rect 48412 24946 48468 25340
rect 48636 24948 48692 24958
rect 48412 24894 48414 24946
rect 48466 24894 48468 24946
rect 48412 24882 48468 24894
rect 48524 24892 48636 24948
rect 47964 24658 48020 24668
rect 47516 24210 47572 24220
rect 48524 24050 48580 24892
rect 48636 24854 48692 24892
rect 48748 24724 48804 24734
rect 48748 24630 48804 24668
rect 48524 23998 48526 24050
rect 48578 23998 48580 24050
rect 48524 23986 48580 23998
rect 47180 23650 47236 23660
rect 47516 23716 47572 23726
rect 47516 23622 47572 23660
rect 48972 23716 49028 25340
rect 49084 23828 49140 23838
rect 49196 23828 49252 25452
rect 49084 23826 49252 23828
rect 49084 23774 49086 23826
rect 49138 23774 49252 23826
rect 49084 23772 49252 23774
rect 49084 23762 49140 23772
rect 47068 22990 47070 23042
rect 47122 22990 47124 23042
rect 47068 22978 47124 22990
rect 47180 23154 47236 23166
rect 47180 23102 47182 23154
rect 47234 23102 47236 23154
rect 47180 22820 47236 23102
rect 46956 22764 47236 22820
rect 47852 23042 47908 23054
rect 47852 22990 47854 23042
rect 47906 22990 47908 23042
rect 46732 22542 46734 22594
rect 46786 22542 46788 22594
rect 46396 22484 46452 22494
rect 46172 22316 46340 22372
rect 46060 22278 46116 22316
rect 45948 22146 46004 22158
rect 45948 22094 45950 22146
rect 46002 22094 46004 22146
rect 45948 21700 46004 22094
rect 46172 22148 46228 22158
rect 46172 22054 46228 22092
rect 45948 21586 46004 21644
rect 45948 21534 45950 21586
rect 46002 21534 46004 21586
rect 45948 21522 46004 21534
rect 45836 20972 46004 21028
rect 45724 20916 45780 20926
rect 45612 20914 45780 20916
rect 45612 20862 45726 20914
rect 45778 20862 45780 20914
rect 45612 20860 45780 20862
rect 45724 20850 45780 20860
rect 44716 19124 44772 19134
rect 44716 19030 44772 19068
rect 45836 19122 45892 19134
rect 45836 19070 45838 19122
rect 45890 19070 45892 19122
rect 43484 18622 43486 18674
rect 43538 18622 43540 18674
rect 41804 18134 41860 18172
rect 42028 18226 42420 18228
rect 42028 18174 42142 18226
rect 42194 18174 42420 18226
rect 42028 18172 42420 18174
rect 42700 18396 43092 18452
rect 43148 18452 43204 18462
rect 41468 17500 41972 17556
rect 41468 17220 41524 17230
rect 41468 17106 41524 17164
rect 41468 17054 41470 17106
rect 41522 17054 41524 17106
rect 41468 17042 41524 17054
rect 41132 13906 41188 13916
rect 41244 16212 41300 16222
rect 41692 16212 41748 17500
rect 41916 17106 41972 17500
rect 41916 17054 41918 17106
rect 41970 17054 41972 17106
rect 41916 17042 41972 17054
rect 41244 16210 41748 16212
rect 41244 16158 41246 16210
rect 41298 16158 41694 16210
rect 41746 16158 41748 16210
rect 41244 16156 41748 16158
rect 40460 12402 40628 12404
rect 40460 12350 40462 12402
rect 40514 12350 40628 12402
rect 40460 12348 40628 12350
rect 40460 12338 40516 12348
rect 40572 12292 40628 12348
rect 40572 12226 40628 12236
rect 40796 13412 40852 13422
rect 40796 12962 40852 13356
rect 41244 13412 41300 16156
rect 41692 16146 41748 16156
rect 41804 15428 41860 15438
rect 41804 15334 41860 15372
rect 41244 13346 41300 13356
rect 41356 14980 41412 14990
rect 40796 12910 40798 12962
rect 40850 12910 40852 12962
rect 40684 12178 40740 12190
rect 40684 12126 40686 12178
rect 40738 12126 40740 12178
rect 40348 11890 40404 11900
rect 40572 12066 40628 12078
rect 40572 12014 40574 12066
rect 40626 12014 40628 12066
rect 40460 11844 40516 11854
rect 40460 11394 40516 11788
rect 40460 11342 40462 11394
rect 40514 11342 40516 11394
rect 40460 11330 40516 11342
rect 40572 11396 40628 12014
rect 40572 11330 40628 11340
rect 40124 11230 40126 11282
rect 40178 11230 40180 11282
rect 39788 10836 39844 10846
rect 39340 10834 39844 10836
rect 39340 10782 39342 10834
rect 39394 10782 39790 10834
rect 39842 10782 39844 10834
rect 39340 10780 39844 10782
rect 39340 10770 39396 10780
rect 39788 10770 39844 10780
rect 40124 10836 40180 11230
rect 40124 10770 40180 10780
rect 40348 11172 40404 11182
rect 40684 11172 40740 12126
rect 40796 11844 40852 12910
rect 41244 12964 41300 12974
rect 41244 12180 41300 12908
rect 41356 12850 41412 14924
rect 42028 14532 42084 18172
rect 42140 18162 42196 18172
rect 42476 17780 42532 17790
rect 42140 17220 42196 17230
rect 42140 16210 42196 17164
rect 42140 16158 42142 16210
rect 42194 16158 42196 16210
rect 42140 16146 42196 16158
rect 42364 15428 42420 15438
rect 42364 15334 42420 15372
rect 42028 14476 42196 14532
rect 42028 14306 42084 14318
rect 42028 14254 42030 14306
rect 42082 14254 42084 14306
rect 41468 13634 41524 13646
rect 41468 13582 41470 13634
rect 41522 13582 41524 13634
rect 41468 13412 41524 13582
rect 42028 13412 42084 14254
rect 41468 13346 41524 13356
rect 41916 13356 42028 13412
rect 41916 13074 41972 13356
rect 42028 13346 42084 13356
rect 41916 13022 41918 13074
rect 41970 13022 41972 13074
rect 41916 13010 41972 13022
rect 41356 12798 41358 12850
rect 41410 12798 41412 12850
rect 41356 12786 41412 12798
rect 41580 12738 41636 12750
rect 41580 12686 41582 12738
rect 41634 12686 41636 12738
rect 41580 12404 41636 12686
rect 41580 12338 41636 12348
rect 42028 12404 42084 12414
rect 42028 12310 42084 12348
rect 41804 12292 41860 12302
rect 41580 12180 41636 12190
rect 41244 12178 41636 12180
rect 41244 12126 41582 12178
rect 41634 12126 41636 12178
rect 41244 12124 41636 12126
rect 41580 12114 41636 12124
rect 41692 12066 41748 12078
rect 41692 12014 41694 12066
rect 41746 12014 41748 12066
rect 40796 11778 40852 11788
rect 41132 11956 41188 11966
rect 41132 11508 41188 11900
rect 41580 11844 41636 11854
rect 41244 11620 41300 11630
rect 41468 11620 41524 11630
rect 41244 11618 41524 11620
rect 41244 11566 41246 11618
rect 41298 11566 41470 11618
rect 41522 11566 41524 11618
rect 41244 11564 41524 11566
rect 41244 11554 41300 11564
rect 41468 11554 41524 11564
rect 40348 11170 40740 11172
rect 40348 11118 40350 11170
rect 40402 11118 40740 11170
rect 40348 11116 40740 11118
rect 40908 11506 41188 11508
rect 40908 11454 41134 11506
rect 41186 11454 41188 11506
rect 40908 11452 41188 11454
rect 40236 10498 40292 10510
rect 40236 10446 40238 10498
rect 40290 10446 40292 10498
rect 39228 10388 39284 10398
rect 39116 10386 39284 10388
rect 39116 10334 39230 10386
rect 39282 10334 39284 10386
rect 39116 10332 39284 10334
rect 39228 10322 39284 10332
rect 40236 10386 40292 10446
rect 40236 10334 40238 10386
rect 40290 10334 40292 10386
rect 40236 10322 40292 10334
rect 38556 9874 38612 9884
rect 38892 10052 38948 10062
rect 38780 9044 38836 9082
rect 38780 8978 38836 8988
rect 38892 8428 38948 9996
rect 39340 10052 39396 10062
rect 39228 9828 39284 9838
rect 39340 9828 39396 9996
rect 40348 10052 40404 11116
rect 40684 10836 40740 10846
rect 40684 10742 40740 10780
rect 40348 9986 40404 9996
rect 40460 9940 40516 9950
rect 39228 9826 39396 9828
rect 39228 9774 39230 9826
rect 39282 9774 39396 9826
rect 39228 9772 39396 9774
rect 39228 9762 39284 9772
rect 39004 9602 39060 9614
rect 39004 9550 39006 9602
rect 39058 9550 39060 9602
rect 39004 9156 39060 9550
rect 39116 9156 39172 9166
rect 39004 9154 39172 9156
rect 39004 9102 39118 9154
rect 39170 9102 39172 9154
rect 39004 9100 39172 9102
rect 39116 9090 39172 9100
rect 39228 9042 39284 9054
rect 39228 8990 39230 9042
rect 39282 8990 39284 9042
rect 39004 8932 39060 8942
rect 39228 8932 39284 8990
rect 39004 8930 39284 8932
rect 39004 8878 39006 8930
rect 39058 8878 39284 8930
rect 39004 8876 39284 8878
rect 39004 8866 39060 8876
rect 38892 8372 39172 8428
rect 39116 8258 39172 8372
rect 39116 8206 39118 8258
rect 39170 8206 39172 8258
rect 39116 8194 39172 8206
rect 39340 8258 39396 9772
rect 40012 9828 40068 9838
rect 40012 9734 40068 9772
rect 40460 9826 40516 9884
rect 40460 9774 40462 9826
rect 40514 9774 40516 9826
rect 40460 9762 40516 9774
rect 40908 9828 40964 11452
rect 41132 11442 41188 11452
rect 40684 9716 40740 9726
rect 40908 9696 40964 9772
rect 41020 11284 41076 11294
rect 39564 9042 39620 9054
rect 39564 8990 39566 9042
rect 39618 8990 39620 9042
rect 39564 8482 39620 8990
rect 40460 9044 40516 9054
rect 40460 8950 40516 8988
rect 40684 9042 40740 9660
rect 40684 8990 40686 9042
rect 40738 8990 40740 9042
rect 40684 8978 40740 8990
rect 40796 9602 40852 9614
rect 40796 9550 40798 9602
rect 40850 9550 40852 9602
rect 39564 8430 39566 8482
rect 39618 8430 39620 8482
rect 39564 8418 39620 8430
rect 39788 8930 39844 8942
rect 39788 8878 39790 8930
rect 39842 8878 39844 8930
rect 39340 8206 39342 8258
rect 39394 8206 39396 8258
rect 39340 8194 39396 8206
rect 39676 8258 39732 8270
rect 39676 8206 39678 8258
rect 39730 8206 39732 8258
rect 38556 8146 38612 8158
rect 38556 8094 38558 8146
rect 38610 8094 38612 8146
rect 38556 7476 38612 8094
rect 39564 7700 39620 7710
rect 39676 7700 39732 8206
rect 39788 8260 39844 8878
rect 40796 8428 40852 9550
rect 41020 9604 41076 11228
rect 41580 10834 41636 11788
rect 41580 10782 41582 10834
rect 41634 10782 41636 10834
rect 41580 10770 41636 10782
rect 41132 9828 41188 9838
rect 41132 9826 41636 9828
rect 41132 9774 41134 9826
rect 41186 9774 41636 9826
rect 41132 9772 41636 9774
rect 41132 9762 41188 9772
rect 41020 9548 41412 9604
rect 40796 8372 41188 8428
rect 39788 8194 39844 8204
rect 40124 8260 40180 8270
rect 39900 8036 39956 8046
rect 39900 7942 39956 7980
rect 39564 7698 39732 7700
rect 39564 7646 39566 7698
rect 39618 7646 39732 7698
rect 39564 7644 39732 7646
rect 39564 7634 39620 7644
rect 38556 7410 38612 7420
rect 39452 5908 39508 5918
rect 39676 5908 39732 7644
rect 39900 7476 39956 7486
rect 39900 7382 39956 7420
rect 40124 7474 40180 8204
rect 40796 8260 40852 8270
rect 40796 8166 40852 8204
rect 40572 8036 40628 8046
rect 40572 7942 40628 7980
rect 40908 8034 40964 8046
rect 40908 7982 40910 8034
rect 40962 7982 40964 8034
rect 40124 7422 40126 7474
rect 40178 7422 40180 7474
rect 40124 7410 40180 7422
rect 39508 5852 39620 5908
rect 39452 5814 39508 5852
rect 37660 5124 37716 5134
rect 37660 5030 37716 5068
rect 38108 5124 38164 5134
rect 38220 5124 38276 5180
rect 39228 5794 39284 5806
rect 39228 5742 39230 5794
rect 39282 5742 39284 5794
rect 38108 5122 38276 5124
rect 38108 5070 38110 5122
rect 38162 5070 38276 5122
rect 38108 5068 38276 5070
rect 38556 5124 38612 5134
rect 38108 5058 38164 5068
rect 38556 5030 38612 5068
rect 39228 5124 39284 5742
rect 39564 5124 39620 5852
rect 39676 5906 39956 5908
rect 39676 5854 39678 5906
rect 39730 5854 39956 5906
rect 39676 5852 39956 5854
rect 39676 5842 39732 5852
rect 39676 5124 39732 5134
rect 39564 5122 39732 5124
rect 39564 5070 39678 5122
rect 39730 5070 39732 5122
rect 39564 5068 39732 5070
rect 39228 4992 39284 5068
rect 39676 5058 39732 5068
rect 39900 5122 39956 5852
rect 39900 5070 39902 5122
rect 39954 5070 39956 5122
rect 39900 5058 39956 5070
rect 40124 5682 40180 5694
rect 40124 5630 40126 5682
rect 40178 5630 40180 5682
rect 39788 4900 39844 4910
rect 39788 4806 39844 4844
rect 40124 4564 40180 5630
rect 40908 5348 40964 7982
rect 41020 8034 41076 8046
rect 41020 7982 41022 8034
rect 41074 7982 41076 8034
rect 41020 7476 41076 7982
rect 41020 7410 41076 7420
rect 41132 6804 41188 8372
rect 41356 6916 41412 9548
rect 41580 9492 41636 9772
rect 41692 9716 41748 12014
rect 41804 11618 41860 12236
rect 42140 12068 42196 14476
rect 41804 11566 41806 11618
rect 41858 11566 41860 11618
rect 41804 11506 41860 11566
rect 41804 11454 41806 11506
rect 41858 11454 41860 11506
rect 41804 11442 41860 11454
rect 42028 12012 42196 12068
rect 42252 13412 42308 13422
rect 41692 9622 41748 9660
rect 41916 10052 41972 10062
rect 41804 9602 41860 9614
rect 41804 9550 41806 9602
rect 41858 9550 41860 9602
rect 41804 9492 41860 9550
rect 41580 9436 41860 9492
rect 41916 9156 41972 9996
rect 41916 9024 41972 9100
rect 42028 9826 42084 12012
rect 42252 11956 42308 13356
rect 42140 11508 42196 11518
rect 42252 11508 42308 11900
rect 42140 11506 42308 11508
rect 42140 11454 42142 11506
rect 42194 11454 42308 11506
rect 42140 11452 42308 11454
rect 42364 11732 42420 11742
rect 42140 11442 42196 11452
rect 42364 10834 42420 11676
rect 42476 11396 42532 17724
rect 42588 17666 42644 17678
rect 42588 17614 42590 17666
rect 42642 17614 42644 17666
rect 42588 17220 42644 17614
rect 42588 17154 42644 17164
rect 42700 16884 42756 18396
rect 42812 18228 42868 18238
rect 42812 17666 42868 18172
rect 42812 17614 42814 17666
rect 42866 17614 42868 17666
rect 42812 17556 42868 17614
rect 43036 17668 43092 17678
rect 42812 17490 42868 17500
rect 42924 17554 42980 17566
rect 42924 17502 42926 17554
rect 42978 17502 42980 17554
rect 42924 17108 42980 17502
rect 42924 17042 42980 17052
rect 43036 17106 43092 17612
rect 43036 17054 43038 17106
rect 43090 17054 43092 17106
rect 43036 17042 43092 17054
rect 43148 17106 43204 18396
rect 43484 17780 43540 18622
rect 44044 18732 44324 18788
rect 44380 19010 44436 19022
rect 44380 18958 44382 19010
rect 44434 18958 44436 19010
rect 43596 18452 43652 18462
rect 43596 18358 43652 18396
rect 43708 18450 43764 18462
rect 43708 18398 43710 18450
rect 43762 18398 43764 18450
rect 43484 17714 43540 17724
rect 43708 17668 43764 18398
rect 43820 17780 43876 17790
rect 43820 17686 43876 17724
rect 43708 17574 43764 17612
rect 44044 17332 44100 18732
rect 44156 18452 44212 18462
rect 44380 18452 44436 18958
rect 44156 18450 44436 18452
rect 44156 18398 44158 18450
rect 44210 18398 44436 18450
rect 44156 18396 44436 18398
rect 45500 18676 45556 18686
rect 44156 18386 44212 18396
rect 44492 18340 44548 18350
rect 44044 17266 44100 17276
rect 44380 18284 44492 18340
rect 44380 17556 44436 18284
rect 44492 18246 44548 18284
rect 44492 17780 44548 17790
rect 44492 17686 44548 17724
rect 45500 17556 45556 18620
rect 45612 18564 45668 18574
rect 45836 18564 45892 19070
rect 45668 18508 45892 18564
rect 45612 18450 45668 18508
rect 45612 18398 45614 18450
rect 45666 18398 45668 18450
rect 45612 18386 45668 18398
rect 45948 18340 46004 20972
rect 46060 20244 46116 20254
rect 46060 20150 46116 20188
rect 45948 18274 46004 18284
rect 46060 19460 46116 19470
rect 46060 18338 46116 19404
rect 46060 18286 46062 18338
rect 46114 18286 46116 18338
rect 46060 18274 46116 18286
rect 45500 17500 45780 17556
rect 43148 17054 43150 17106
rect 43202 17054 43204 17106
rect 43148 16996 43204 17054
rect 43260 17108 43316 17118
rect 43260 17014 43316 17052
rect 44268 17108 44324 17118
rect 43148 16930 43204 16940
rect 43484 16996 43540 17006
rect 42700 16818 42756 16828
rect 42812 16882 42868 16894
rect 42812 16830 42814 16882
rect 42866 16830 42868 16882
rect 42812 16322 42868 16830
rect 42924 16884 42980 16894
rect 42980 16828 43092 16884
rect 42924 16790 42980 16828
rect 42812 16270 42814 16322
rect 42866 16270 42868 16322
rect 42812 16258 42868 16270
rect 42924 16100 42980 16110
rect 42700 15986 42756 15998
rect 42700 15934 42702 15986
rect 42754 15934 42756 15986
rect 42588 15316 42644 15326
rect 42588 15222 42644 15260
rect 42700 14980 42756 15934
rect 42812 15988 42868 15998
rect 42812 15894 42868 15932
rect 42924 15538 42980 16044
rect 42924 15486 42926 15538
rect 42978 15486 42980 15538
rect 42924 15474 42980 15486
rect 42700 13858 42756 14924
rect 43036 14084 43092 16828
rect 43372 16100 43428 16110
rect 43372 16006 43428 16044
rect 43484 15876 43540 16940
rect 43820 16884 43876 16894
rect 43820 16790 43876 16828
rect 43708 16660 43764 16670
rect 43708 16100 43764 16604
rect 43708 16098 43988 16100
rect 43708 16046 43710 16098
rect 43762 16046 43988 16098
rect 43708 16044 43988 16046
rect 43708 16034 43764 16044
rect 43260 15820 43540 15876
rect 43708 15876 43764 15886
rect 43148 15428 43204 15438
rect 43148 14754 43204 15372
rect 43148 14702 43150 14754
rect 43202 14702 43204 14754
rect 43148 14642 43204 14702
rect 43148 14590 43150 14642
rect 43202 14590 43204 14642
rect 43148 14578 43204 14590
rect 43036 14028 43204 14084
rect 42700 13806 42702 13858
rect 42754 13806 42756 13858
rect 42700 13794 42756 13806
rect 43036 13860 43092 13870
rect 43036 13766 43092 13804
rect 43148 12962 43204 14028
rect 43260 13746 43316 15820
rect 43708 15782 43764 15820
rect 43932 15538 43988 16044
rect 44044 15988 44100 15998
rect 44044 15986 44212 15988
rect 44044 15934 44046 15986
rect 44098 15934 44212 15986
rect 44044 15932 44212 15934
rect 44044 15922 44100 15932
rect 43932 15486 43934 15538
rect 43986 15486 43988 15538
rect 43932 15474 43988 15486
rect 43708 15428 43764 15438
rect 43708 15334 43764 15372
rect 43484 15316 43540 15326
rect 43484 15222 43540 15260
rect 43596 15202 43652 15214
rect 43596 15150 43598 15202
rect 43650 15150 43652 15202
rect 43260 13694 43262 13746
rect 43314 13694 43316 13746
rect 43260 13412 43316 13694
rect 43260 13346 43316 13356
rect 43484 14754 43540 14766
rect 43484 14702 43486 14754
rect 43538 14702 43540 14754
rect 43148 12910 43150 12962
rect 43202 12910 43204 12962
rect 43036 12404 43092 12414
rect 43148 12404 43204 12910
rect 43484 12628 43540 14702
rect 43596 14532 43652 15150
rect 44044 14532 44100 14542
rect 43596 14530 44100 14532
rect 43596 14478 44046 14530
rect 44098 14478 44100 14530
rect 43596 14476 44100 14478
rect 44044 14466 44100 14476
rect 44156 14308 44212 15932
rect 44268 15148 44324 17052
rect 44380 17106 44436 17500
rect 44380 17054 44382 17106
rect 44434 17054 44436 17106
rect 44380 17042 44436 17054
rect 45164 17108 45220 17118
rect 45164 17014 45220 17052
rect 45612 17108 45668 17118
rect 45612 17014 45668 17052
rect 44716 16996 44772 17006
rect 44716 16902 44772 16940
rect 45724 16322 45780 17500
rect 45724 16270 45726 16322
rect 45778 16270 45780 16322
rect 44604 15988 44660 15998
rect 44604 15428 44660 15932
rect 45052 15428 45108 15438
rect 44604 15372 45052 15428
rect 44604 15148 44660 15372
rect 45052 15296 45108 15372
rect 45612 15428 45668 15438
rect 45724 15428 45780 16270
rect 45948 17108 46004 17118
rect 45948 15986 46004 17052
rect 46284 17108 46340 22316
rect 46396 20914 46452 22428
rect 46732 22484 46788 22542
rect 46732 22418 46788 22428
rect 47740 22260 47796 22270
rect 47740 22166 47796 22204
rect 46844 22146 46900 22158
rect 46844 22094 46846 22146
rect 46898 22094 46900 22146
rect 46844 21812 46900 22094
rect 46844 21746 46900 21756
rect 46956 22146 47012 22158
rect 46956 22094 46958 22146
rect 47010 22094 47012 22146
rect 46620 21474 46676 21486
rect 46620 21422 46622 21474
rect 46674 21422 46676 21474
rect 46620 21140 46676 21422
rect 46620 21074 46676 21084
rect 46396 20862 46398 20914
rect 46450 20862 46452 20914
rect 46396 20850 46452 20862
rect 46508 20804 46564 20814
rect 46956 20804 47012 22094
rect 47628 22148 47684 22158
rect 47628 22054 47684 22092
rect 47404 21812 47460 21822
rect 47852 21812 47908 22990
rect 48300 23044 48356 23054
rect 48300 22950 48356 22988
rect 48188 22484 48244 22494
rect 48244 22428 48356 22484
rect 48188 22390 48244 22428
rect 47404 21718 47460 21756
rect 47740 21756 47908 21812
rect 47180 21586 47236 21598
rect 47180 21534 47182 21586
rect 47234 21534 47236 21586
rect 47180 21140 47236 21534
rect 47292 21588 47348 21598
rect 47292 21494 47348 21532
rect 47180 21074 47236 21084
rect 46508 20802 47012 20804
rect 46508 20750 46510 20802
rect 46562 20750 47012 20802
rect 46508 20748 47012 20750
rect 46508 20244 46564 20748
rect 46508 20178 46564 20188
rect 46396 19348 46452 19358
rect 46396 19346 46900 19348
rect 46396 19294 46398 19346
rect 46450 19294 46900 19346
rect 46396 19292 46900 19294
rect 46396 19282 46452 19292
rect 46844 19234 46900 19292
rect 46844 19182 46846 19234
rect 46898 19182 46900 19234
rect 46844 19170 46900 19182
rect 47404 19124 47460 19134
rect 47404 19030 47460 19068
rect 46508 19012 46564 19022
rect 46508 18450 46564 18956
rect 47292 19012 47348 19022
rect 47292 18918 47348 18956
rect 47516 19010 47572 19022
rect 47516 18958 47518 19010
rect 47570 18958 47572 19010
rect 46508 18398 46510 18450
rect 46562 18398 46564 18450
rect 46508 17666 46564 18398
rect 46620 17780 46676 17790
rect 46620 17686 46676 17724
rect 47516 17780 47572 18958
rect 47740 18452 47796 21756
rect 48300 21700 48356 22428
rect 48636 22148 48692 22158
rect 48524 22146 48692 22148
rect 48524 22094 48638 22146
rect 48690 22094 48692 22146
rect 48524 22092 48692 22094
rect 47964 21698 48356 21700
rect 47964 21646 48302 21698
rect 48354 21646 48356 21698
rect 47964 21644 48356 21646
rect 47852 21586 47908 21598
rect 47852 21534 47854 21586
rect 47906 21534 47908 21586
rect 47852 21474 47908 21534
rect 47852 21422 47854 21474
rect 47906 21422 47908 21474
rect 47852 21410 47908 21422
rect 47852 21140 47908 21150
rect 47852 20802 47908 21084
rect 47852 20750 47854 20802
rect 47906 20750 47908 20802
rect 47852 20738 47908 20750
rect 47852 20244 47908 20254
rect 47964 20244 48020 21644
rect 48300 21634 48356 21644
rect 48412 21700 48468 21710
rect 48524 21700 48580 22092
rect 48636 22082 48692 22092
rect 48412 21698 48580 21700
rect 48412 21646 48414 21698
rect 48466 21646 48580 21698
rect 48412 21644 48580 21646
rect 48412 21634 48468 21644
rect 48076 21474 48132 21486
rect 48076 21422 48078 21474
rect 48130 21422 48132 21474
rect 48076 21364 48132 21422
rect 48412 21364 48468 21374
rect 48076 21362 48468 21364
rect 48076 21310 48414 21362
rect 48466 21310 48468 21362
rect 48076 21308 48468 21310
rect 48412 21298 48468 21308
rect 47852 20242 48020 20244
rect 47852 20190 47854 20242
rect 47906 20190 48020 20242
rect 47852 20188 48020 20190
rect 48300 20244 48356 20254
rect 48524 20244 48580 21644
rect 48356 20188 48580 20244
rect 48636 20690 48692 20702
rect 48636 20638 48638 20690
rect 48690 20638 48692 20690
rect 47852 20178 47908 20188
rect 48300 20150 48356 20188
rect 48636 19236 48692 20638
rect 48636 19170 48692 19180
rect 47852 18452 47908 18462
rect 47740 18450 47908 18452
rect 47740 18398 47854 18450
rect 47906 18398 47908 18450
rect 47740 18396 47908 18398
rect 47516 17714 47572 17724
rect 46508 17614 46510 17666
rect 46562 17614 46564 17666
rect 46508 17602 46564 17614
rect 47852 17668 47908 18396
rect 47852 17602 47908 17612
rect 48076 18452 48132 18462
rect 46284 17042 46340 17052
rect 47404 17554 47460 17566
rect 47404 17502 47406 17554
rect 47458 17502 47460 17554
rect 46060 16212 46116 16222
rect 46620 16212 46676 16222
rect 46060 16210 46676 16212
rect 46060 16158 46062 16210
rect 46114 16158 46622 16210
rect 46674 16158 46676 16210
rect 46060 16156 46676 16158
rect 46060 16146 46116 16156
rect 45948 15934 45950 15986
rect 46002 15934 46004 15986
rect 45948 15922 46004 15934
rect 45612 15426 45780 15428
rect 45612 15374 45614 15426
rect 45666 15374 45780 15426
rect 45612 15372 45780 15374
rect 45836 15538 45892 15550
rect 45836 15486 45838 15538
rect 45890 15486 45892 15538
rect 45612 15362 45668 15372
rect 44268 15092 44436 15148
rect 44268 14642 44324 14654
rect 44268 14590 44270 14642
rect 44322 14590 44324 14642
rect 44268 14308 44324 14590
rect 43820 14252 44324 14308
rect 43708 13860 43764 13870
rect 43596 13522 43652 13534
rect 43596 13470 43598 13522
rect 43650 13470 43652 13522
rect 43596 12962 43652 13470
rect 43596 12910 43598 12962
rect 43650 12910 43652 12962
rect 43596 12898 43652 12910
rect 43708 12852 43764 13804
rect 43820 13074 43876 14252
rect 44156 13972 44212 13982
rect 44380 13972 44436 15092
rect 44156 13970 44436 13972
rect 44156 13918 44158 13970
rect 44210 13918 44436 13970
rect 44156 13916 44436 13918
rect 44492 15092 44660 15148
rect 44156 13860 44212 13916
rect 44156 13794 44212 13804
rect 43820 13022 43822 13074
rect 43874 13022 43876 13074
rect 43820 13010 43876 13022
rect 43708 12796 43876 12852
rect 43484 12572 43652 12628
rect 43484 12404 43540 12414
rect 43036 12402 43540 12404
rect 43036 12350 43038 12402
rect 43090 12350 43486 12402
rect 43538 12350 43540 12402
rect 43036 12348 43540 12350
rect 43036 12338 43092 12348
rect 42588 12292 42644 12302
rect 42588 12198 42644 12236
rect 42812 11732 42868 11742
rect 42812 11618 42868 11676
rect 42812 11566 42814 11618
rect 42866 11566 42868 11618
rect 42812 11554 42868 11566
rect 43484 11508 43540 12348
rect 43596 12404 43652 12572
rect 43596 11732 43652 12348
rect 43596 11666 43652 11676
rect 43484 11442 43540 11452
rect 42476 11340 43092 11396
rect 42364 10782 42366 10834
rect 42418 10782 42420 10834
rect 42364 10770 42420 10782
rect 42700 10834 42756 11340
rect 43036 11282 43092 11340
rect 43036 11230 43038 11282
rect 43090 11230 43092 11282
rect 43036 11218 43092 11230
rect 42924 11172 42980 11182
rect 42924 11078 42980 11116
rect 43708 11172 43764 11182
rect 42700 10782 42702 10834
rect 42754 10782 42756 10834
rect 42028 9774 42030 9826
rect 42082 9774 42084 9826
rect 42028 9492 42084 9774
rect 42028 9266 42084 9436
rect 42028 9214 42030 9266
rect 42082 9214 42084 9266
rect 42028 9044 42084 9214
rect 42252 9380 42308 9390
rect 42700 9380 42756 10782
rect 43708 10722 43764 11116
rect 43708 10670 43710 10722
rect 43762 10670 43764 10722
rect 43708 10658 43764 10670
rect 43148 10500 43204 10510
rect 43148 10498 43316 10500
rect 43148 10446 43150 10498
rect 43202 10446 43316 10498
rect 43148 10444 43316 10446
rect 43148 10434 43204 10444
rect 43260 9938 43316 10444
rect 43260 9886 43262 9938
rect 43314 9886 43316 9938
rect 43036 9828 43092 9838
rect 43036 9604 43092 9772
rect 43036 9538 43092 9548
rect 43260 9716 43316 9886
rect 43148 9380 43204 9390
rect 42700 9324 42980 9380
rect 42252 9266 42308 9324
rect 42252 9214 42254 9266
rect 42306 9214 42308 9266
rect 42252 9202 42308 9214
rect 42028 8428 42084 8988
rect 41580 8372 42084 8428
rect 42588 9156 42644 9166
rect 42700 9156 42756 9166
rect 42644 9154 42756 9156
rect 42644 9102 42702 9154
rect 42754 9102 42756 9154
rect 42644 9100 42756 9102
rect 41580 8370 41636 8372
rect 41580 8318 41582 8370
rect 41634 8318 41636 8370
rect 41580 8306 41636 8318
rect 42028 8260 42084 8270
rect 41580 7700 41636 7710
rect 42028 7700 42084 8204
rect 42476 8260 42532 8270
rect 42588 8260 42644 9100
rect 42700 9090 42756 9100
rect 42924 9044 42980 9324
rect 43148 9266 43204 9324
rect 43148 9214 43150 9266
rect 43202 9214 43204 9266
rect 43148 9202 43204 9214
rect 43260 9268 43316 9660
rect 43260 9202 43316 9212
rect 43708 9714 43764 9726
rect 43708 9662 43710 9714
rect 43762 9662 43764 9714
rect 43708 9156 43764 9662
rect 43708 9090 43764 9100
rect 43820 9154 43876 12796
rect 43932 12404 43988 12414
rect 43932 12310 43988 12348
rect 43932 11620 43988 11630
rect 43932 10722 43988 11564
rect 44044 11508 44100 11518
rect 44044 11394 44100 11452
rect 44044 11342 44046 11394
rect 44098 11342 44100 11394
rect 44044 11330 44100 11342
rect 44492 11172 44548 15092
rect 44716 14644 44772 14654
rect 44716 14550 44772 14588
rect 45724 14084 45780 14094
rect 45612 13636 45668 13646
rect 45612 13542 45668 13580
rect 45724 13074 45780 14028
rect 45724 13022 45726 13074
rect 45778 13022 45780 13074
rect 45724 13010 45780 13022
rect 45164 12066 45220 12078
rect 45164 12014 45166 12066
rect 45218 12014 45220 12066
rect 45164 11508 45220 12014
rect 45164 11442 45220 11452
rect 45500 11508 45556 11518
rect 45500 11414 45556 11452
rect 43932 10670 43934 10722
rect 43986 10670 43988 10722
rect 43932 10658 43988 10670
rect 44044 11116 44548 11172
rect 44604 11396 44660 11406
rect 43820 9102 43822 9154
rect 43874 9102 43876 9154
rect 42924 9042 43092 9044
rect 42924 8990 42926 9042
rect 42978 8990 43092 9042
rect 42924 8988 43092 8990
rect 42924 8978 42980 8988
rect 42812 8930 42868 8942
rect 42812 8878 42814 8930
rect 42866 8878 42868 8930
rect 42476 8258 42644 8260
rect 42476 8206 42478 8258
rect 42530 8206 42644 8258
rect 42476 8204 42644 8206
rect 42700 8260 42756 8270
rect 42812 8260 42868 8878
rect 42924 8260 42980 8270
rect 42812 8258 42980 8260
rect 42812 8206 42926 8258
rect 42978 8206 42980 8258
rect 42812 8204 42980 8206
rect 42476 8194 42532 8204
rect 42700 8166 42756 8204
rect 41580 7698 42084 7700
rect 41580 7646 41582 7698
rect 41634 7646 42030 7698
rect 42082 7646 42084 7698
rect 41580 7644 42084 7646
rect 41580 7634 41636 7644
rect 42028 7634 42084 7644
rect 42588 8034 42644 8046
rect 42588 7982 42590 8034
rect 42642 7982 42644 8034
rect 42476 7362 42532 7374
rect 42476 7310 42478 7362
rect 42530 7310 42532 7362
rect 41356 6860 41972 6916
rect 40908 5282 40964 5292
rect 41020 6748 41636 6804
rect 41020 5122 41076 6748
rect 41580 6018 41636 6748
rect 41580 5966 41582 6018
rect 41634 5966 41636 6018
rect 41580 5954 41636 5966
rect 41804 5682 41860 5694
rect 41804 5630 41806 5682
rect 41858 5630 41860 5682
rect 41468 5348 41524 5358
rect 41804 5348 41860 5630
rect 41468 5254 41524 5292
rect 41580 5292 41860 5348
rect 41356 5124 41412 5134
rect 41580 5124 41636 5292
rect 41916 5236 41972 6860
rect 42476 6020 42532 7310
rect 42588 6580 42644 7982
rect 42924 7362 42980 8204
rect 43036 8260 43092 8988
rect 43148 8372 43204 8382
rect 43148 8278 43204 8316
rect 43036 8194 43092 8204
rect 43148 7476 43204 7486
rect 43148 7382 43204 7420
rect 43820 7476 43876 9102
rect 43932 8820 43988 8830
rect 44044 8820 44100 11116
rect 44156 10836 44212 10846
rect 44604 10836 44660 11340
rect 45724 11396 45780 11406
rect 45724 11302 45780 11340
rect 44716 11284 44772 11294
rect 45836 11284 45892 15486
rect 45948 15428 46004 15438
rect 45948 15334 46004 15372
rect 46172 15426 46228 16156
rect 46620 16146 46676 16156
rect 46172 15374 46174 15426
rect 46226 15374 46228 15426
rect 46172 15362 46228 15374
rect 46732 15874 46788 15886
rect 46732 15822 46734 15874
rect 46786 15822 46788 15874
rect 46732 15148 46788 15822
rect 47180 15428 47236 15438
rect 46844 15426 47236 15428
rect 46844 15374 47182 15426
rect 47234 15374 47236 15426
rect 46844 15372 47236 15374
rect 46844 15148 46900 15372
rect 47180 15362 47236 15372
rect 46732 15092 46900 15148
rect 47292 15204 47348 15242
rect 47292 15138 47348 15148
rect 46508 14644 46564 14654
rect 46508 14550 46564 14588
rect 46844 14530 46900 15092
rect 46956 15090 47012 15102
rect 46956 15038 46958 15090
rect 47010 15038 47012 15090
rect 46956 14644 47012 15038
rect 47404 14644 47460 17502
rect 48076 17556 48132 18396
rect 48748 18338 48804 18350
rect 48748 18286 48750 18338
rect 48802 18286 48804 18338
rect 48748 17780 48804 18286
rect 48972 18340 49028 23660
rect 49196 23044 49252 23772
rect 49308 23380 49364 25788
rect 49420 25508 49476 26124
rect 49532 25956 49588 26852
rect 49756 26852 49812 26862
rect 49868 26852 49924 27918
rect 50092 28642 50148 28654
rect 50092 28590 50094 28642
rect 50146 28590 50148 28642
rect 50092 27748 50148 28590
rect 50316 28420 50372 30044
rect 50764 30006 50820 30044
rect 50876 29988 50932 30942
rect 50988 30884 51044 31612
rect 51212 32564 51268 32574
rect 51100 30884 51156 30894
rect 50988 30882 51156 30884
rect 50988 30830 51102 30882
rect 51154 30830 51156 30882
rect 50988 30828 51156 30830
rect 51100 30818 51156 30828
rect 51212 29988 51268 32508
rect 51548 32450 51604 32462
rect 51548 32398 51550 32450
rect 51602 32398 51604 32450
rect 51548 31948 51604 32398
rect 51548 31892 51828 31948
rect 51772 31778 51828 31892
rect 51772 31726 51774 31778
rect 51826 31726 51828 31778
rect 51548 31108 51604 31118
rect 51548 31014 51604 31052
rect 51772 30884 51828 31726
rect 51772 30818 51828 30828
rect 50876 29986 51268 29988
rect 50876 29934 51214 29986
rect 51266 29934 51268 29986
rect 50876 29932 51268 29934
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 50428 28644 50484 28654
rect 50428 28550 50484 28588
rect 50876 28644 50932 28654
rect 50316 28364 50484 28420
rect 50092 27682 50148 27692
rect 50428 27412 50484 28364
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 50652 27860 50708 27870
rect 50428 27356 50596 27412
rect 50428 27188 50484 27198
rect 50428 27094 50484 27132
rect 50540 26964 50596 27356
rect 50652 27300 50708 27804
rect 50652 27168 50708 27244
rect 50876 27186 50932 28588
rect 51100 27860 51156 27898
rect 51100 27794 51156 27804
rect 50876 27134 50878 27186
rect 50930 27134 50932 27186
rect 50876 27122 50932 27134
rect 51100 27636 51156 27646
rect 51100 27074 51156 27580
rect 51212 27524 51268 29932
rect 51324 30660 51380 30670
rect 51324 28084 51380 30604
rect 51324 28028 51492 28084
rect 51212 27458 51268 27468
rect 51212 27188 51268 27198
rect 51212 27094 51268 27132
rect 51100 27022 51102 27074
rect 51154 27022 51156 27074
rect 51100 27010 51156 27022
rect 49756 26850 49924 26852
rect 49756 26798 49758 26850
rect 49810 26798 49924 26850
rect 49756 26796 49924 26798
rect 49756 26786 49812 26796
rect 49868 26180 49924 26796
rect 50428 26908 50540 26964
rect 50428 26514 50484 26908
rect 50540 26832 50596 26908
rect 51324 26964 51380 26974
rect 51324 26870 51380 26908
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 50428 26462 50430 26514
rect 50482 26462 50484 26514
rect 50428 26450 50484 26462
rect 49868 26086 49924 26124
rect 50540 26180 50596 26190
rect 49532 25900 49924 25956
rect 49420 25442 49476 25452
rect 49756 25394 49812 25406
rect 49756 25342 49758 25394
rect 49810 25342 49812 25394
rect 49756 24724 49812 25342
rect 49868 24724 49924 25900
rect 50540 25620 50596 26124
rect 50540 25506 50596 25564
rect 51324 25620 51380 25630
rect 51324 25526 51380 25564
rect 50540 25454 50542 25506
rect 50594 25454 50596 25506
rect 50540 25442 50596 25454
rect 50764 25508 50820 25518
rect 50764 25414 50820 25452
rect 50316 25396 50372 25406
rect 50092 25394 50372 25396
rect 50092 25342 50318 25394
rect 50370 25342 50372 25394
rect 50092 25340 50372 25342
rect 49980 24948 50036 24958
rect 49980 24854 50036 24892
rect 50092 24946 50148 25340
rect 50316 25330 50372 25340
rect 50876 25396 50932 25406
rect 50876 25302 50932 25340
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 50092 24894 50094 24946
rect 50146 24894 50148 24946
rect 50092 24882 50148 24894
rect 49868 24668 50372 24724
rect 49756 24500 49812 24668
rect 50204 24500 50260 24510
rect 49756 24498 50260 24500
rect 49756 24446 50206 24498
rect 50258 24446 50260 24498
rect 49756 24444 50260 24446
rect 50204 23938 50260 24444
rect 50204 23886 50206 23938
rect 50258 23886 50260 23938
rect 50204 23874 50260 23886
rect 49308 23314 49364 23324
rect 49196 20692 49252 22988
rect 49308 21700 49364 21710
rect 49308 20914 49364 21644
rect 49644 21700 49700 21710
rect 49644 21586 49700 21644
rect 49644 21534 49646 21586
rect 49698 21534 49700 21586
rect 49644 21364 49700 21534
rect 49868 21588 49924 21598
rect 49868 21494 49924 21532
rect 49644 21298 49700 21308
rect 49308 20862 49310 20914
rect 49362 20862 49364 20914
rect 49308 20850 49364 20862
rect 49196 20636 49364 20692
rect 49084 19236 49140 19246
rect 49084 19142 49140 19180
rect 49196 19124 49252 19134
rect 49196 19030 49252 19068
rect 48972 18284 49140 18340
rect 48972 17892 49028 17902
rect 48972 17798 49028 17836
rect 48748 17714 48804 17724
rect 48860 17668 48916 17678
rect 48860 17574 48916 17612
rect 48076 17490 48132 17500
rect 48972 17556 49028 17566
rect 48972 17462 49028 17500
rect 48636 15876 48692 15886
rect 48636 15538 48692 15820
rect 48636 15486 48638 15538
rect 48690 15486 48692 15538
rect 48636 15474 48692 15486
rect 49084 15316 49140 18284
rect 48636 15260 49140 15316
rect 49196 15876 49252 15886
rect 49308 15876 49364 20636
rect 50316 20132 50372 24668
rect 50652 23826 50708 23838
rect 50652 23774 50654 23826
rect 50706 23774 50708 23826
rect 50652 23716 50708 23774
rect 50652 23660 50932 23716
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 50876 23156 50932 23660
rect 51100 23266 51156 23278
rect 51100 23214 51102 23266
rect 51154 23214 51156 23266
rect 50988 23156 51044 23166
rect 50876 23154 51044 23156
rect 50876 23102 50990 23154
rect 51042 23102 51044 23154
rect 50876 23100 51044 23102
rect 50540 22372 50596 22382
rect 50540 22278 50596 22316
rect 50988 22370 51044 23100
rect 50988 22318 50990 22370
rect 51042 22318 51044 22370
rect 50988 22306 51044 22318
rect 51100 22372 51156 23214
rect 51324 23268 51380 23278
rect 51324 23174 51380 23212
rect 51100 22306 51156 22316
rect 51212 22260 51268 22270
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 50540 21700 50596 21710
rect 50540 20914 50596 21644
rect 51100 21588 51156 21598
rect 51100 21494 51156 21532
rect 50540 20862 50542 20914
rect 50594 20862 50596 20914
rect 50540 20850 50596 20862
rect 50876 20804 50932 20814
rect 51212 20804 51268 22204
rect 51324 21364 51380 21374
rect 51324 21270 51380 21308
rect 50876 20802 51268 20804
rect 50876 20750 50878 20802
rect 50930 20750 51268 20802
rect 50876 20748 51268 20750
rect 50876 20738 50932 20748
rect 51324 20690 51380 20702
rect 51324 20638 51326 20690
rect 51378 20638 51380 20690
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 50316 20066 50372 20076
rect 49420 19236 49476 19246
rect 49868 19236 49924 19246
rect 49420 19234 49924 19236
rect 49420 19182 49422 19234
rect 49474 19182 49870 19234
rect 49922 19182 49924 19234
rect 49420 19180 49924 19182
rect 49420 19170 49476 19180
rect 49868 19170 49924 19180
rect 50092 19236 50148 19246
rect 49980 19124 50036 19134
rect 49980 18450 50036 19068
rect 49980 18398 49982 18450
rect 50034 18398 50036 18450
rect 49980 18386 50036 18398
rect 50092 18338 50148 19180
rect 51324 19122 51380 20638
rect 51436 19236 51492 28028
rect 51772 27748 51828 27758
rect 51772 27654 51828 27692
rect 51772 27524 51828 27534
rect 51772 24612 51828 27468
rect 51884 24836 51940 34636
rect 51996 34242 52052 34748
rect 51996 34190 51998 34242
rect 52050 34190 52052 34242
rect 52108 34356 52164 34860
rect 52108 34224 52164 34300
rect 52332 34354 52388 36428
rect 53340 36418 53396 36428
rect 53452 36260 53508 40348
rect 53564 40338 53620 40348
rect 53900 39618 53956 39630
rect 53900 39566 53902 39618
rect 53954 39566 53956 39618
rect 53564 39508 53620 39518
rect 53564 38948 53620 39452
rect 53564 38882 53620 38892
rect 53676 39394 53732 39406
rect 53676 39342 53678 39394
rect 53730 39342 53732 39394
rect 53676 38164 53732 39342
rect 53564 38108 53732 38164
rect 53788 38834 53844 38846
rect 53788 38782 53790 38834
rect 53842 38782 53844 38834
rect 53564 38050 53620 38108
rect 53564 37998 53566 38050
rect 53618 37998 53620 38050
rect 53564 37986 53620 37998
rect 53676 37940 53732 37950
rect 53788 37940 53844 38782
rect 53900 38724 53956 39566
rect 53900 38630 53956 38668
rect 53900 38164 53956 38174
rect 54012 38164 54068 41468
rect 54236 41458 54292 41468
rect 54348 41748 54404 41758
rect 54348 41410 54404 41692
rect 54348 41358 54350 41410
rect 54402 41358 54404 41410
rect 54348 41346 54404 41358
rect 54460 41746 54516 41758
rect 54460 41694 54462 41746
rect 54514 41694 54516 41746
rect 54460 41300 54516 41694
rect 54572 41748 54628 41758
rect 54572 41654 54628 41692
rect 54684 41410 54740 42028
rect 54684 41358 54686 41410
rect 54738 41358 54740 41410
rect 54684 41346 54740 41358
rect 55020 42530 55188 42532
rect 55020 42478 55134 42530
rect 55186 42478 55188 42530
rect 55020 42476 55188 42478
rect 54460 41234 54516 41244
rect 54908 41300 54964 41310
rect 55020 41300 55076 42476
rect 55132 42466 55188 42476
rect 55468 42532 55524 42542
rect 54908 41298 55076 41300
rect 54908 41246 54910 41298
rect 54962 41246 55076 41298
rect 54908 41244 55076 41246
rect 54908 41234 54964 41244
rect 54124 41186 54180 41198
rect 54124 41134 54126 41186
rect 54178 41134 54180 41186
rect 54124 40626 54180 41134
rect 54124 40574 54126 40626
rect 54178 40574 54180 40626
rect 54124 40562 54180 40574
rect 54460 40964 54516 40974
rect 54460 40626 54516 40908
rect 55020 40964 55076 41244
rect 55356 41300 55412 41310
rect 55468 41300 55524 42476
rect 55916 42532 55972 42542
rect 55916 42196 55972 42476
rect 55916 41746 55972 42140
rect 56028 41972 56084 43486
rect 56140 43538 56308 43540
rect 56140 43486 56254 43538
rect 56306 43486 56308 43538
rect 56140 43484 56308 43486
rect 56140 42532 56196 43484
rect 56252 43474 56308 43484
rect 56476 43540 56532 45164
rect 56588 44882 56644 44894
rect 56588 44830 56590 44882
rect 56642 44830 56644 44882
rect 56588 44434 56644 44830
rect 56588 44382 56590 44434
rect 56642 44382 56644 44434
rect 56700 44548 56756 45164
rect 56700 44416 56756 44492
rect 56588 43764 56644 44382
rect 56588 43698 56644 43708
rect 56812 44322 56868 44334
rect 56812 44270 56814 44322
rect 56866 44270 56868 44322
rect 56476 43446 56532 43484
rect 56812 43540 56868 44270
rect 56812 43474 56868 43484
rect 56476 42980 56532 42990
rect 56924 42980 56980 46508
rect 57372 47460 57428 49756
rect 57484 49746 57540 49756
rect 57596 49026 57652 49038
rect 57596 48974 57598 49026
rect 57650 48974 57652 49026
rect 57484 48804 57540 48814
rect 57596 48804 57652 48974
rect 57820 49026 57876 49982
rect 57820 48974 57822 49026
rect 57874 48974 57876 49026
rect 57820 48962 57876 48974
rect 58156 50370 58212 50382
rect 58156 50318 58158 50370
rect 58210 50318 58212 50370
rect 58156 49810 58212 50318
rect 58268 49924 58324 51212
rect 58380 51266 58660 51268
rect 58380 51214 58382 51266
rect 58434 51214 58660 51266
rect 58380 51212 58660 51214
rect 58380 51154 58436 51212
rect 58380 51102 58382 51154
rect 58434 51102 58436 51154
rect 58380 51090 58436 51102
rect 58380 49924 58436 49934
rect 58268 49922 58436 49924
rect 58268 49870 58382 49922
rect 58434 49870 58436 49922
rect 58268 49868 58436 49870
rect 58156 49758 58158 49810
rect 58210 49758 58212 49810
rect 58156 48804 58212 49758
rect 58268 49028 58324 49038
rect 58268 48934 58324 48972
rect 57596 48748 58212 48804
rect 57484 48354 57540 48748
rect 57484 48302 57486 48354
rect 57538 48302 57540 48354
rect 57484 48290 57540 48302
rect 57596 48242 57652 48254
rect 57596 48190 57598 48242
rect 57650 48190 57652 48242
rect 57596 47796 57652 48190
rect 57932 48244 57988 48254
rect 57932 48150 57988 48188
rect 58380 48244 58436 49868
rect 58492 49924 58548 49934
rect 58492 49830 58548 49868
rect 58380 48178 58436 48188
rect 57596 47730 57652 47740
rect 57372 46116 57428 47404
rect 57484 47236 57540 47246
rect 57484 46786 57540 47180
rect 57484 46734 57486 46786
rect 57538 46734 57540 46786
rect 57484 46722 57540 46734
rect 58156 46674 58212 46686
rect 58156 46622 58158 46674
rect 58210 46622 58212 46674
rect 57820 46562 57876 46574
rect 57820 46510 57822 46562
rect 57874 46510 57876 46562
rect 57484 46116 57540 46126
rect 57372 46114 57540 46116
rect 57372 46062 57486 46114
rect 57538 46062 57540 46114
rect 57372 46060 57540 46062
rect 57484 46050 57540 46060
rect 57820 46114 57876 46510
rect 57820 46062 57822 46114
rect 57874 46062 57876 46114
rect 56140 42438 56196 42476
rect 56252 42642 56308 42654
rect 56252 42590 56254 42642
rect 56306 42590 56308 42642
rect 56252 41972 56308 42590
rect 56028 41916 56308 41972
rect 55916 41694 55918 41746
rect 55970 41694 55972 41746
rect 55916 41682 55972 41694
rect 56252 41858 56308 41916
rect 56364 42532 56420 42542
rect 56364 42084 56420 42476
rect 56364 41970 56420 42028
rect 56364 41918 56366 41970
rect 56418 41918 56420 41970
rect 56364 41906 56420 41918
rect 56252 41806 56254 41858
rect 56306 41806 56308 41858
rect 55356 41298 55524 41300
rect 55356 41246 55358 41298
rect 55410 41246 55524 41298
rect 55356 41244 55524 41246
rect 55356 41234 55412 41244
rect 55020 40898 55076 40908
rect 55804 40964 55860 40974
rect 55804 40870 55860 40908
rect 54460 40574 54462 40626
rect 54514 40574 54516 40626
rect 54460 40562 54516 40574
rect 54684 39508 54740 39518
rect 54348 39396 54404 39406
rect 53900 38162 54068 38164
rect 53900 38110 53902 38162
rect 53954 38110 54068 38162
rect 53900 38108 54068 38110
rect 54124 39394 54404 39396
rect 54124 39342 54350 39394
rect 54402 39342 54404 39394
rect 54124 39340 54404 39342
rect 53900 38098 53956 38108
rect 54124 38050 54180 39340
rect 54348 39330 54404 39340
rect 54572 39394 54628 39406
rect 54572 39342 54574 39394
rect 54626 39342 54628 39394
rect 54572 38724 54628 39342
rect 54684 38836 54740 39452
rect 54796 38836 54852 38846
rect 54684 38834 54852 38836
rect 54684 38782 54798 38834
rect 54850 38782 54852 38834
rect 54684 38780 54852 38782
rect 54796 38770 54852 38780
rect 54572 38500 54628 38668
rect 55580 38724 55636 38734
rect 55580 38630 55636 38668
rect 54572 38444 55076 38500
rect 54124 37998 54126 38050
rect 54178 37998 54180 38050
rect 54124 37986 54180 37998
rect 53676 37938 53844 37940
rect 53676 37886 53678 37938
rect 53730 37886 53844 37938
rect 53676 37884 53844 37886
rect 53676 37874 53732 37884
rect 53788 36596 53844 37884
rect 54908 37940 54964 37950
rect 54348 37492 54404 37502
rect 54348 37398 54404 37436
rect 54908 37490 54964 37884
rect 54908 37438 54910 37490
rect 54962 37438 54964 37490
rect 54908 37426 54964 37438
rect 53900 36596 53956 36606
rect 53788 36594 53956 36596
rect 53788 36542 53902 36594
rect 53954 36542 53956 36594
rect 53788 36540 53956 36542
rect 53900 36530 53956 36540
rect 55020 36594 55076 38444
rect 55244 38162 55300 38174
rect 55244 38110 55246 38162
rect 55298 38110 55300 38162
rect 55244 37492 55300 38110
rect 56252 38164 56308 41806
rect 56476 39058 56532 42924
rect 56700 42924 56980 42980
rect 57036 46004 57092 46014
rect 56700 42866 56756 42924
rect 56700 42814 56702 42866
rect 56754 42814 56756 42866
rect 56700 42196 56756 42814
rect 56700 42130 56756 42140
rect 57036 42532 57092 45948
rect 57820 45332 57876 46062
rect 58044 45892 58100 45902
rect 58156 45892 58212 46622
rect 58044 45890 58212 45892
rect 58044 45838 58046 45890
rect 58098 45838 58212 45890
rect 58044 45836 58212 45838
rect 58044 45826 58100 45836
rect 57932 45332 57988 45342
rect 57820 45330 57988 45332
rect 57820 45278 57934 45330
rect 57986 45278 57988 45330
rect 57820 45276 57988 45278
rect 57932 45266 57988 45276
rect 57596 45218 57652 45230
rect 57596 45166 57598 45218
rect 57650 45166 57652 45218
rect 57484 43764 57540 43774
rect 57484 43650 57540 43708
rect 57484 43598 57486 43650
rect 57538 43598 57540 43650
rect 57484 43586 57540 43598
rect 57260 43540 57316 43550
rect 57148 42532 57204 42542
rect 57036 42530 57204 42532
rect 57036 42478 57150 42530
rect 57202 42478 57204 42530
rect 57036 42476 57204 42478
rect 56588 41412 56644 41422
rect 56588 41298 56644 41356
rect 56588 41246 56590 41298
rect 56642 41246 56644 41298
rect 56588 41234 56644 41246
rect 57036 40964 57092 42476
rect 57148 42466 57204 42476
rect 57260 41298 57316 43484
rect 57596 42756 57652 45166
rect 57820 45108 57876 45118
rect 57708 45052 57820 45108
rect 57708 44436 57764 45052
rect 57820 44976 57876 45052
rect 58044 45106 58100 45118
rect 58044 45054 58046 45106
rect 58098 45054 58100 45106
rect 57708 43708 57764 44380
rect 57708 43652 57988 43708
rect 57932 43538 57988 43652
rect 57932 43486 57934 43538
rect 57986 43486 57988 43538
rect 57932 43474 57988 43486
rect 58044 43428 58100 45054
rect 58156 43708 58212 45836
rect 58492 45108 58548 45118
rect 58492 45014 58548 45052
rect 58156 43652 58548 43708
rect 58380 43428 58436 43438
rect 58044 43426 58436 43428
rect 58044 43374 58382 43426
rect 58434 43374 58436 43426
rect 58044 43372 58436 43374
rect 57596 42700 57876 42756
rect 57596 42532 57652 42542
rect 57260 41246 57262 41298
rect 57314 41246 57316 41298
rect 57260 41234 57316 41246
rect 57372 42530 57652 42532
rect 57372 42478 57598 42530
rect 57650 42478 57652 42530
rect 57372 42476 57652 42478
rect 57372 41412 57428 42476
rect 57596 42466 57652 42476
rect 57484 42084 57540 42094
rect 57484 41990 57540 42028
rect 56812 39620 56868 39630
rect 56588 39396 56644 39406
rect 56812 39396 56868 39564
rect 56588 39394 56868 39396
rect 56588 39342 56590 39394
rect 56642 39342 56868 39394
rect 56588 39340 56868 39342
rect 56588 39330 56644 39340
rect 56476 39006 56478 39058
rect 56530 39006 56532 39058
rect 56476 38994 56532 39006
rect 56700 38836 56756 38846
rect 56700 38742 56756 38780
rect 56364 38724 56420 38734
rect 56364 38630 56420 38668
rect 56364 38164 56420 38174
rect 56252 38162 56420 38164
rect 56252 38110 56366 38162
rect 56418 38110 56420 38162
rect 56252 38108 56420 38110
rect 56364 38098 56420 38108
rect 55244 37426 55300 37436
rect 56140 38050 56196 38062
rect 56140 37998 56142 38050
rect 56194 37998 56196 38050
rect 55916 37044 55972 37054
rect 55020 36542 55022 36594
rect 55074 36542 55076 36594
rect 55020 36530 55076 36542
rect 55468 37042 55972 37044
rect 55468 36990 55918 37042
rect 55970 36990 55972 37042
rect 55468 36988 55972 36990
rect 54572 36372 54628 36382
rect 54124 36370 54628 36372
rect 54124 36318 54574 36370
rect 54626 36318 54628 36370
rect 54124 36316 54628 36318
rect 53116 36204 53508 36260
rect 53788 36258 53844 36270
rect 53788 36206 53790 36258
rect 53842 36206 53844 36258
rect 53004 35700 53060 35710
rect 53004 35606 53060 35644
rect 52556 34916 52612 34926
rect 52556 34822 52612 34860
rect 52332 34302 52334 34354
rect 52386 34302 52388 34354
rect 52332 34290 52388 34302
rect 52668 34356 52724 34366
rect 52668 34262 52724 34300
rect 51996 34178 52052 34190
rect 53116 31948 53172 36204
rect 53228 35698 53284 35710
rect 53228 35646 53230 35698
rect 53282 35646 53284 35698
rect 53228 35252 53284 35646
rect 53676 35700 53732 35710
rect 53284 35196 53508 35252
rect 53228 35186 53284 35196
rect 53452 34130 53508 35196
rect 53564 34916 53620 34926
rect 53564 34822 53620 34860
rect 53452 34078 53454 34130
rect 53506 34078 53508 34130
rect 53452 34066 53508 34078
rect 53676 34130 53732 35644
rect 53788 34914 53844 36206
rect 54012 36258 54068 36270
rect 54012 36206 54014 36258
rect 54066 36206 54068 36258
rect 53900 35812 53956 35822
rect 53900 35718 53956 35756
rect 53788 34862 53790 34914
rect 53842 34862 53844 34914
rect 53788 34804 53844 34862
rect 54012 34916 54068 36206
rect 54012 34850 54068 34860
rect 53788 34738 53844 34748
rect 54012 34356 54068 34366
rect 54124 34356 54180 36316
rect 54572 36306 54628 36316
rect 54796 36370 54852 36382
rect 54796 36318 54798 36370
rect 54850 36318 54852 36370
rect 54796 35812 54852 36318
rect 54796 35698 54852 35756
rect 54796 35646 54798 35698
rect 54850 35646 54852 35698
rect 54796 35634 54852 35646
rect 55132 36370 55188 36382
rect 55132 36318 55134 36370
rect 55186 36318 55188 36370
rect 54684 35586 54740 35598
rect 54684 35534 54686 35586
rect 54738 35534 54740 35586
rect 54684 35476 54740 35534
rect 55132 35476 55188 36318
rect 54684 35420 55188 35476
rect 55468 35476 55524 36988
rect 55916 36978 55972 36988
rect 56140 36820 56196 37998
rect 56476 38050 56532 38062
rect 56476 37998 56478 38050
rect 56530 37998 56532 38050
rect 56364 37156 56420 37166
rect 56476 37156 56532 37998
rect 56364 37154 56532 37156
rect 56364 37102 56366 37154
rect 56418 37102 56532 37154
rect 56364 37100 56532 37102
rect 56700 37154 56756 37166
rect 56700 37102 56702 37154
rect 56754 37102 56756 37154
rect 56364 37042 56420 37100
rect 56364 36990 56366 37042
rect 56418 36990 56420 37042
rect 56364 36978 56420 36990
rect 56700 36820 56756 37102
rect 55692 36764 56756 36820
rect 55580 35700 55636 35710
rect 55580 35606 55636 35644
rect 55468 35420 55636 35476
rect 54460 35028 54516 35038
rect 54684 35028 54740 35420
rect 54460 35026 54740 35028
rect 54460 34974 54462 35026
rect 54514 34974 54740 35026
rect 54460 34972 54740 34974
rect 54460 34962 54516 34972
rect 54012 34354 54180 34356
rect 54012 34302 54014 34354
rect 54066 34302 54180 34354
rect 54012 34300 54180 34302
rect 54012 34290 54068 34300
rect 53676 34078 53678 34130
rect 53730 34078 53732 34130
rect 53676 34066 53732 34078
rect 54460 33460 54516 33470
rect 54460 32674 54516 33404
rect 54460 32622 54462 32674
rect 54514 32622 54516 32674
rect 54460 32610 54516 32622
rect 54796 33122 54852 33134
rect 54796 33070 54798 33122
rect 54850 33070 54852 33122
rect 53788 32562 53844 32574
rect 53788 32510 53790 32562
rect 53842 32510 53844 32562
rect 53116 31892 53284 31948
rect 52444 31778 52500 31790
rect 52444 31726 52446 31778
rect 52498 31726 52500 31778
rect 52444 31108 52500 31726
rect 52668 31668 52724 31678
rect 52668 31574 52724 31612
rect 52780 31220 52836 31230
rect 52780 31126 52836 31164
rect 52444 30976 52500 31052
rect 52556 31106 52612 31118
rect 52556 31054 52558 31106
rect 52610 31054 52612 31106
rect 52556 30884 52612 31054
rect 52556 30818 52612 30828
rect 52668 30996 52724 31006
rect 52668 30212 52724 30940
rect 53116 30884 53172 30894
rect 53116 30790 53172 30828
rect 52108 30100 52164 30110
rect 52668 30080 52724 30156
rect 52108 29428 52164 30044
rect 53004 29540 53060 29550
rect 53004 29446 53060 29484
rect 52108 29426 52276 29428
rect 52108 29374 52110 29426
rect 52162 29374 52276 29426
rect 52108 29372 52276 29374
rect 52108 29362 52164 29372
rect 52220 28868 52276 29372
rect 52444 29426 52500 29438
rect 52444 29374 52446 29426
rect 52498 29374 52500 29426
rect 52332 28868 52388 28878
rect 52220 28866 52388 28868
rect 52220 28814 52334 28866
rect 52386 28814 52388 28866
rect 52220 28812 52388 28814
rect 52332 28802 52388 28812
rect 52108 28644 52164 28654
rect 52444 28644 52500 29374
rect 52668 28868 52724 28878
rect 52668 28774 52724 28812
rect 52164 28588 52500 28644
rect 52108 28512 52164 28588
rect 52668 27858 52724 27870
rect 52668 27806 52670 27858
rect 52722 27806 52724 27858
rect 52444 27748 52500 27758
rect 52444 27654 52500 27692
rect 52108 27076 52164 27086
rect 51996 26964 52052 26974
rect 51996 26870 52052 26908
rect 52108 26514 52164 27020
rect 52668 26964 52724 27806
rect 52668 26898 52724 26908
rect 52780 27076 52836 27086
rect 52108 26462 52110 26514
rect 52162 26462 52164 26514
rect 52108 26450 52164 26462
rect 52780 26292 52836 27020
rect 52892 26292 52948 26302
rect 52780 26290 52948 26292
rect 52780 26238 52894 26290
rect 52946 26238 52948 26290
rect 52780 26236 52948 26238
rect 52892 26226 52948 26236
rect 51884 24770 51940 24780
rect 52780 25284 52836 25294
rect 52780 24834 52836 25228
rect 53228 24836 53284 31892
rect 53340 31778 53396 31790
rect 53340 31726 53342 31778
rect 53394 31726 53396 31778
rect 53340 31220 53396 31726
rect 53340 31154 53396 31164
rect 53788 31554 53844 32510
rect 54796 32564 54852 33070
rect 54796 32498 54852 32508
rect 55356 32564 55412 32574
rect 54012 32450 54068 32462
rect 54012 32398 54014 32450
rect 54066 32398 54068 32450
rect 53900 32004 53956 32014
rect 53900 31890 53956 31948
rect 53900 31838 53902 31890
rect 53954 31838 53956 31890
rect 53900 31826 53956 31838
rect 54012 31668 54068 32398
rect 55132 32450 55188 32462
rect 55132 32398 55134 32450
rect 55186 32398 55188 32450
rect 54460 31892 54516 31902
rect 54460 31798 54516 31836
rect 54796 31892 54852 31902
rect 54012 31574 54068 31612
rect 53788 31502 53790 31554
rect 53842 31502 53844 31554
rect 53676 30212 53732 30222
rect 53452 30098 53508 30110
rect 53452 30046 53454 30098
rect 53506 30046 53508 30098
rect 53452 28868 53508 30046
rect 53676 29428 53732 30156
rect 53788 29986 53844 31502
rect 54796 31218 54852 31836
rect 55132 31892 55188 32398
rect 55356 31948 55412 32508
rect 55132 31826 55188 31836
rect 55244 31892 55412 31948
rect 55468 31892 55524 31902
rect 54796 31166 54798 31218
rect 54850 31166 54852 31218
rect 54796 31154 54852 31166
rect 55244 31778 55300 31892
rect 55468 31798 55524 31836
rect 55244 31726 55246 31778
rect 55298 31726 55300 31778
rect 55244 31556 55300 31726
rect 55244 31218 55300 31500
rect 55244 31166 55246 31218
rect 55298 31166 55300 31218
rect 55244 31154 55300 31166
rect 53788 29934 53790 29986
rect 53842 29934 53844 29986
rect 53788 29922 53844 29934
rect 54124 30210 54180 30222
rect 54124 30158 54126 30210
rect 54178 30158 54180 30210
rect 54124 29540 54180 30158
rect 53900 29428 53956 29438
rect 53452 28802 53508 28812
rect 53564 29426 53956 29428
rect 53564 29374 53902 29426
rect 53954 29374 53956 29426
rect 53564 29372 53956 29374
rect 53564 28756 53620 29372
rect 53900 29362 53956 29372
rect 54124 29314 54180 29484
rect 54908 30212 54964 30222
rect 54908 29986 54964 30156
rect 55468 30212 55524 30222
rect 55468 30118 55524 30156
rect 54908 29934 54910 29986
rect 54962 29934 54964 29986
rect 54124 29262 54126 29314
rect 54178 29262 54180 29314
rect 54124 29250 54180 29262
rect 54572 29316 54628 29326
rect 54908 29316 54964 29934
rect 55132 29316 55188 29326
rect 54908 29314 55188 29316
rect 54908 29262 55134 29314
rect 55186 29262 55188 29314
rect 54908 29260 55188 29262
rect 54572 29222 54628 29260
rect 53340 28644 53396 28654
rect 53564 28644 53620 28700
rect 54348 29092 54404 29102
rect 54348 28754 54404 29036
rect 54348 28702 54350 28754
rect 54402 28702 54404 28754
rect 54348 28690 54404 28702
rect 55132 29092 55188 29260
rect 55132 28754 55188 29036
rect 55132 28702 55134 28754
rect 55186 28702 55188 28754
rect 55132 28690 55188 28702
rect 55356 29316 55412 29326
rect 53340 28642 53620 28644
rect 53340 28590 53342 28642
rect 53394 28590 53620 28642
rect 53340 28588 53620 28590
rect 55020 28642 55076 28654
rect 55020 28590 55022 28642
rect 55074 28590 55076 28642
rect 53340 28578 53396 28588
rect 55020 28532 55076 28590
rect 55356 28644 55412 29260
rect 55356 28578 55412 28588
rect 53340 27748 53396 27758
rect 53340 27746 53508 27748
rect 53340 27694 53342 27746
rect 53394 27694 53508 27746
rect 53340 27692 53508 27694
rect 53340 27682 53396 27692
rect 53452 26962 53508 27692
rect 55020 27188 55076 28476
rect 55020 27122 55076 27132
rect 53676 27076 53732 27114
rect 53676 27010 53732 27020
rect 53452 26910 53454 26962
rect 53506 26910 53508 26962
rect 53452 26178 53508 26910
rect 54012 26964 54068 26974
rect 54012 26962 54516 26964
rect 54012 26910 54014 26962
rect 54066 26910 54516 26962
rect 54012 26908 54516 26910
rect 54012 26898 54068 26908
rect 53676 26852 53732 26862
rect 53676 26758 53732 26796
rect 54460 26514 54516 26908
rect 54460 26462 54462 26514
rect 54514 26462 54516 26514
rect 54460 26450 54516 26462
rect 53452 26126 53454 26178
rect 53506 26126 53508 26178
rect 53452 26114 53508 26126
rect 54572 26402 54628 26414
rect 54572 26350 54574 26402
rect 54626 26350 54628 26402
rect 53676 26068 53732 26078
rect 53676 25974 53732 26012
rect 54348 26068 54404 26078
rect 54348 25618 54404 26012
rect 54348 25566 54350 25618
rect 54402 25566 54404 25618
rect 54348 25554 54404 25566
rect 53900 25508 53956 25518
rect 53900 25414 53956 25452
rect 54572 25508 54628 26350
rect 55580 26292 55636 35420
rect 55692 30436 55748 36764
rect 56252 35924 56308 35934
rect 55916 34130 55972 34142
rect 55916 34078 55918 34130
rect 55970 34078 55972 34130
rect 55804 31892 55860 31902
rect 55916 31892 55972 34078
rect 56140 34130 56196 34142
rect 56140 34078 56142 34130
rect 56194 34078 56196 34130
rect 56140 33348 56196 34078
rect 56252 34132 56308 35868
rect 56588 35810 56644 35822
rect 56588 35758 56590 35810
rect 56642 35758 56644 35810
rect 56364 35700 56420 35710
rect 56364 35476 56420 35644
rect 56364 35474 56532 35476
rect 56364 35422 56366 35474
rect 56418 35422 56532 35474
rect 56364 35420 56532 35422
rect 56364 35410 56420 35420
rect 56476 35026 56532 35420
rect 56476 34974 56478 35026
rect 56530 34974 56532 35026
rect 56476 34962 56532 34974
rect 56588 34916 56644 35758
rect 56700 35700 56756 35710
rect 56700 35586 56756 35644
rect 56700 35534 56702 35586
rect 56754 35534 56756 35586
rect 56700 35522 56756 35534
rect 56700 34916 56756 34926
rect 56588 34914 56756 34916
rect 56588 34862 56702 34914
rect 56754 34862 56756 34914
rect 56588 34860 56756 34862
rect 56364 34356 56420 34366
rect 56700 34356 56756 34860
rect 56364 34354 56756 34356
rect 56364 34302 56366 34354
rect 56418 34302 56756 34354
rect 56364 34300 56756 34302
rect 56364 34290 56420 34300
rect 56252 34076 56420 34132
rect 56252 33348 56308 33358
rect 56028 33346 56308 33348
rect 56028 33294 56254 33346
rect 56306 33294 56308 33346
rect 56028 33292 56308 33294
rect 56028 32674 56084 33292
rect 56252 33282 56308 33292
rect 56028 32622 56030 32674
rect 56082 32622 56084 32674
rect 56028 32610 56084 32622
rect 56364 31948 56420 34076
rect 56476 34130 56532 34142
rect 56476 34078 56478 34130
rect 56530 34078 56532 34130
rect 56476 33460 56532 34078
rect 56476 33366 56532 33404
rect 56812 31948 56868 39340
rect 56924 33234 56980 33246
rect 56924 33182 56926 33234
rect 56978 33182 56980 33234
rect 56924 32564 56980 33182
rect 56924 32498 56980 32508
rect 55804 31890 55972 31892
rect 55804 31838 55806 31890
rect 55858 31838 55972 31890
rect 55804 31836 55972 31838
rect 56252 31892 56420 31948
rect 56476 31892 56868 31948
rect 55804 31826 55860 31836
rect 55692 30380 55860 30436
rect 55692 30210 55748 30222
rect 55692 30158 55694 30210
rect 55746 30158 55748 30210
rect 55692 29428 55748 30158
rect 55692 29362 55748 29372
rect 55692 29204 55748 29214
rect 55692 29110 55748 29148
rect 54572 25442 54628 25452
rect 55468 26236 55636 26292
rect 53452 25396 53508 25406
rect 52780 24782 52782 24834
rect 52834 24782 52836 24834
rect 52780 24770 52836 24782
rect 53116 24780 53284 24836
rect 53340 25394 53508 25396
rect 53340 25342 53454 25394
rect 53506 25342 53508 25394
rect 53340 25340 53508 25342
rect 53004 24722 53060 24734
rect 53004 24670 53006 24722
rect 53058 24670 53060 24722
rect 51772 24556 51940 24612
rect 51772 22258 51828 22270
rect 51772 22206 51774 22258
rect 51826 22206 51828 22258
rect 51660 21812 51716 21822
rect 51772 21812 51828 22206
rect 51660 21810 51828 21812
rect 51660 21758 51662 21810
rect 51714 21758 51828 21810
rect 51660 21756 51828 21758
rect 51660 21746 51716 21756
rect 51884 20188 51940 24556
rect 52668 23828 52724 23838
rect 52668 23154 52724 23772
rect 53004 23828 53060 24670
rect 53116 24388 53172 24780
rect 53340 24722 53396 25340
rect 53452 25330 53508 25340
rect 53340 24670 53342 24722
rect 53394 24670 53396 24722
rect 53228 24612 53284 24622
rect 53228 24518 53284 24556
rect 53116 24332 53284 24388
rect 53004 23762 53060 23772
rect 52668 23102 52670 23154
rect 52722 23102 52724 23154
rect 52668 23090 52724 23102
rect 51996 22260 52052 22270
rect 51996 22166 52052 22204
rect 52220 22260 52276 22270
rect 52220 22166 52276 22204
rect 52332 22258 52388 22270
rect 52332 22206 52334 22258
rect 52386 22206 52388 22258
rect 52332 21700 52388 22206
rect 52332 21634 52388 21644
rect 52108 21474 52164 21486
rect 52108 21422 52110 21474
rect 52162 21422 52164 21474
rect 52108 21364 52164 21422
rect 52108 21298 52164 21308
rect 51884 20132 52276 20188
rect 51436 19170 51492 19180
rect 52220 19906 52276 20132
rect 52892 19908 52948 19918
rect 52220 19854 52222 19906
rect 52274 19854 52276 19906
rect 51324 19070 51326 19122
rect 51378 19070 51380 19122
rect 50316 19012 50372 19022
rect 50092 18286 50094 18338
rect 50146 18286 50148 18338
rect 50092 18274 50148 18286
rect 50204 19010 50372 19012
rect 50204 18958 50318 19010
rect 50370 18958 50372 19010
rect 50204 18956 50372 18958
rect 50092 17892 50148 17902
rect 50204 17892 50260 18956
rect 50316 18946 50372 18956
rect 50428 19012 50484 19022
rect 50428 18918 50484 18956
rect 50540 19012 50596 19022
rect 50540 19010 50932 19012
rect 50540 18958 50542 19010
rect 50594 18958 50932 19010
rect 50540 18956 50932 18958
rect 50540 18946 50596 18956
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 50092 17890 50260 17892
rect 50092 17838 50094 17890
rect 50146 17838 50260 17890
rect 50092 17836 50260 17838
rect 50316 18228 50372 18238
rect 50092 17826 50148 17836
rect 49980 17780 50036 17790
rect 49980 16884 50036 17724
rect 50092 16884 50148 16894
rect 49980 16882 50148 16884
rect 49980 16830 50094 16882
rect 50146 16830 50148 16882
rect 49980 16828 50148 16830
rect 50092 16818 50148 16828
rect 50316 16770 50372 18172
rect 50876 18228 50932 18956
rect 50876 18162 50932 18172
rect 51324 17778 51380 19070
rect 52220 19124 52276 19854
rect 52780 19852 52892 19908
rect 52220 19058 52276 19068
rect 52668 19124 52724 19134
rect 52668 19030 52724 19068
rect 51324 17726 51326 17778
rect 51378 17726 51380 17778
rect 51324 17714 51380 17726
rect 51436 19012 51492 19022
rect 51436 17666 51492 18956
rect 51660 19010 51716 19022
rect 51660 18958 51662 19010
rect 51714 18958 51716 19010
rect 51660 18450 51716 18958
rect 52780 18564 52836 19852
rect 52892 19776 52948 19852
rect 52780 18470 52836 18508
rect 51660 18398 51662 18450
rect 51714 18398 51716 18450
rect 51660 18386 51716 18398
rect 52108 18450 52164 18462
rect 52108 18398 52110 18450
rect 52162 18398 52164 18450
rect 52108 17892 52164 18398
rect 52108 17826 52164 17836
rect 52220 18338 52276 18350
rect 52220 18286 52222 18338
rect 52274 18286 52276 18338
rect 51436 17614 51438 17666
rect 51490 17614 51492 17666
rect 51436 17602 51492 17614
rect 51996 17668 52052 17678
rect 52220 17668 52276 18286
rect 51996 17666 52276 17668
rect 51996 17614 51998 17666
rect 52050 17614 52276 17666
rect 51996 17612 52276 17614
rect 52332 17892 52388 17902
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 51996 16882 52052 17612
rect 51996 16830 51998 16882
rect 52050 16830 52052 16882
rect 51996 16818 52052 16830
rect 52332 16882 52388 17836
rect 53228 17108 53284 24332
rect 53340 23154 53396 24670
rect 55132 24836 55188 24846
rect 54684 24050 54740 24062
rect 54684 23998 54686 24050
rect 54738 23998 54740 24050
rect 54124 23938 54180 23950
rect 54124 23886 54126 23938
rect 54178 23886 54180 23938
rect 54012 23268 54068 23278
rect 53340 23102 53342 23154
rect 53394 23102 53396 23154
rect 53340 23090 53396 23102
rect 53564 23156 53620 23166
rect 53452 23044 53508 23054
rect 53452 22950 53508 22988
rect 53564 22260 53620 23100
rect 53564 21698 53620 22204
rect 53564 21646 53566 21698
rect 53618 21646 53620 21698
rect 53564 21634 53620 21646
rect 53788 23044 53844 23054
rect 53788 21586 53844 22988
rect 54012 22370 54068 23212
rect 54012 22318 54014 22370
rect 54066 22318 54068 22370
rect 54012 22306 54068 22318
rect 54124 21810 54180 23886
rect 54460 23938 54516 23950
rect 54460 23886 54462 23938
rect 54514 23886 54516 23938
rect 54460 23268 54516 23886
rect 54460 23202 54516 23212
rect 54348 23156 54404 23166
rect 54348 23062 54404 23100
rect 54460 23044 54516 23054
rect 54460 22950 54516 22988
rect 54684 22930 54740 23998
rect 55132 23828 55188 24780
rect 55468 24500 55524 26236
rect 55804 25618 55860 30380
rect 56028 29986 56084 29998
rect 56028 29934 56030 29986
rect 56082 29934 56084 29986
rect 56028 29540 56084 29934
rect 56028 29474 56084 29484
rect 56140 29314 56196 29326
rect 56140 29262 56142 29314
rect 56194 29262 56196 29314
rect 56140 29092 56196 29262
rect 56140 29026 56196 29036
rect 56252 26628 56308 31892
rect 56364 30882 56420 30894
rect 56364 30830 56366 30882
rect 56418 30830 56420 30882
rect 56364 28980 56420 30830
rect 56476 29092 56532 31892
rect 56812 30882 56868 30894
rect 56812 30830 56814 30882
rect 56866 30830 56868 30882
rect 56588 30772 56644 30782
rect 56588 30322 56644 30716
rect 56812 30772 56868 30830
rect 56812 30706 56868 30716
rect 56588 30270 56590 30322
rect 56642 30270 56644 30322
rect 56588 30258 56644 30270
rect 56700 29314 56756 29326
rect 56700 29262 56702 29314
rect 56754 29262 56756 29314
rect 56476 29036 56644 29092
rect 56364 28914 56420 28924
rect 56364 28644 56420 28654
rect 56364 28550 56420 28588
rect 55804 25566 55806 25618
rect 55858 25566 55860 25618
rect 55804 25554 55860 25566
rect 56140 26572 56308 26628
rect 56476 26852 56532 26862
rect 55692 25508 55748 25518
rect 55580 25506 55748 25508
rect 55580 25454 55694 25506
rect 55746 25454 55748 25506
rect 55580 25452 55748 25454
rect 55580 24836 55636 25452
rect 55692 25442 55748 25452
rect 56028 25396 56084 25406
rect 55804 25340 56028 25396
rect 55580 24742 55636 24780
rect 55692 24836 55748 24846
rect 55804 24836 55860 25340
rect 56028 25302 56084 25340
rect 55692 24834 55860 24836
rect 55692 24782 55694 24834
rect 55746 24782 55860 24834
rect 55692 24780 55860 24782
rect 55692 24770 55748 24780
rect 55580 24500 55636 24510
rect 55468 24498 55636 24500
rect 55468 24446 55582 24498
rect 55634 24446 55636 24498
rect 55468 24444 55636 24446
rect 55580 24434 55636 24444
rect 55132 23734 55188 23772
rect 56140 23826 56196 26572
rect 56476 26514 56532 26796
rect 56476 26462 56478 26514
rect 56530 26462 56532 26514
rect 56476 26450 56532 26462
rect 56588 26514 56644 29036
rect 56700 28980 56756 29262
rect 56700 28914 56756 28924
rect 56588 26462 56590 26514
rect 56642 26462 56644 26514
rect 56588 26450 56644 26462
rect 56252 26402 56308 26414
rect 56252 26350 56254 26402
rect 56306 26350 56308 26402
rect 56252 24948 56308 26350
rect 56700 26292 56756 26302
rect 56700 26198 56756 26236
rect 56924 26292 56980 26302
rect 56924 25506 56980 26236
rect 56924 25454 56926 25506
rect 56978 25454 56980 25506
rect 56924 25442 56980 25454
rect 57036 25172 57092 40908
rect 57148 41188 57204 41198
rect 57148 39618 57204 41132
rect 57372 41186 57428 41356
rect 57372 41134 57374 41186
rect 57426 41134 57428 41186
rect 57372 41122 57428 41134
rect 57596 41970 57652 41982
rect 57596 41918 57598 41970
rect 57650 41918 57652 41970
rect 57596 41188 57652 41918
rect 57596 41122 57652 41132
rect 57596 40962 57652 40974
rect 57596 40910 57598 40962
rect 57650 40910 57652 40962
rect 57484 40628 57540 40638
rect 57596 40628 57652 40910
rect 57484 40626 57652 40628
rect 57484 40574 57486 40626
rect 57538 40574 57652 40626
rect 57484 40572 57652 40574
rect 57820 40628 57876 42700
rect 57932 41970 57988 41982
rect 57932 41918 57934 41970
rect 57986 41918 57988 41970
rect 57932 41412 57988 41918
rect 57932 41346 57988 41356
rect 57820 40572 57988 40628
rect 57484 40562 57540 40572
rect 57708 40516 57764 40526
rect 57708 40422 57764 40460
rect 57820 40402 57876 40414
rect 57820 40350 57822 40402
rect 57874 40350 57876 40402
rect 57820 40292 57876 40350
rect 57596 40236 57876 40292
rect 57372 39620 57428 39630
rect 57596 39620 57652 40236
rect 57932 40180 57988 40572
rect 57148 39566 57150 39618
rect 57202 39566 57204 39618
rect 57148 39554 57204 39566
rect 57260 39618 57652 39620
rect 57260 39566 57374 39618
rect 57426 39566 57652 39618
rect 57260 39564 57652 39566
rect 57708 40124 57988 40180
rect 58268 40514 58324 40526
rect 58268 40462 58270 40514
rect 58322 40462 58324 40514
rect 58268 40292 58324 40462
rect 57260 34244 57316 39564
rect 57372 39554 57428 39564
rect 57596 38724 57652 38734
rect 57596 38630 57652 38668
rect 57708 38500 57764 40124
rect 57820 39620 57876 39630
rect 57820 39526 57876 39564
rect 58268 39620 58324 40236
rect 58268 39554 58324 39564
rect 57596 38444 57764 38500
rect 57932 38836 57988 38846
rect 57484 37492 57540 37502
rect 57596 37492 57652 38444
rect 57820 38162 57876 38174
rect 57820 38110 57822 38162
rect 57874 38110 57876 38162
rect 57484 37490 57652 37492
rect 57484 37438 57486 37490
rect 57538 37438 57652 37490
rect 57484 37436 57652 37438
rect 57708 38050 57764 38062
rect 57708 37998 57710 38050
rect 57762 37998 57764 38050
rect 57484 37426 57540 37436
rect 57708 37378 57764 37998
rect 57708 37326 57710 37378
rect 57762 37326 57764 37378
rect 57372 36764 57652 36820
rect 57372 36482 57428 36764
rect 57372 36430 57374 36482
rect 57426 36430 57428 36482
rect 57372 36418 57428 36430
rect 57484 36594 57540 36606
rect 57484 36542 57486 36594
rect 57538 36542 57540 36594
rect 57484 35810 57540 36542
rect 57484 35758 57486 35810
rect 57538 35758 57540 35810
rect 57372 35028 57428 35038
rect 57484 35028 57540 35758
rect 57372 35026 57540 35028
rect 57372 34974 57374 35026
rect 57426 34974 57540 35026
rect 57372 34972 57540 34974
rect 57596 35700 57652 36764
rect 57708 36148 57764 37326
rect 57820 37378 57876 38110
rect 57820 37326 57822 37378
rect 57874 37326 57876 37378
rect 57820 36594 57876 37326
rect 57820 36542 57822 36594
rect 57874 36542 57876 36594
rect 57820 36530 57876 36542
rect 57932 36372 57988 38780
rect 58380 38050 58436 43372
rect 58492 38946 58548 43652
rect 58492 38894 58494 38946
rect 58546 38894 58548 38946
rect 58492 38882 58548 38894
rect 58380 37998 58382 38050
rect 58434 37998 58436 38050
rect 58380 37986 58436 37998
rect 57708 36082 57764 36092
rect 57820 36316 57988 36372
rect 57708 35924 57764 35934
rect 57820 35924 57876 36316
rect 57708 35922 57876 35924
rect 57708 35870 57710 35922
rect 57762 35870 57876 35922
rect 57708 35868 57876 35870
rect 58044 36036 58100 36046
rect 57708 35858 57764 35868
rect 57708 35700 57764 35710
rect 57596 35698 57764 35700
rect 57596 35646 57710 35698
rect 57762 35646 57764 35698
rect 57596 35644 57764 35646
rect 57372 34962 57428 34972
rect 57484 34244 57540 34254
rect 57260 34242 57540 34244
rect 57260 34190 57486 34242
rect 57538 34190 57540 34242
rect 57260 34188 57540 34190
rect 57484 34178 57540 34188
rect 57596 34020 57652 35644
rect 57708 35634 57764 35644
rect 57932 35700 57988 35710
rect 57932 35606 57988 35644
rect 57372 33964 57652 34020
rect 57708 34188 57988 34244
rect 57372 32004 57428 33964
rect 57484 33346 57540 33358
rect 57484 33294 57486 33346
rect 57538 33294 57540 33346
rect 57484 32786 57540 33294
rect 57708 33124 57764 34188
rect 57932 34130 57988 34188
rect 57932 34078 57934 34130
rect 57986 34078 57988 34130
rect 57932 34066 57988 34078
rect 58044 33908 58100 35980
rect 58268 34020 58324 34030
rect 57932 33852 58100 33908
rect 58156 34018 58324 34020
rect 58156 33966 58270 34018
rect 58322 33966 58324 34018
rect 58156 33964 58324 33966
rect 57932 33458 57988 33852
rect 57932 33406 57934 33458
rect 57986 33406 57988 33458
rect 57932 33394 57988 33406
rect 58044 33348 58100 33358
rect 58156 33348 58212 33964
rect 58268 33954 58324 33964
rect 58044 33346 58212 33348
rect 58044 33294 58046 33346
rect 58098 33294 58212 33346
rect 58044 33292 58212 33294
rect 58044 33282 58100 33292
rect 57820 33124 57876 33134
rect 57708 33122 57876 33124
rect 57708 33070 57822 33122
rect 57874 33070 57876 33122
rect 57708 33068 57876 33070
rect 57484 32734 57486 32786
rect 57538 32734 57540 32786
rect 57484 32722 57540 32734
rect 57820 32788 57876 33068
rect 57820 32732 57988 32788
rect 57708 32676 57764 32686
rect 57372 31938 57428 31948
rect 57596 32674 57764 32676
rect 57596 32622 57710 32674
rect 57762 32622 57764 32674
rect 57596 32620 57764 32622
rect 57596 31778 57652 32620
rect 57708 32610 57764 32620
rect 57820 32564 57876 32574
rect 57820 32452 57876 32508
rect 57708 32396 57876 32452
rect 57708 31890 57764 32396
rect 57932 31948 57988 32732
rect 57708 31838 57710 31890
rect 57762 31838 57764 31890
rect 57708 31826 57764 31838
rect 57820 31892 57988 31948
rect 58156 32002 58212 33292
rect 58156 31950 58158 32002
rect 58210 31950 58212 32002
rect 58156 31938 58212 31950
rect 57596 31726 57598 31778
rect 57650 31726 57652 31778
rect 57484 30882 57540 30894
rect 57484 30830 57486 30882
rect 57538 30830 57540 30882
rect 57372 30772 57428 30782
rect 57372 30322 57428 30716
rect 57372 30270 57374 30322
rect 57426 30270 57428 30322
rect 57372 30258 57428 30270
rect 57260 30210 57316 30222
rect 57260 30158 57262 30210
rect 57314 30158 57316 30210
rect 57260 30100 57316 30158
rect 57484 30100 57540 30830
rect 57260 30044 57540 30100
rect 57260 28980 57316 30044
rect 57484 29540 57540 29550
rect 57484 29446 57540 29484
rect 57260 28914 57316 28924
rect 57596 28756 57652 31726
rect 57708 30772 57764 30782
rect 57708 30678 57764 30716
rect 57820 29650 57876 31892
rect 58044 30772 58100 30782
rect 58044 30770 58324 30772
rect 58044 30718 58046 30770
rect 58098 30718 58324 30770
rect 58044 30716 58324 30718
rect 58044 30706 58100 30716
rect 57820 29598 57822 29650
rect 57874 29598 57876 29650
rect 57820 29586 57876 29598
rect 58156 30098 58212 30110
rect 58156 30046 58158 30098
rect 58210 30046 58212 30098
rect 57708 29426 57764 29438
rect 57708 29374 57710 29426
rect 57762 29374 57764 29426
rect 57708 28980 57764 29374
rect 58044 29426 58100 29438
rect 58044 29374 58046 29426
rect 58098 29374 58100 29426
rect 58044 29204 58100 29374
rect 58044 29138 58100 29148
rect 57708 28914 57764 28924
rect 57820 28756 57876 28766
rect 57596 28754 57876 28756
rect 57596 28702 57822 28754
rect 57874 28702 57876 28754
rect 57596 28700 57876 28702
rect 57820 28690 57876 28700
rect 57932 28644 57988 28654
rect 58156 28644 58212 30046
rect 57932 28642 58212 28644
rect 57932 28590 57934 28642
rect 57986 28590 58212 28642
rect 57932 28588 58212 28590
rect 58268 28642 58324 30716
rect 58268 28590 58270 28642
rect 58322 28590 58324 28642
rect 57932 28578 57988 28588
rect 57148 28532 57204 28542
rect 57708 28532 57764 28542
rect 57148 28530 57764 28532
rect 57148 28478 57150 28530
rect 57202 28478 57710 28530
rect 57762 28478 57764 28530
rect 57148 28476 57764 28478
rect 57148 28466 57204 28476
rect 57372 27186 57428 28476
rect 57708 28466 57764 28476
rect 57372 27134 57374 27186
rect 57426 27134 57428 27186
rect 57372 27122 57428 27134
rect 58044 27074 58100 28588
rect 58268 28578 58324 28590
rect 58044 27022 58046 27074
rect 58098 27022 58100 27074
rect 58044 27010 58100 27022
rect 56252 24882 56308 24892
rect 56924 25116 57092 25172
rect 57148 26962 57204 26974
rect 57148 26910 57150 26962
rect 57202 26910 57204 26962
rect 57148 25618 57204 26910
rect 57932 26852 57988 26862
rect 57596 26292 57652 26302
rect 57596 26198 57652 26236
rect 57932 26290 57988 26796
rect 57932 26238 57934 26290
rect 57986 26238 57988 26290
rect 57932 26226 57988 26238
rect 57148 25566 57150 25618
rect 57202 25566 57204 25618
rect 56140 23774 56142 23826
rect 56194 23774 56196 23826
rect 55692 23380 55748 23390
rect 56140 23380 56196 23774
rect 55692 23378 56196 23380
rect 55692 23326 55694 23378
rect 55746 23326 56142 23378
rect 56194 23326 56196 23378
rect 55692 23324 56196 23326
rect 55692 23314 55748 23324
rect 54684 22878 54686 22930
rect 54738 22878 54740 22930
rect 54460 22372 54516 22382
rect 54684 22372 54740 22878
rect 54460 22370 54740 22372
rect 54460 22318 54462 22370
rect 54514 22318 54740 22370
rect 54460 22316 54740 22318
rect 54460 22306 54516 22316
rect 55132 22260 55188 22270
rect 55132 22258 55412 22260
rect 55132 22206 55134 22258
rect 55186 22206 55412 22258
rect 55132 22204 55412 22206
rect 55132 22194 55188 22204
rect 54124 21758 54126 21810
rect 54178 21758 54180 21810
rect 54124 21746 54180 21758
rect 53788 21534 53790 21586
rect 53842 21534 53844 21586
rect 53788 21522 53844 21534
rect 55356 21586 55412 22204
rect 56028 22258 56084 23324
rect 56140 23314 56196 23324
rect 56364 23938 56420 23950
rect 56364 23886 56366 23938
rect 56418 23886 56420 23938
rect 56364 23828 56420 23886
rect 56364 22482 56420 23772
rect 56364 22430 56366 22482
rect 56418 22430 56420 22482
rect 56364 22418 56420 22430
rect 56028 22206 56030 22258
rect 56082 22206 56084 22258
rect 56028 22194 56084 22206
rect 55356 21534 55358 21586
rect 55410 21534 55412 21586
rect 54348 21364 54404 21374
rect 54348 20802 54404 21308
rect 54348 20750 54350 20802
rect 54402 20750 54404 20802
rect 54348 20738 54404 20750
rect 54796 21364 54852 21374
rect 54684 20692 54740 20702
rect 54684 20598 54740 20636
rect 53788 20578 53844 20590
rect 53788 20526 53790 20578
rect 53842 20526 53844 20578
rect 53676 20468 53732 20478
rect 53452 20130 53508 20142
rect 53452 20078 53454 20130
rect 53506 20078 53508 20130
rect 53452 19124 53508 20078
rect 53676 19234 53732 20412
rect 53788 20132 53844 20526
rect 53788 19796 53844 20076
rect 54460 20578 54516 20590
rect 54460 20526 54462 20578
rect 54514 20526 54516 20578
rect 54460 19908 54516 20526
rect 54460 19842 54516 19852
rect 54796 20130 54852 21308
rect 55020 21362 55076 21374
rect 55020 21310 55022 21362
rect 55074 21310 55076 21362
rect 55020 20468 55076 21310
rect 55356 21364 55412 21534
rect 56364 22148 56420 22158
rect 55356 21298 55412 21308
rect 55580 21474 55636 21486
rect 55580 21422 55582 21474
rect 55634 21422 55636 21474
rect 55020 20402 55076 20412
rect 55580 20188 55636 21422
rect 56140 21362 56196 21374
rect 56140 21310 56142 21362
rect 56194 21310 56196 21362
rect 56028 20692 56084 20702
rect 56028 20598 56084 20636
rect 55580 20132 55748 20188
rect 54796 20078 54798 20130
rect 54850 20078 54852 20130
rect 53788 19730 53844 19740
rect 54012 19796 54068 19806
rect 53676 19182 53678 19234
rect 53730 19182 53732 19234
rect 53676 19170 53732 19182
rect 53788 19236 53844 19246
rect 53452 19058 53508 19068
rect 53564 18676 53620 18686
rect 53452 18564 53508 18574
rect 53452 18338 53508 18508
rect 53452 18286 53454 18338
rect 53506 18286 53508 18338
rect 53452 18274 53508 18286
rect 53452 17780 53508 17790
rect 53564 17780 53620 18620
rect 53452 17778 53620 17780
rect 53452 17726 53454 17778
rect 53506 17726 53620 17778
rect 53452 17724 53620 17726
rect 53788 17778 53844 19180
rect 53900 19124 53956 19134
rect 53900 19030 53956 19068
rect 54012 18676 54068 19740
rect 54348 19236 54404 19246
rect 54348 19142 54404 19180
rect 54012 18562 54068 18620
rect 54012 18510 54014 18562
rect 54066 18510 54068 18562
rect 54012 18498 54068 18510
rect 54124 19010 54180 19022
rect 54124 18958 54126 19010
rect 54178 18958 54180 19010
rect 54124 18452 54180 18958
rect 54796 18452 54852 20078
rect 55692 20020 55748 20132
rect 55692 19954 55748 19964
rect 56028 20018 56084 20030
rect 56028 19966 56030 20018
rect 56082 19966 56084 20018
rect 55020 19908 55076 19918
rect 55020 19814 55076 19852
rect 55468 19908 55524 19918
rect 56028 19908 56084 19966
rect 55468 19906 55636 19908
rect 55468 19854 55470 19906
rect 55522 19854 55636 19906
rect 55468 19852 55636 19854
rect 55468 19842 55524 19852
rect 55468 19236 55524 19246
rect 55468 19142 55524 19180
rect 55356 19124 55412 19134
rect 55356 19030 55412 19068
rect 55580 19124 55636 19852
rect 56028 19842 56084 19852
rect 56140 19236 56196 21310
rect 56364 20802 56420 22092
rect 56588 21476 56644 21486
rect 56476 21364 56532 21374
rect 56476 21270 56532 21308
rect 56364 20750 56366 20802
rect 56418 20750 56420 20802
rect 56140 19170 56196 19180
rect 56252 20018 56308 20030
rect 56252 19966 56254 20018
rect 56306 19966 56308 20018
rect 55580 19058 55636 19068
rect 56028 19010 56084 19022
rect 56028 18958 56030 19010
rect 56082 18958 56084 19010
rect 56028 18564 56084 18958
rect 56084 18508 56196 18564
rect 56028 18498 56084 18508
rect 54908 18452 54964 18462
rect 54796 18450 54964 18452
rect 54796 18398 54910 18450
rect 54962 18398 54964 18450
rect 54796 18396 54964 18398
rect 54124 18386 54180 18396
rect 54908 18386 54964 18396
rect 55916 18452 55972 18462
rect 53788 17726 53790 17778
rect 53842 17726 53844 17778
rect 53452 17714 53508 17724
rect 53788 17332 53844 17726
rect 53228 17052 53620 17108
rect 53340 16884 53396 16894
rect 52332 16830 52334 16882
rect 52386 16830 52388 16882
rect 52332 16818 52388 16830
rect 53004 16882 53396 16884
rect 53004 16830 53342 16882
rect 53394 16830 53396 16882
rect 53004 16828 53396 16830
rect 50316 16718 50318 16770
rect 50370 16718 50372 16770
rect 50316 16706 50372 16718
rect 50764 16772 50820 16782
rect 52892 16772 52948 16782
rect 50764 16770 50932 16772
rect 50764 16718 50766 16770
rect 50818 16718 50932 16770
rect 50764 16716 50932 16718
rect 50764 16706 50820 16716
rect 49196 15874 49364 15876
rect 49196 15822 49198 15874
rect 49250 15822 49364 15874
rect 49196 15820 49364 15822
rect 49756 15876 49812 15886
rect 49196 15428 49252 15820
rect 49756 15538 49812 15820
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 49756 15486 49758 15538
rect 49810 15486 49812 15538
rect 49756 15474 49812 15486
rect 48412 15204 48468 15242
rect 48412 15138 48468 15148
rect 46956 14578 47012 14588
rect 47292 14588 47460 14644
rect 46844 14478 46846 14530
rect 46898 14478 46900 14530
rect 46844 14466 46900 14478
rect 46060 14084 46116 14094
rect 46060 13970 46116 14028
rect 46060 13918 46062 13970
rect 46114 13918 46116 13970
rect 46060 13906 46116 13918
rect 46620 14084 46676 14094
rect 46620 13858 46676 14028
rect 46620 13806 46622 13858
rect 46674 13806 46676 13858
rect 45948 13636 46004 13646
rect 45948 12402 46004 13580
rect 46396 13636 46452 13646
rect 45948 12350 45950 12402
rect 46002 12350 46004 12402
rect 45948 12338 46004 12350
rect 46060 13076 46116 13086
rect 46060 11396 46116 13020
rect 46396 12962 46452 13580
rect 46620 13074 46676 13806
rect 46844 13858 46900 13870
rect 46844 13806 46846 13858
rect 46898 13806 46900 13858
rect 46844 13636 46900 13806
rect 46844 13570 46900 13580
rect 46620 13022 46622 13074
rect 46674 13022 46676 13074
rect 46620 13010 46676 13022
rect 46956 13522 47012 13534
rect 46956 13470 46958 13522
rect 47010 13470 47012 13522
rect 46396 12910 46398 12962
rect 46450 12910 46452 12962
rect 46396 12898 46452 12910
rect 46956 12292 47012 13470
rect 47292 13076 47348 14588
rect 47404 14420 47460 14430
rect 48636 14420 48692 15260
rect 49196 15204 49252 15372
rect 49980 15428 50036 15438
rect 48860 15148 49252 15204
rect 49532 15314 49588 15326
rect 49532 15262 49534 15314
rect 49586 15262 49588 15314
rect 49532 15204 49588 15262
rect 49644 15316 49700 15326
rect 49644 15222 49700 15260
rect 48748 15090 48804 15102
rect 48748 15038 48750 15090
rect 48802 15038 48804 15090
rect 48748 14644 48804 15038
rect 48748 14578 48804 14588
rect 48860 14642 48916 15148
rect 49532 15138 49588 15148
rect 48860 14590 48862 14642
rect 48914 14590 48916 14642
rect 48860 14578 48916 14590
rect 49644 14644 49700 14654
rect 49644 14550 49700 14588
rect 49980 14530 50036 15372
rect 50876 14756 50932 16716
rect 52668 16770 52948 16772
rect 52668 16718 52894 16770
rect 52946 16718 52948 16770
rect 52668 16716 52948 16718
rect 52444 15988 52500 15998
rect 52444 15894 52500 15932
rect 52668 15988 52724 16716
rect 52892 16706 52948 16716
rect 53004 16436 53060 16828
rect 53340 16818 53396 16828
rect 52780 16380 53060 16436
rect 52780 16098 52836 16380
rect 52780 16046 52782 16098
rect 52834 16046 52836 16098
rect 52780 16034 52836 16046
rect 52668 15922 52724 15932
rect 53452 15988 53508 15998
rect 53452 15894 53508 15932
rect 52556 15876 52612 15886
rect 52556 15426 52612 15820
rect 52556 15374 52558 15426
rect 52610 15374 52612 15426
rect 52556 15362 52612 15374
rect 52444 15316 52500 15326
rect 52220 15314 52500 15316
rect 52220 15262 52446 15314
rect 52498 15262 52500 15314
rect 52220 15260 52500 15262
rect 50876 14690 50932 14700
rect 51884 14756 51940 14766
rect 51884 14662 51940 14700
rect 52220 14754 52276 15260
rect 52444 15250 52500 15260
rect 52668 15316 52724 15326
rect 53340 15316 53396 15326
rect 52220 14702 52222 14754
rect 52274 14702 52276 14754
rect 52220 14690 52276 14702
rect 52332 14756 52388 14766
rect 49980 14478 49982 14530
rect 50034 14478 50036 14530
rect 49980 14466 50036 14478
rect 50316 14642 50372 14654
rect 50316 14590 50318 14642
rect 50370 14590 50372 14642
rect 47404 14418 47572 14420
rect 47404 14366 47406 14418
rect 47458 14366 47572 14418
rect 47404 14364 47572 14366
rect 48636 14364 48804 14420
rect 47404 14354 47460 14364
rect 47292 13010 47348 13020
rect 47404 13746 47460 13758
rect 47404 13694 47406 13746
rect 47458 13694 47460 13746
rect 47180 12292 47236 12302
rect 46956 12290 47236 12292
rect 46956 12238 47182 12290
rect 47234 12238 47236 12290
rect 46956 12236 47236 12238
rect 47180 12226 47236 12236
rect 47404 12290 47460 13694
rect 47516 12964 47572 14364
rect 47852 14308 47908 14318
rect 47628 14306 47908 14308
rect 47628 14254 47854 14306
rect 47906 14254 47908 14306
rect 47628 14252 47908 14254
rect 47628 13858 47684 14252
rect 47852 14242 47908 14252
rect 47628 13806 47630 13858
rect 47682 13806 47684 13858
rect 47628 13636 47684 13806
rect 47740 14084 47796 14094
rect 47740 13858 47796 14028
rect 48188 14084 48244 14094
rect 48188 13970 48244 14028
rect 48188 13918 48190 13970
rect 48242 13918 48244 13970
rect 48188 13906 48244 13918
rect 47740 13806 47742 13858
rect 47794 13806 47796 13858
rect 47740 13794 47796 13806
rect 47628 13570 47684 13580
rect 47740 12964 47796 12974
rect 47516 12962 47796 12964
rect 47516 12910 47742 12962
rect 47794 12910 47796 12962
rect 47516 12908 47796 12910
rect 47628 12404 47684 12414
rect 47628 12310 47684 12348
rect 47404 12238 47406 12290
rect 47458 12238 47460 12290
rect 47404 12226 47460 12238
rect 47740 12290 47796 12908
rect 47740 12238 47742 12290
rect 47794 12238 47796 12290
rect 47740 12226 47796 12238
rect 48524 12850 48580 12862
rect 48524 12798 48526 12850
rect 48578 12798 48580 12850
rect 44716 11282 45108 11284
rect 44716 11230 44718 11282
rect 44770 11230 45108 11282
rect 44716 11228 45108 11230
rect 44716 11218 44772 11228
rect 44156 10834 44660 10836
rect 44156 10782 44158 10834
rect 44210 10782 44660 10834
rect 44156 10780 44660 10782
rect 44156 10770 44212 10780
rect 44268 10612 44324 10622
rect 44716 10612 44772 10622
rect 44156 10610 44772 10612
rect 44156 10558 44270 10610
rect 44322 10558 44718 10610
rect 44770 10558 44772 10610
rect 44156 10556 44772 10558
rect 44156 9604 44212 10556
rect 44268 10546 44324 10556
rect 44716 10546 44772 10556
rect 44268 10052 44324 10062
rect 44268 9716 44324 9996
rect 44604 9828 44660 9838
rect 44604 9734 44660 9772
rect 44268 9650 44324 9660
rect 44156 9538 44212 9548
rect 44380 9602 44436 9614
rect 44380 9550 44382 9602
rect 44434 9550 44436 9602
rect 43932 8818 44100 8820
rect 43932 8766 43934 8818
rect 43986 8766 44100 8818
rect 43932 8764 44100 8766
rect 44156 9156 44212 9166
rect 44380 9156 44436 9550
rect 44492 9156 44548 9166
rect 44380 9154 44548 9156
rect 44380 9102 44494 9154
rect 44546 9102 44548 9154
rect 44380 9100 44548 9102
rect 43932 8372 43988 8764
rect 43932 7700 43988 8316
rect 44156 8258 44212 9100
rect 44492 9090 44548 9100
rect 44716 9156 44772 9166
rect 44716 9062 44772 9100
rect 44940 9156 44996 9166
rect 44940 9062 44996 9100
rect 45052 9154 45108 11228
rect 45836 11218 45892 11228
rect 45948 11340 46116 11396
rect 45164 10498 45220 10510
rect 45164 10446 45166 10498
rect 45218 10446 45220 10498
rect 45164 9828 45220 10446
rect 45612 10498 45668 10510
rect 45612 10446 45614 10498
rect 45666 10446 45668 10498
rect 45612 10052 45668 10446
rect 45612 9986 45668 9996
rect 45164 9762 45220 9772
rect 45388 9604 45444 9614
rect 45388 9268 45444 9548
rect 45500 9268 45556 9278
rect 45388 9266 45556 9268
rect 45388 9214 45502 9266
rect 45554 9214 45556 9266
rect 45388 9212 45556 9214
rect 45500 9202 45556 9212
rect 45052 9102 45054 9154
rect 45106 9102 45108 9154
rect 45052 8428 45108 9102
rect 44156 8206 44158 8258
rect 44210 8206 44212 8258
rect 44156 8194 44212 8206
rect 44604 8372 45108 8428
rect 45948 9156 46004 11340
rect 47068 11284 47124 11294
rect 46060 11172 46116 11182
rect 46620 11172 46676 11182
rect 46060 11170 46676 11172
rect 46060 11118 46062 11170
rect 46114 11118 46622 11170
rect 46674 11118 46676 11170
rect 46060 11116 46676 11118
rect 46060 11106 46116 11116
rect 46284 10050 46340 11116
rect 46620 11106 46676 11116
rect 46732 11172 46788 11182
rect 46732 11078 46788 11116
rect 46844 11170 46900 11182
rect 46844 11118 46846 11170
rect 46898 11118 46900 11170
rect 46844 11060 46900 11118
rect 46284 9998 46286 10050
rect 46338 9998 46340 10050
rect 46284 9986 46340 9998
rect 46620 10610 46676 10622
rect 46620 10558 46622 10610
rect 46674 10558 46676 10610
rect 46620 10050 46676 10558
rect 46620 9998 46622 10050
rect 46674 9998 46676 10050
rect 46620 9986 46676 9998
rect 46620 9828 46676 9838
rect 46844 9828 46900 11004
rect 47068 10498 47124 11228
rect 47068 10446 47070 10498
rect 47122 10446 47124 10498
rect 47068 10434 47124 10446
rect 47404 10610 47460 10622
rect 47404 10558 47406 10610
rect 47458 10558 47460 10610
rect 46620 9826 46900 9828
rect 46620 9774 46622 9826
rect 46674 9774 46900 9826
rect 46620 9772 46900 9774
rect 47068 9828 47124 9838
rect 46620 9762 46676 9772
rect 47068 9734 47124 9772
rect 46284 9156 46340 9166
rect 45948 9154 46340 9156
rect 45948 9102 46286 9154
rect 46338 9102 46340 9154
rect 45948 9100 46340 9102
rect 44604 8258 44660 8372
rect 44604 8206 44606 8258
rect 44658 8206 44660 8258
rect 44604 8194 44660 8206
rect 44716 8146 44772 8158
rect 44716 8094 44718 8146
rect 44770 8094 44772 8146
rect 43932 7634 43988 7644
rect 44492 7700 44548 7710
rect 44492 7606 44548 7644
rect 42924 7310 42926 7362
rect 42978 7310 42980 7362
rect 42924 7298 42980 7310
rect 43820 7364 43876 7420
rect 43932 7364 43988 7374
rect 43820 7362 43988 7364
rect 43820 7310 43934 7362
rect 43986 7310 43988 7362
rect 43820 7308 43988 7310
rect 43820 6802 43876 7308
rect 43932 7298 43988 7308
rect 43820 6750 43822 6802
rect 43874 6750 43876 6802
rect 43820 6738 43876 6750
rect 42588 6524 43204 6580
rect 42476 5954 42532 5964
rect 42140 5684 42196 5694
rect 42140 5682 43092 5684
rect 42140 5630 42142 5682
rect 42194 5630 43092 5682
rect 42140 5628 43092 5630
rect 42140 5618 42196 5628
rect 42924 5236 42980 5246
rect 41916 5180 42084 5236
rect 41020 5070 41022 5122
rect 41074 5070 41076 5122
rect 41020 5058 41076 5070
rect 41132 5122 41636 5124
rect 41132 5070 41358 5122
rect 41410 5070 41636 5122
rect 41132 5068 41636 5070
rect 41692 5122 41748 5134
rect 41692 5070 41694 5122
rect 41746 5070 41748 5122
rect 40124 4498 40180 4508
rect 40572 4900 40628 4910
rect 40572 4450 40628 4844
rect 41132 4788 41188 5068
rect 41356 5058 41412 5068
rect 41692 4900 41748 5070
rect 41804 5124 41860 5134
rect 41804 5030 41860 5068
rect 41916 5012 41972 5022
rect 41916 4918 41972 4956
rect 41692 4834 41748 4844
rect 40908 4732 41188 4788
rect 40684 4564 40740 4574
rect 40684 4470 40740 4508
rect 40908 4562 40964 4732
rect 40908 4510 40910 4562
rect 40962 4510 40964 4562
rect 40908 4498 40964 4510
rect 42028 4564 42084 5180
rect 42924 5142 42980 5180
rect 43036 5122 43092 5628
rect 43036 5070 43038 5122
rect 43090 5070 43092 5122
rect 43036 5058 43092 5070
rect 42476 5012 42532 5022
rect 42532 4956 42644 5012
rect 42476 4918 42532 4956
rect 40572 4398 40574 4450
rect 40626 4398 40628 4450
rect 40572 4386 40628 4398
rect 37436 4338 37604 4340
rect 37436 4286 37438 4338
rect 37490 4286 37604 4338
rect 37436 4284 37604 4286
rect 37436 4274 37492 4284
rect 37100 3554 37268 3556
rect 37100 3502 37102 3554
rect 37154 3502 37268 3554
rect 37100 3500 37268 3502
rect 37324 4228 37380 4238
rect 37324 3554 37380 4172
rect 37324 3502 37326 3554
rect 37378 3502 37380 3554
rect 37100 3490 37156 3500
rect 37324 3490 37380 3502
rect 37436 3892 37492 3902
rect 34972 3444 35028 3482
rect 34972 3378 35028 3388
rect 33628 3266 33684 3276
rect 37212 3332 37268 3342
rect 37436 3332 37492 3836
rect 37548 3442 37604 4284
rect 42028 4338 42084 4508
rect 42028 4286 42030 4338
rect 42082 4286 42084 4338
rect 38780 4226 38836 4238
rect 38780 4174 38782 4226
rect 38834 4174 38836 4226
rect 37884 4116 37940 4126
rect 37884 4022 37940 4060
rect 38780 3892 38836 4174
rect 41916 4226 41972 4238
rect 41916 4174 41918 4226
rect 41970 4174 41972 4226
rect 39004 4116 39060 4126
rect 39004 4022 39060 4060
rect 39340 4116 39396 4126
rect 39340 4022 39396 4060
rect 41020 4116 41076 4126
rect 38780 3826 38836 3836
rect 39452 3668 39508 3678
rect 39452 3574 39508 3612
rect 41020 3554 41076 4060
rect 41916 4116 41972 4174
rect 41916 4050 41972 4060
rect 41020 3502 41022 3554
rect 41074 3502 41076 3554
rect 41020 3490 41076 3502
rect 41916 3892 41972 3902
rect 37548 3390 37550 3442
rect 37602 3390 37604 3442
rect 37548 3378 37604 3390
rect 38556 3444 38612 3454
rect 40348 3444 40404 3454
rect 38556 3442 38836 3444
rect 38556 3390 38558 3442
rect 38610 3390 38836 3442
rect 38556 3388 38836 3390
rect 38556 3378 38612 3388
rect 37212 3330 37492 3332
rect 37212 3278 37214 3330
rect 37266 3278 37492 3330
rect 37212 3276 37492 3278
rect 38780 3332 38836 3388
rect 40348 3350 40404 3388
rect 41132 3444 41188 3454
rect 41132 3350 41188 3388
rect 41356 3444 41412 3454
rect 41804 3444 41860 3454
rect 41356 3442 41860 3444
rect 41356 3390 41358 3442
rect 41410 3390 41806 3442
rect 41858 3390 41860 3442
rect 41356 3388 41860 3390
rect 41356 3378 41412 3388
rect 41804 3378 41860 3388
rect 41916 3442 41972 3836
rect 41916 3390 41918 3442
rect 41970 3390 41972 3442
rect 41916 3378 41972 3390
rect 42028 3444 42084 4286
rect 42140 4788 42196 4798
rect 42140 3554 42196 4732
rect 42588 4226 42644 4956
rect 42700 5010 42756 5022
rect 42700 4958 42702 5010
rect 42754 4958 42756 5010
rect 42700 4900 42756 4958
rect 43148 5012 43204 6524
rect 44492 6244 44548 6254
rect 44044 6132 44100 6142
rect 43820 5906 43876 5918
rect 43820 5854 43822 5906
rect 43874 5854 43876 5906
rect 43260 5796 43316 5806
rect 43260 5702 43316 5740
rect 43820 5236 43876 5854
rect 43820 5170 43876 5180
rect 43932 5908 43988 5918
rect 43148 4946 43204 4956
rect 42700 4834 42756 4844
rect 43148 4564 43204 4574
rect 43148 4470 43204 4508
rect 43932 4452 43988 5852
rect 44044 5796 44100 6076
rect 44492 6130 44548 6188
rect 44492 6078 44494 6130
rect 44546 6078 44548 6130
rect 44492 6066 44548 6078
rect 44044 5122 44100 5740
rect 44380 5906 44436 5918
rect 44380 5854 44382 5906
rect 44434 5854 44436 5906
rect 44044 5070 44046 5122
rect 44098 5070 44100 5122
rect 44044 5058 44100 5070
rect 44156 5682 44212 5694
rect 44156 5630 44158 5682
rect 44210 5630 44212 5682
rect 44156 5124 44212 5630
rect 44156 5058 44212 5068
rect 44380 4788 44436 5854
rect 44604 5908 44660 5918
rect 44604 5814 44660 5852
rect 44716 5684 44772 8094
rect 45948 8036 46004 9100
rect 46284 9090 46340 9100
rect 46508 9156 46564 9166
rect 45948 8034 46116 8036
rect 45948 7982 45950 8034
rect 46002 7982 46116 8034
rect 45948 7980 46116 7982
rect 45948 7970 46004 7980
rect 45388 7588 45444 7598
rect 46060 7588 46116 7980
rect 45388 7586 46116 7588
rect 45388 7534 45390 7586
rect 45442 7534 46116 7586
rect 45388 7532 46116 7534
rect 45388 7522 45444 7532
rect 46060 7474 46116 7532
rect 46060 7422 46062 7474
rect 46114 7422 46116 7474
rect 46060 7410 46116 7422
rect 46508 7474 46564 9100
rect 46956 9156 47012 9166
rect 46620 9044 46676 9054
rect 46620 8930 46676 8988
rect 46620 8878 46622 8930
rect 46674 8878 46676 8930
rect 46620 8866 46676 8878
rect 46956 8258 47012 9100
rect 47404 9156 47460 10558
rect 48524 10164 48580 12798
rect 48748 10836 48804 14364
rect 49308 13076 49364 13086
rect 49308 12292 49364 13020
rect 49756 12962 49812 12974
rect 49756 12910 49758 12962
rect 49810 12910 49812 12962
rect 49644 12852 49700 12862
rect 49644 12402 49700 12796
rect 49644 12350 49646 12402
rect 49698 12350 49700 12402
rect 49644 12338 49700 12350
rect 49756 12404 49812 12910
rect 50316 12964 50372 14590
rect 51660 14530 51716 14542
rect 51660 14478 51662 14530
rect 51714 14478 51716 14530
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 51660 13636 51716 14478
rect 52332 13860 52388 14700
rect 51996 13636 52052 13646
rect 51660 13634 52164 13636
rect 51660 13582 51998 13634
rect 52050 13582 52164 13634
rect 51660 13580 52164 13582
rect 51996 13570 52052 13580
rect 51212 13076 51268 13086
rect 51212 12982 51268 13020
rect 52108 13076 52164 13580
rect 52332 13186 52388 13804
rect 52668 13858 52724 15260
rect 52668 13806 52670 13858
rect 52722 13806 52724 13858
rect 52668 13794 52724 13806
rect 52780 15314 53396 15316
rect 52780 15262 53342 15314
rect 53394 15262 53396 15314
rect 52780 15260 53396 15262
rect 52332 13134 52334 13186
rect 52386 13134 52388 13186
rect 52332 13122 52388 13134
rect 52668 13188 52724 13198
rect 52780 13188 52836 15260
rect 53340 15250 53396 15260
rect 53564 14868 53620 17052
rect 53788 17106 53844 17276
rect 53788 17054 53790 17106
rect 53842 17054 53844 17106
rect 53788 17042 53844 17054
rect 55468 17666 55524 17678
rect 55468 17614 55470 17666
rect 55522 17614 55524 17666
rect 53900 16996 53956 17006
rect 53900 16902 53956 16940
rect 53676 16884 53732 16894
rect 53676 16210 53732 16828
rect 54012 16884 54068 16894
rect 54012 16790 54068 16828
rect 55020 16884 55076 16894
rect 53676 16158 53678 16210
rect 53730 16158 53732 16210
rect 53676 16146 53732 16158
rect 55020 16098 55076 16828
rect 55020 16046 55022 16098
rect 55074 16046 55076 16098
rect 55020 16034 55076 16046
rect 55244 16882 55300 16894
rect 55244 16830 55246 16882
rect 55298 16830 55300 16882
rect 54460 15988 54516 15998
rect 53676 15876 53732 15886
rect 53676 15782 53732 15820
rect 54236 15876 54292 15886
rect 53564 14802 53620 14812
rect 54236 15314 54292 15820
rect 54236 15262 54238 15314
rect 54290 15262 54292 15314
rect 54236 14530 54292 15262
rect 54236 14478 54238 14530
rect 54290 14478 54292 14530
rect 54236 14466 54292 14478
rect 54460 15090 54516 15932
rect 55244 15988 55300 16830
rect 55244 15894 55300 15932
rect 54796 15316 54852 15326
rect 54796 15222 54852 15260
rect 54460 15038 54462 15090
rect 54514 15038 54516 15090
rect 54460 14530 54516 15038
rect 54684 14644 54740 14654
rect 55468 14644 55524 17614
rect 55692 17554 55748 17566
rect 55692 17502 55694 17554
rect 55746 17502 55748 17554
rect 55580 16884 55636 16894
rect 55580 16790 55636 16828
rect 55692 16212 55748 17502
rect 55916 16770 55972 18396
rect 56028 18338 56084 18350
rect 56028 18286 56030 18338
rect 56082 18286 56084 18338
rect 56028 16884 56084 18286
rect 56028 16818 56084 16828
rect 55916 16718 55918 16770
rect 55970 16718 55972 16770
rect 55916 16706 55972 16718
rect 55916 16212 55972 16222
rect 55692 16210 55972 16212
rect 55692 16158 55918 16210
rect 55970 16158 55972 16210
rect 55692 16156 55972 16158
rect 55916 16146 55972 16156
rect 56140 16098 56196 18508
rect 56252 18452 56308 19966
rect 56252 18386 56308 18396
rect 56364 18004 56420 20750
rect 56476 20244 56532 20282
rect 56476 20178 56532 20188
rect 56588 20130 56644 21420
rect 56700 21476 56756 21486
rect 56700 21474 56868 21476
rect 56700 21422 56702 21474
rect 56754 21422 56868 21474
rect 56700 21420 56868 21422
rect 56700 21410 56756 21420
rect 56588 20078 56590 20130
rect 56642 20078 56644 20130
rect 56588 20066 56644 20078
rect 56700 20690 56756 20702
rect 56700 20638 56702 20690
rect 56754 20638 56756 20690
rect 56588 19906 56644 19918
rect 56588 19854 56590 19906
rect 56642 19854 56644 19906
rect 56588 18676 56644 19854
rect 56700 18788 56756 20638
rect 56812 20020 56868 21420
rect 56812 19954 56868 19964
rect 56700 18722 56756 18732
rect 56588 18610 56644 18620
rect 56252 17948 56420 18004
rect 56476 18452 56532 18462
rect 56252 16882 56308 17948
rect 56476 17108 56532 18396
rect 56924 17442 56980 25116
rect 57148 24724 57204 25566
rect 57484 26178 57540 26190
rect 57484 26126 57486 26178
rect 57538 26126 57540 26178
rect 57484 25508 57540 26126
rect 57148 24658 57204 24668
rect 57260 25452 57540 25508
rect 57820 25508 57876 25518
rect 57820 25506 58100 25508
rect 57820 25454 57822 25506
rect 57874 25454 58100 25506
rect 57820 25452 58100 25454
rect 57260 25396 57316 25452
rect 57820 25442 57876 25452
rect 57260 23938 57316 25340
rect 57484 24948 57540 24958
rect 57484 24854 57540 24892
rect 57820 24724 57876 24734
rect 57820 24630 57876 24668
rect 58044 24612 58100 25452
rect 58044 24518 58100 24556
rect 57260 23886 57262 23938
rect 57314 23886 57316 23938
rect 57260 22370 57316 23886
rect 57260 22318 57262 22370
rect 57314 22318 57316 22370
rect 57260 22306 57316 22318
rect 57932 23826 57988 23838
rect 57932 23774 57934 23826
rect 57986 23774 57988 23826
rect 57260 21588 57316 21598
rect 57484 21588 57540 21598
rect 57260 20802 57316 21532
rect 57260 20750 57262 20802
rect 57314 20750 57316 20802
rect 57260 19796 57316 20750
rect 57372 21586 57540 21588
rect 57372 21534 57486 21586
rect 57538 21534 57540 21586
rect 57372 21532 57540 21534
rect 57372 20914 57428 21532
rect 57484 21522 57540 21532
rect 57708 21588 57764 21598
rect 57708 21494 57764 21532
rect 57596 21476 57652 21486
rect 57596 21382 57652 21420
rect 57372 20862 57374 20914
rect 57426 20862 57428 20914
rect 57372 20132 57428 20862
rect 57596 21252 57652 21262
rect 57484 20132 57540 20142
rect 57372 20130 57540 20132
rect 57372 20078 57486 20130
rect 57538 20078 57540 20130
rect 57372 20076 57540 20078
rect 57484 20066 57540 20076
rect 57596 20018 57652 21196
rect 57932 20132 57988 23774
rect 58156 22148 58212 22158
rect 58156 22054 58212 22092
rect 58044 21586 58100 21598
rect 58044 21534 58046 21586
rect 58098 21534 58100 21586
rect 58044 20692 58100 21534
rect 58492 21588 58548 21598
rect 58492 21494 58548 21532
rect 58044 20626 58100 20636
rect 57596 19966 57598 20018
rect 57650 19966 57652 20018
rect 57596 19954 57652 19966
rect 57820 20020 57876 20030
rect 57820 19926 57876 19964
rect 57260 19730 57316 19740
rect 57932 19234 57988 20076
rect 58380 20468 58436 20478
rect 57932 19182 57934 19234
rect 57986 19182 57988 19234
rect 57932 19170 57988 19182
rect 58156 19908 58212 19918
rect 57372 18788 57428 18798
rect 56924 17390 56926 17442
rect 56978 17390 56980 17442
rect 56924 17378 56980 17390
rect 57036 17666 57092 17678
rect 57036 17614 57038 17666
rect 57090 17614 57092 17666
rect 56476 17042 56532 17052
rect 56364 16996 56420 17006
rect 56364 16902 56420 16940
rect 57036 16996 57092 17614
rect 57372 17668 57428 18732
rect 57708 18788 57764 18798
rect 57596 18676 57652 18686
rect 57596 18582 57652 18620
rect 57708 18674 57764 18732
rect 57708 18622 57710 18674
rect 57762 18622 57764 18674
rect 57708 18610 57764 18622
rect 57820 18564 57876 18574
rect 57820 18470 57876 18508
rect 57932 18450 57988 18462
rect 57932 18398 57934 18450
rect 57986 18398 57988 18450
rect 57372 17666 57876 17668
rect 57372 17614 57374 17666
rect 57426 17614 57876 17666
rect 57372 17612 57876 17614
rect 57372 17602 57428 17612
rect 57036 16930 57092 16940
rect 57260 17332 57316 17342
rect 56252 16830 56254 16882
rect 56306 16830 56308 16882
rect 56252 16818 56308 16830
rect 56140 16046 56142 16098
rect 56194 16046 56196 16098
rect 56140 16034 56196 16046
rect 56812 16660 56868 16670
rect 55692 15988 55748 15998
rect 55692 15538 55748 15932
rect 55692 15486 55694 15538
rect 55746 15486 55748 15538
rect 55692 15474 55748 15486
rect 56364 15540 56420 15550
rect 56364 15426 56420 15484
rect 56364 15374 56366 15426
rect 56418 15374 56420 15426
rect 55580 15316 55636 15326
rect 55580 15222 55636 15260
rect 55580 14644 55636 14654
rect 55468 14642 55636 14644
rect 55468 14590 55582 14642
rect 55634 14590 55636 14642
rect 55468 14588 55636 14590
rect 54684 14550 54740 14588
rect 55580 14578 55636 14588
rect 56252 14532 56308 14542
rect 56364 14532 56420 15374
rect 56700 15316 56756 15326
rect 54460 14478 54462 14530
rect 54514 14478 54516 14530
rect 54460 14466 54516 14478
rect 55804 14530 56420 14532
rect 55804 14478 56254 14530
rect 56306 14478 56420 14530
rect 56476 15260 56700 15316
rect 56476 14644 56532 15260
rect 56700 15222 56756 15260
rect 56476 14512 56532 14588
rect 55804 14476 56420 14478
rect 55356 13972 55412 13982
rect 55804 13972 55860 14476
rect 56252 14466 56308 14476
rect 55356 13970 55860 13972
rect 55356 13918 55358 13970
rect 55410 13918 55806 13970
rect 55858 13918 55860 13970
rect 55356 13916 55860 13918
rect 55356 13906 55412 13916
rect 55804 13906 55860 13916
rect 56588 13972 56644 13982
rect 53788 13860 53844 13870
rect 53788 13766 53844 13804
rect 54796 13524 54852 13534
rect 54796 13430 54852 13468
rect 55468 13524 55524 13534
rect 52668 13186 52836 13188
rect 52668 13134 52670 13186
rect 52722 13134 52836 13186
rect 52668 13132 52836 13134
rect 52668 13122 52724 13132
rect 50316 12898 50372 12908
rect 50988 12964 51044 12974
rect 52108 12944 52164 13020
rect 50204 12850 50260 12862
rect 50204 12798 50206 12850
rect 50258 12798 50260 12850
rect 50204 12740 50260 12798
rect 50764 12852 50820 12862
rect 50764 12758 50820 12796
rect 50204 12674 50260 12684
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 49756 12310 49812 12348
rect 49532 12292 49588 12302
rect 49308 12290 49588 12292
rect 49308 12238 49534 12290
rect 49586 12238 49588 12290
rect 49308 12236 49588 12238
rect 49532 12226 49588 12236
rect 50988 11394 51044 12908
rect 50988 11342 50990 11394
rect 51042 11342 51044 11394
rect 49532 11172 49588 11182
rect 48748 10704 48804 10780
rect 49196 10836 49252 10846
rect 48524 10098 48580 10108
rect 48300 9940 48356 9950
rect 48300 9846 48356 9884
rect 49196 9940 49252 10780
rect 49532 10724 49588 11116
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 49756 10836 49812 10846
rect 49756 10742 49812 10780
rect 49196 9826 49252 9884
rect 49420 10722 49588 10724
rect 49420 10670 49534 10722
rect 49586 10670 49588 10722
rect 49420 10668 49588 10670
rect 49420 9938 49476 10668
rect 49532 10658 49588 10668
rect 50988 10610 51044 11342
rect 50988 10558 50990 10610
rect 51042 10558 51044 10610
rect 50988 10546 51044 10558
rect 51324 12850 51380 12862
rect 51324 12798 51326 12850
rect 51378 12798 51380 12850
rect 51324 12740 51380 12798
rect 51324 11506 51380 12684
rect 53900 12290 53956 12302
rect 53900 12238 53902 12290
rect 53954 12238 53956 12290
rect 51324 11454 51326 11506
rect 51378 11454 51380 11506
rect 51324 10610 51380 11454
rect 53676 11954 53732 11966
rect 53676 11902 53678 11954
rect 53730 11902 53732 11954
rect 51660 11284 51716 11294
rect 51660 11190 51716 11228
rect 53116 11284 53172 11294
rect 51324 10558 51326 10610
rect 51378 10558 51380 10610
rect 51324 10546 51380 10558
rect 53116 10610 53172 11228
rect 53676 11284 53732 11902
rect 53676 11218 53732 11228
rect 53116 10558 53118 10610
rect 53170 10558 53172 10610
rect 53116 10546 53172 10558
rect 53340 10610 53396 10622
rect 53340 10558 53342 10610
rect 53394 10558 53396 10610
rect 51548 10498 51604 10510
rect 51548 10446 51550 10498
rect 51602 10446 51604 10498
rect 49868 10388 49924 10398
rect 49868 10294 49924 10332
rect 49420 9886 49422 9938
rect 49474 9886 49476 9938
rect 49420 9874 49476 9886
rect 49532 10164 49588 10174
rect 49196 9774 49198 9826
rect 49250 9774 49252 9826
rect 49196 9762 49252 9774
rect 47180 9044 47236 9054
rect 47404 9024 47460 9100
rect 47628 9156 47684 9166
rect 47628 9062 47684 9100
rect 49084 9156 49140 9166
rect 47740 9042 47796 9054
rect 47180 8950 47236 8988
rect 47740 8990 47742 9042
rect 47794 8990 47796 9042
rect 46956 8206 46958 8258
rect 47010 8206 47012 8258
rect 46956 8194 47012 8206
rect 47068 8372 47124 8382
rect 46956 7588 47012 7598
rect 47068 7588 47124 8316
rect 47740 8372 47796 8990
rect 47740 8306 47796 8316
rect 49084 8258 49140 9100
rect 49084 8206 49086 8258
rect 49138 8206 49140 8258
rect 49084 8194 49140 8206
rect 49532 9154 49588 10108
rect 51548 9828 51604 10446
rect 53340 10500 53396 10558
rect 51660 10388 51716 10398
rect 51660 9938 51716 10332
rect 51660 9886 51662 9938
rect 51714 9886 51716 9938
rect 51660 9874 51716 9886
rect 51548 9762 51604 9772
rect 52108 9828 52164 9838
rect 49868 9716 49924 9726
rect 49868 9622 49924 9660
rect 50428 9716 50484 9726
rect 49532 9102 49534 9154
rect 49586 9102 49588 9154
rect 49532 8258 49588 9102
rect 49756 9156 49812 9166
rect 49756 9062 49812 9100
rect 50428 9156 50484 9660
rect 50876 9604 50932 9614
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 50876 9268 50932 9548
rect 51548 9604 51604 9614
rect 51548 9510 51604 9548
rect 49868 8818 49924 8830
rect 49868 8766 49870 8818
rect 49922 8766 49924 8818
rect 49868 8428 49924 8766
rect 49868 8372 50036 8428
rect 49532 8206 49534 8258
rect 49586 8206 49588 8258
rect 49532 8194 49588 8206
rect 46956 7586 47124 7588
rect 46956 7534 46958 7586
rect 47010 7534 47124 7586
rect 46956 7532 47124 7534
rect 47852 8146 47908 8158
rect 47852 8094 47854 8146
rect 47906 8094 47908 8146
rect 46956 7522 47012 7532
rect 46508 7422 46510 7474
rect 46562 7422 46564 7474
rect 46508 7410 46564 7422
rect 45388 6466 45444 6478
rect 45388 6414 45390 6466
rect 45442 6414 45444 6466
rect 45276 6132 45332 6142
rect 45388 6132 45444 6414
rect 45332 6076 45444 6132
rect 45276 6000 45332 6076
rect 45500 6020 45556 6030
rect 45500 5926 45556 5964
rect 46284 6020 46340 6030
rect 46284 5926 46340 5964
rect 47068 6020 47124 6058
rect 47068 5954 47124 5964
rect 45164 5906 45220 5918
rect 45164 5854 45166 5906
rect 45218 5854 45220 5906
rect 45164 5684 45220 5854
rect 44604 5628 45220 5684
rect 45388 5908 45444 5918
rect 46172 5908 46228 5918
rect 44604 5122 44660 5628
rect 45388 5348 45444 5852
rect 45948 5852 46172 5908
rect 45500 5348 45556 5358
rect 45388 5346 45556 5348
rect 45388 5294 45502 5346
rect 45554 5294 45556 5346
rect 45388 5292 45556 5294
rect 45500 5282 45556 5292
rect 45836 5236 45892 5246
rect 45836 5142 45892 5180
rect 44604 5070 44606 5122
rect 44658 5070 44660 5122
rect 44604 5058 44660 5070
rect 44380 4722 44436 4732
rect 44492 5012 44548 5022
rect 44492 4564 44548 4956
rect 44716 5012 44772 5022
rect 44716 5010 44884 5012
rect 44716 4958 44718 5010
rect 44770 4958 44884 5010
rect 44716 4956 44884 4958
rect 44716 4946 44772 4956
rect 44044 4452 44100 4462
rect 43932 4450 44100 4452
rect 43932 4398 44046 4450
rect 44098 4398 44100 4450
rect 43932 4396 44100 4398
rect 44044 4386 44100 4396
rect 44492 4338 44548 4508
rect 44492 4286 44494 4338
rect 44546 4286 44548 4338
rect 44492 4274 44548 4286
rect 44828 4452 44884 4956
rect 45724 4898 45780 4910
rect 45724 4846 45726 4898
rect 45778 4846 45780 4898
rect 45724 4788 45780 4846
rect 45724 4722 45780 4732
rect 45724 4564 45780 4574
rect 45724 4470 45780 4508
rect 45948 4562 46004 5852
rect 46172 5814 46228 5852
rect 46956 5908 47012 5918
rect 46956 5814 47012 5852
rect 47852 5906 47908 8094
rect 49756 8146 49812 8158
rect 49756 8094 49758 8146
rect 49810 8094 49812 8146
rect 49756 8036 49812 8094
rect 49756 7970 49812 7980
rect 49644 7700 49700 7710
rect 48636 6468 48692 6478
rect 47964 6132 48020 6142
rect 47964 6038 48020 6076
rect 47852 5854 47854 5906
rect 47906 5854 47908 5906
rect 46284 5684 46340 5694
rect 46284 5590 46340 5628
rect 47292 5684 47348 5694
rect 47292 5234 47348 5628
rect 47292 5182 47294 5234
rect 47346 5182 47348 5234
rect 47292 5170 47348 5182
rect 47740 5124 47796 5134
rect 47852 5124 47908 5854
rect 48524 5348 48580 5358
rect 47740 5122 47908 5124
rect 47740 5070 47742 5122
rect 47794 5070 47908 5122
rect 47740 5068 47908 5070
rect 48076 5236 48132 5246
rect 47740 5058 47796 5068
rect 45948 4510 45950 4562
rect 46002 4510 46004 4562
rect 45948 4498 46004 4510
rect 42588 4174 42590 4226
rect 42642 4174 42644 4226
rect 42588 4162 42644 4174
rect 44828 4226 44884 4396
rect 45612 4452 45668 4462
rect 45612 4358 45668 4396
rect 48076 4338 48132 5180
rect 48076 4286 48078 4338
rect 48130 4286 48132 4338
rect 48076 4274 48132 4286
rect 48188 5124 48244 5134
rect 48188 5010 48244 5068
rect 48188 4958 48190 5010
rect 48242 4958 48244 5010
rect 48188 4340 48244 4958
rect 48300 4340 48356 4350
rect 48188 4338 48356 4340
rect 48188 4286 48302 4338
rect 48354 4286 48356 4338
rect 48188 4284 48356 4286
rect 48300 4274 48356 4284
rect 48524 4338 48580 5292
rect 48636 4450 48692 6412
rect 48748 6244 48804 6254
rect 48748 5348 48804 6188
rect 48748 5234 48804 5292
rect 49644 5346 49700 7644
rect 49980 7474 50036 8372
rect 50428 7700 50484 9100
rect 50764 9212 50932 9268
rect 50652 9044 50708 9054
rect 50652 8036 50708 8988
rect 50764 8146 50820 9212
rect 51660 9156 51716 9166
rect 51660 9062 51716 9100
rect 51548 9044 51604 9054
rect 51548 8950 51604 8988
rect 51884 9042 51940 9054
rect 51884 8990 51886 9042
rect 51938 8990 51940 9042
rect 50988 8818 51044 8830
rect 50988 8766 50990 8818
rect 51042 8766 51044 8818
rect 50988 8428 51044 8766
rect 50876 8372 51044 8428
rect 51100 8820 51156 8830
rect 50876 8260 50932 8372
rect 51100 8260 51156 8764
rect 51884 8372 51940 8990
rect 51884 8306 51940 8316
rect 50876 8194 50932 8204
rect 50988 8258 51156 8260
rect 50988 8206 51102 8258
rect 51154 8206 51156 8258
rect 50988 8204 51156 8206
rect 50764 8094 50766 8146
rect 50818 8094 50820 8146
rect 50764 8082 50820 8094
rect 50652 7970 50708 7980
rect 50876 8036 50932 8046
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 50428 7644 50708 7700
rect 50652 7586 50708 7644
rect 50652 7534 50654 7586
rect 50706 7534 50708 7586
rect 50652 7522 50708 7534
rect 49980 7422 49982 7474
rect 50034 7422 50036 7474
rect 49980 7410 50036 7422
rect 50876 7474 50932 7980
rect 50876 7422 50878 7474
rect 50930 7422 50932 7474
rect 50876 7410 50932 7422
rect 50988 7362 51044 8204
rect 51100 8194 51156 8204
rect 52108 8258 52164 9772
rect 52780 9828 52836 9838
rect 52780 9042 52836 9772
rect 52780 8990 52782 9042
rect 52834 8990 52836 9042
rect 52780 8978 52836 8990
rect 53004 9044 53060 9054
rect 53340 9044 53396 10444
rect 53900 10500 53956 12238
rect 55468 12180 55524 13468
rect 56476 12964 56532 12974
rect 56140 12962 56532 12964
rect 56140 12910 56478 12962
rect 56530 12910 56532 12962
rect 56140 12908 56532 12910
rect 56028 12292 56084 12302
rect 56028 12198 56084 12236
rect 55580 12180 55636 12190
rect 55468 12124 55580 12180
rect 54012 11956 54068 11966
rect 54012 11954 54964 11956
rect 54012 11902 54014 11954
rect 54066 11902 54964 11954
rect 54012 11900 54964 11902
rect 54012 11890 54068 11900
rect 53900 10434 53956 10444
rect 54012 11394 54068 11406
rect 54012 11342 54014 11394
rect 54066 11342 54068 11394
rect 54012 10498 54068 11342
rect 54908 11394 54964 11900
rect 55468 11788 55524 12124
rect 55580 12048 55636 12124
rect 56140 12068 56196 12908
rect 56476 12898 56532 12908
rect 54908 11342 54910 11394
rect 54962 11342 54964 11394
rect 54908 11330 54964 11342
rect 55356 11732 55524 11788
rect 56028 12012 56196 12068
rect 56252 12738 56308 12750
rect 56252 12686 56254 12738
rect 56306 12686 56308 12738
rect 55356 11394 55412 11676
rect 55356 11342 55358 11394
rect 55410 11342 55412 11394
rect 55356 11330 55412 11342
rect 54012 10446 54014 10498
rect 54066 10446 54068 10498
rect 54012 10276 54068 10446
rect 54124 11282 54180 11294
rect 54124 11230 54126 11282
rect 54178 11230 54180 11282
rect 54124 10388 54180 11230
rect 54684 11284 54740 11294
rect 54684 11190 54740 11228
rect 54796 11172 54852 11182
rect 54796 10610 54852 11116
rect 56028 11172 56084 12012
rect 56028 11106 56084 11116
rect 56140 11844 56196 11854
rect 55804 10724 55860 10734
rect 55804 10722 55972 10724
rect 55804 10670 55806 10722
rect 55858 10670 55972 10722
rect 55804 10668 55972 10670
rect 55804 10658 55860 10668
rect 54796 10558 54798 10610
rect 54850 10558 54852 10610
rect 54796 10546 54852 10558
rect 55692 10610 55748 10622
rect 55692 10558 55694 10610
rect 55746 10558 55748 10610
rect 54572 10500 54628 10510
rect 54572 10406 54628 10444
rect 54124 10322 54180 10332
rect 54460 10388 54516 10398
rect 54012 10210 54068 10220
rect 54348 9826 54404 9838
rect 54348 9774 54350 9826
rect 54402 9774 54404 9826
rect 53676 9156 53732 9166
rect 53676 9062 53732 9100
rect 54348 9156 54404 9774
rect 53004 9042 53396 9044
rect 53004 8990 53006 9042
rect 53058 8990 53396 9042
rect 53004 8988 53396 8990
rect 53564 9044 53620 9054
rect 53004 8820 53060 8988
rect 53004 8754 53060 8764
rect 53228 8372 53284 8382
rect 52108 8206 52110 8258
rect 52162 8206 52164 8258
rect 52108 8194 52164 8206
rect 52668 8260 52724 8270
rect 52668 8166 52724 8204
rect 53116 8148 53172 8158
rect 53116 7586 53172 8092
rect 53228 7698 53284 8316
rect 53452 8372 53508 8382
rect 53452 8258 53508 8316
rect 53452 8206 53454 8258
rect 53506 8206 53508 8258
rect 53452 8194 53508 8206
rect 53228 7646 53230 7698
rect 53282 7646 53284 7698
rect 53228 7634 53284 7646
rect 53452 7700 53508 7710
rect 53564 7700 53620 8988
rect 54236 9044 54292 9054
rect 54236 8950 54292 8988
rect 54236 8258 54292 8270
rect 54236 8206 54238 8258
rect 54290 8206 54292 8258
rect 53676 8148 53732 8158
rect 53676 8054 53732 8092
rect 53452 7698 53620 7700
rect 53452 7646 53454 7698
rect 53506 7646 53620 7698
rect 53452 7644 53620 7646
rect 53452 7634 53508 7644
rect 53116 7534 53118 7586
rect 53170 7534 53172 7586
rect 53116 7522 53172 7534
rect 50988 7310 50990 7362
rect 51042 7310 51044 7362
rect 50988 7298 51044 7310
rect 53788 7364 53844 7374
rect 54236 7364 54292 8206
rect 54348 7586 54404 9100
rect 54460 9154 54516 10332
rect 55132 10388 55188 10398
rect 55132 10386 55300 10388
rect 55132 10334 55134 10386
rect 55186 10334 55300 10386
rect 55132 10332 55300 10334
rect 55132 10322 55188 10332
rect 54796 10276 54852 10286
rect 54460 9102 54462 9154
rect 54514 9102 54516 9154
rect 54460 9090 54516 9102
rect 54572 9826 54628 9838
rect 54572 9774 54574 9826
rect 54626 9774 54628 9826
rect 54572 9604 54628 9774
rect 54572 8428 54628 9548
rect 54684 9268 54740 9278
rect 54684 9174 54740 9212
rect 54796 9154 54852 10220
rect 54796 9102 54798 9154
rect 54850 9102 54852 9154
rect 54796 9090 54852 9102
rect 55132 10164 55188 10174
rect 54460 8372 54628 8428
rect 55020 8484 55076 8494
rect 55132 8484 55188 10108
rect 55244 9826 55300 10332
rect 55468 10052 55524 10062
rect 55468 9958 55524 9996
rect 55244 9774 55246 9826
rect 55298 9774 55300 9826
rect 55244 9762 55300 9774
rect 55692 9268 55748 10558
rect 55020 8482 55188 8484
rect 55020 8430 55022 8482
rect 55074 8430 55188 8482
rect 55020 8428 55188 8430
rect 55356 9156 55412 9166
rect 55020 8418 55076 8428
rect 54460 7698 54516 8372
rect 54684 8260 54740 8270
rect 54684 8166 54740 8204
rect 54460 7646 54462 7698
rect 54514 7646 54516 7698
rect 54460 7634 54516 7646
rect 54684 7700 54740 7710
rect 55356 7700 55412 9100
rect 55580 8148 55636 8158
rect 54684 7698 55412 7700
rect 54684 7646 54686 7698
rect 54738 7646 55412 7698
rect 54684 7644 55412 7646
rect 54684 7634 54740 7644
rect 54348 7534 54350 7586
rect 54402 7534 54404 7586
rect 54348 7522 54404 7534
rect 55356 7474 55412 7644
rect 55356 7422 55358 7474
rect 55410 7422 55412 7474
rect 55356 7410 55412 7422
rect 55468 8146 55636 8148
rect 55468 8094 55582 8146
rect 55634 8094 55636 8146
rect 55468 8092 55636 8094
rect 53788 7362 54292 7364
rect 53788 7310 53790 7362
rect 53842 7310 54292 7362
rect 53788 7308 54292 7310
rect 53788 6580 53844 7308
rect 55468 6692 55524 8092
rect 55580 8082 55636 8092
rect 55580 7476 55636 7486
rect 55692 7476 55748 9212
rect 55804 10052 55860 10062
rect 55804 8932 55860 9996
rect 55916 9156 55972 10668
rect 56028 10610 56084 10622
rect 56028 10558 56030 10610
rect 56082 10558 56084 10610
rect 56028 9828 56084 10558
rect 56028 9762 56084 9772
rect 56140 10052 56196 11788
rect 56252 11284 56308 12686
rect 56364 12738 56420 12750
rect 56364 12686 56366 12738
rect 56418 12686 56420 12738
rect 56364 12180 56420 12686
rect 56588 12402 56644 13916
rect 56588 12350 56590 12402
rect 56642 12350 56644 12402
rect 56588 12338 56644 12350
rect 56476 12180 56532 12190
rect 56364 12178 56532 12180
rect 56364 12126 56478 12178
rect 56530 12126 56532 12178
rect 56364 12124 56532 12126
rect 56476 12114 56532 12124
rect 56812 11844 56868 16604
rect 57260 15428 57316 17276
rect 57820 16994 57876 17612
rect 57820 16942 57822 16994
rect 57874 16942 57876 16994
rect 57820 16930 57876 16942
rect 57484 16660 57540 16670
rect 57260 14642 57316 15372
rect 57372 16658 57540 16660
rect 57372 16606 57486 16658
rect 57538 16606 57540 16658
rect 57372 16604 57540 16606
rect 57372 14868 57428 16604
rect 57484 16594 57540 16604
rect 57596 16660 57652 16670
rect 57596 16566 57652 16604
rect 57932 16548 57988 18398
rect 58156 16994 58212 19852
rect 58380 19234 58436 20412
rect 58380 19182 58382 19234
rect 58434 19182 58436 19234
rect 58380 19170 58436 19182
rect 58604 18788 58660 51212
rect 58604 18722 58660 18732
rect 58716 28756 58772 28766
rect 58268 18226 58324 18238
rect 58268 18174 58270 18226
rect 58322 18174 58324 18226
rect 58268 17106 58324 18174
rect 58268 17054 58270 17106
rect 58322 17054 58324 17106
rect 58268 17042 58324 17054
rect 58380 17108 58436 17118
rect 58156 16942 58158 16994
rect 58210 16942 58212 16994
rect 58156 16930 58212 16942
rect 58380 16994 58436 17052
rect 58380 16942 58382 16994
rect 58434 16942 58436 16994
rect 58380 16930 58436 16942
rect 57708 16492 57988 16548
rect 57708 16436 57764 16492
rect 57484 16380 57764 16436
rect 57484 15426 57540 16380
rect 58492 16098 58548 16110
rect 58492 16046 58494 16098
rect 58546 16046 58548 16098
rect 57484 15374 57486 15426
rect 57538 15374 57540 15426
rect 57484 15362 57540 15374
rect 57820 15986 57876 15998
rect 57820 15934 57822 15986
rect 57874 15934 57876 15986
rect 57596 15316 57652 15326
rect 57596 15222 57652 15260
rect 57372 14812 57540 14868
rect 57260 14590 57262 14642
rect 57314 14590 57316 14642
rect 57260 14578 57316 14590
rect 56476 11788 56868 11844
rect 56924 12292 56980 12302
rect 56476 11506 56532 11788
rect 56476 11454 56478 11506
rect 56530 11454 56532 11506
rect 56476 11442 56532 11454
rect 56252 11218 56308 11228
rect 56588 11284 56644 11294
rect 56588 11190 56644 11228
rect 56364 11172 56420 11182
rect 56364 10276 56420 11116
rect 56364 10210 56420 10220
rect 56924 10052 56980 12236
rect 57372 12180 57428 12190
rect 57036 12178 57428 12180
rect 57036 12126 57374 12178
rect 57426 12126 57428 12178
rect 57036 12124 57428 12126
rect 57036 11394 57092 12124
rect 57372 12114 57428 12124
rect 57484 12068 57540 14812
rect 57820 13972 57876 15934
rect 57932 15428 57988 15438
rect 57932 15314 57988 15372
rect 57932 15262 57934 15314
rect 57986 15262 57988 15314
rect 57932 15250 57988 15262
rect 57820 13906 57876 13916
rect 58492 14306 58548 16046
rect 58716 15540 58772 28700
rect 58716 15474 58772 15484
rect 58492 14254 58494 14306
rect 58546 14254 58548 14306
rect 57596 12292 57652 12302
rect 57596 12198 57652 12236
rect 57708 12180 57764 12190
rect 57708 12086 57764 12124
rect 57484 12012 57652 12068
rect 57036 11342 57038 11394
rect 57090 11342 57092 11394
rect 57036 11330 57092 11342
rect 57148 11956 57204 11966
rect 57148 11172 57204 11900
rect 56140 9996 56868 10052
rect 55916 9090 55972 9100
rect 56028 9042 56084 9054
rect 56028 8990 56030 9042
rect 56082 8990 56084 9042
rect 56028 8932 56084 8990
rect 55804 8876 56084 8932
rect 56140 8932 56196 9996
rect 56812 9938 56868 9996
rect 56812 9886 56814 9938
rect 56866 9886 56868 9938
rect 56812 9874 56868 9886
rect 56924 9826 56980 9996
rect 56924 9774 56926 9826
rect 56978 9774 56980 9826
rect 56924 9762 56980 9774
rect 57036 11116 57204 11172
rect 56252 8932 56308 8942
rect 56140 8930 56308 8932
rect 56140 8878 56254 8930
rect 56306 8878 56308 8930
rect 56140 8876 56308 8878
rect 56252 8866 56308 8876
rect 56700 8930 56756 8942
rect 56700 8878 56702 8930
rect 56754 8878 56756 8930
rect 56700 8428 56756 8878
rect 56588 8372 56756 8428
rect 56924 8484 56980 8494
rect 57036 8484 57092 11116
rect 57484 9938 57540 9950
rect 57484 9886 57486 9938
rect 57538 9886 57540 9938
rect 57484 9154 57540 9886
rect 57596 9266 57652 12012
rect 58492 11956 58548 14254
rect 58492 11890 58548 11900
rect 57596 9214 57598 9266
rect 57650 9214 57652 9266
rect 57596 9202 57652 9214
rect 57708 11172 57764 11182
rect 57484 9102 57486 9154
rect 57538 9102 57540 9154
rect 57484 9090 57540 9102
rect 57708 9154 57764 11116
rect 57708 9102 57710 9154
rect 57762 9102 57764 9154
rect 57708 9090 57764 9102
rect 58044 9828 58100 9838
rect 58044 9042 58100 9772
rect 58044 8990 58046 9042
rect 58098 8990 58100 9042
rect 58044 8978 58100 8990
rect 56924 8482 57092 8484
rect 56924 8430 56926 8482
rect 56978 8430 57092 8482
rect 56924 8428 57092 8430
rect 57932 8818 57988 8830
rect 57932 8766 57934 8818
rect 57986 8766 57988 8818
rect 57932 8428 57988 8766
rect 56924 8418 56980 8428
rect 57708 8372 57988 8428
rect 56588 8370 56644 8372
rect 56588 8318 56590 8370
rect 56642 8318 56644 8370
rect 56588 8306 56644 8318
rect 55916 8258 55972 8270
rect 55916 8206 55918 8258
rect 55970 8206 55972 8258
rect 55916 7698 55972 8206
rect 55916 7646 55918 7698
rect 55970 7646 55972 7698
rect 55916 7634 55972 7646
rect 56700 8258 56756 8270
rect 56700 8206 56702 8258
rect 56754 8206 56756 8258
rect 55580 7474 55748 7476
rect 55580 7422 55582 7474
rect 55634 7422 55748 7474
rect 55580 7420 55748 7422
rect 55580 7410 55636 7420
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 53788 6132 53844 6524
rect 55020 6636 55524 6692
rect 55020 6468 55076 6636
rect 56700 6580 56756 8206
rect 57708 8034 57764 8372
rect 57708 7982 57710 8034
rect 57762 7982 57764 8034
rect 57708 7700 57764 7982
rect 57708 7634 57764 7644
rect 56700 6514 56756 6524
rect 55020 6374 55076 6412
rect 55468 6468 55524 6478
rect 55468 6374 55524 6412
rect 53788 6066 53844 6076
rect 49644 5294 49646 5346
rect 49698 5294 49700 5346
rect 49644 5282 49700 5294
rect 48748 5182 48750 5234
rect 48802 5182 48804 5234
rect 48748 5170 48804 5182
rect 49196 5236 49252 5246
rect 49196 5142 49252 5180
rect 48972 5124 49028 5134
rect 48972 5030 49028 5068
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 48636 4398 48638 4450
rect 48690 4398 48692 4450
rect 48636 4386 48692 4398
rect 48524 4286 48526 4338
rect 48578 4286 48580 4338
rect 48524 4274 48580 4286
rect 44828 4174 44830 4226
rect 44882 4174 44884 4226
rect 44828 4162 44884 4174
rect 47516 3780 47572 3790
rect 47516 3666 47572 3724
rect 47516 3614 47518 3666
rect 47570 3614 47572 3666
rect 47516 3602 47572 3614
rect 42140 3502 42142 3554
rect 42194 3502 42196 3554
rect 42140 3490 42196 3502
rect 42028 3378 42084 3388
rect 48076 3444 48132 3454
rect 39004 3332 39060 3342
rect 38780 3330 39060 3332
rect 38780 3278 39006 3330
rect 39058 3278 39060 3330
rect 38780 3276 39060 3278
rect 37212 3266 37268 3276
rect 38780 800 38836 3276
rect 39004 3266 39060 3276
rect 48076 3330 48132 3388
rect 48748 3444 48804 3454
rect 48748 3350 48804 3388
rect 55692 3444 55748 3454
rect 56028 3444 56084 3454
rect 55692 3442 56028 3444
rect 55692 3390 55694 3442
rect 55746 3390 56028 3442
rect 55692 3388 56028 3390
rect 55692 3378 55748 3388
rect 48076 3278 48078 3330
rect 48130 3278 48132 3330
rect 47404 2994 47460 3006
rect 47404 2942 47406 2994
rect 47458 2942 47460 2994
rect 47404 800 47460 2942
rect 48076 2994 48132 3278
rect 55356 3332 55412 3342
rect 55356 3238 55412 3276
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 48076 2942 48078 2994
rect 48130 2942 48132 2994
rect 48076 2930 48132 2942
rect 56028 800 56084 3388
rect 56588 3444 56644 3454
rect 56588 3350 56644 3388
rect 4256 0 4368 800
rect 12880 0 12992 800
rect 21504 0 21616 800
rect 30128 0 30240 800
rect 38752 0 38864 800
rect 47376 0 47488 800
rect 56000 0 56112 800
<< via2 >>
rect 1372 60732 1428 60788
rect 1148 56924 1204 56980
rect 1036 52332 1092 52388
rect 924 49868 980 49924
rect 1036 43260 1092 43316
rect 924 40012 980 40068
rect 1036 33852 1092 33908
rect 1036 23324 1092 23380
rect 1260 52220 1316 52276
rect 1260 48524 1316 48580
rect 1708 60620 1764 60676
rect 1484 55916 1540 55972
rect 4476 60394 4532 60396
rect 4476 60342 4478 60394
rect 4478 60342 4530 60394
rect 4530 60342 4532 60394
rect 4476 60340 4532 60342
rect 4580 60394 4636 60396
rect 4580 60342 4582 60394
rect 4582 60342 4634 60394
rect 4634 60342 4636 60394
rect 4580 60340 4636 60342
rect 4684 60394 4740 60396
rect 4684 60342 4686 60394
rect 4686 60342 4738 60394
rect 4738 60342 4740 60394
rect 4684 60340 4740 60342
rect 25340 60844 25396 60900
rect 4620 60002 4676 60004
rect 4620 59950 4622 60002
rect 4622 59950 4674 60002
rect 4674 59950 4676 60002
rect 4620 59948 4676 59950
rect 4956 59948 5012 60004
rect 3724 59778 3780 59780
rect 3724 59726 3726 59778
rect 3726 59726 3778 59778
rect 3778 59726 3780 59778
rect 3724 59724 3780 59726
rect 2716 58940 2772 58996
rect 2492 58268 2548 58324
rect 1596 52220 1652 52276
rect 1708 55356 1764 55412
rect 3612 58940 3668 58996
rect 4620 59442 4676 59444
rect 4620 59390 4622 59442
rect 4622 59390 4674 59442
rect 4674 59390 4676 59442
rect 4620 59388 4676 59390
rect 4060 58940 4116 58996
rect 3388 58210 3444 58212
rect 3388 58158 3390 58210
rect 3390 58158 3442 58210
rect 3442 58158 3444 58210
rect 3388 58156 3444 58158
rect 2940 57708 2996 57764
rect 2156 56252 2212 56308
rect 2380 57260 2436 57316
rect 2380 55804 2436 55860
rect 2380 55580 2436 55636
rect 2268 55468 2324 55524
rect 1820 54626 1876 54628
rect 1820 54574 1822 54626
rect 1822 54574 1874 54626
rect 1874 54574 1876 54626
rect 1820 54572 1876 54574
rect 1932 53900 1988 53956
rect 2044 53618 2100 53620
rect 2044 53566 2046 53618
rect 2046 53566 2098 53618
rect 2098 53566 2100 53618
rect 2044 53564 2100 53566
rect 2716 56306 2772 56308
rect 2716 56254 2718 56306
rect 2718 56254 2770 56306
rect 2770 56254 2772 56306
rect 2716 56252 2772 56254
rect 2940 56252 2996 56308
rect 3164 57596 3220 57652
rect 4060 57874 4116 57876
rect 4060 57822 4062 57874
rect 4062 57822 4114 57874
rect 4114 57822 4116 57874
rect 4060 57820 4116 57822
rect 4844 59052 4900 59108
rect 4476 58826 4532 58828
rect 4476 58774 4478 58826
rect 4478 58774 4530 58826
rect 4530 58774 4532 58826
rect 4476 58772 4532 58774
rect 4580 58826 4636 58828
rect 4580 58774 4582 58826
rect 4582 58774 4634 58826
rect 4634 58774 4636 58826
rect 4580 58772 4636 58774
rect 4684 58826 4740 58828
rect 4684 58774 4686 58826
rect 4686 58774 4738 58826
rect 4738 58774 4740 58826
rect 4684 58772 4740 58774
rect 3724 57538 3780 57540
rect 3724 57486 3726 57538
rect 3726 57486 3778 57538
rect 3778 57486 3780 57538
rect 3724 57484 3780 57486
rect 3500 56642 3556 56644
rect 3500 56590 3502 56642
rect 3502 56590 3554 56642
rect 3554 56590 3556 56642
rect 3500 56588 3556 56590
rect 3164 55970 3220 55972
rect 3164 55918 3166 55970
rect 3166 55918 3218 55970
rect 3218 55918 3220 55970
rect 3164 55916 3220 55918
rect 3052 55580 3108 55636
rect 3388 55804 3444 55860
rect 2604 55244 2660 55300
rect 2828 55132 2884 55188
rect 2604 54796 2660 54852
rect 1820 52274 1876 52276
rect 1820 52222 1822 52274
rect 1822 52222 1874 52274
rect 1874 52222 1876 52274
rect 1820 52220 1876 52222
rect 1932 51884 1988 51940
rect 2380 53004 2436 53060
rect 2156 52668 2212 52724
rect 2268 51884 2324 51940
rect 1932 51266 1988 51268
rect 1932 51214 1934 51266
rect 1934 51214 1986 51266
rect 1986 51214 1988 51266
rect 1932 51212 1988 51214
rect 2156 50594 2212 50596
rect 2156 50542 2158 50594
rect 2158 50542 2210 50594
rect 2210 50542 2212 50594
rect 2156 50540 2212 50542
rect 1820 50428 1876 50484
rect 1484 48188 1540 48244
rect 1596 49196 1652 49252
rect 1372 42812 1428 42868
rect 1372 38780 1428 38836
rect 1596 47628 1652 47684
rect 2044 48636 2100 48692
rect 2380 49810 2436 49812
rect 2380 49758 2382 49810
rect 2382 49758 2434 49810
rect 2434 49758 2436 49810
rect 2380 49756 2436 49758
rect 2268 48412 2324 48468
rect 2380 48300 2436 48356
rect 2268 47292 2324 47348
rect 2380 46956 2436 47012
rect 2156 46732 2212 46788
rect 1820 46396 1876 46452
rect 1932 46060 1988 46116
rect 2716 54738 2772 54740
rect 2716 54686 2718 54738
rect 2718 54686 2770 54738
rect 2770 54686 2772 54738
rect 2716 54684 2772 54686
rect 2716 53116 2772 53172
rect 3612 55580 3668 55636
rect 3724 55020 3780 55076
rect 3276 53842 3332 53844
rect 3276 53790 3278 53842
rect 3278 53790 3330 53842
rect 3330 53790 3332 53842
rect 3276 53788 3332 53790
rect 3164 53676 3220 53732
rect 2940 53340 2996 53396
rect 3052 53452 3108 53508
rect 2828 52892 2884 52948
rect 2940 53116 2996 53172
rect 2604 51938 2660 51940
rect 2604 51886 2606 51938
rect 2606 51886 2658 51938
rect 2658 51886 2660 51938
rect 2604 51884 2660 51886
rect 2604 50706 2660 50708
rect 2604 50654 2606 50706
rect 2606 50654 2658 50706
rect 2658 50654 2660 50706
rect 2604 50652 2660 50654
rect 3164 53340 3220 53396
rect 3052 52780 3108 52836
rect 3164 52220 3220 52276
rect 3276 52892 3332 52948
rect 3052 52108 3108 52164
rect 2940 50092 2996 50148
rect 2940 49698 2996 49700
rect 2940 49646 2942 49698
rect 2942 49646 2994 49698
rect 2994 49646 2996 49698
rect 2940 49644 2996 49646
rect 4060 56028 4116 56084
rect 4060 55580 4116 55636
rect 3948 55074 4004 55076
rect 3948 55022 3950 55074
rect 3950 55022 4002 55074
rect 4002 55022 4004 55074
rect 3948 55020 4004 55022
rect 4508 57932 4564 57988
rect 4620 57538 4676 57540
rect 4620 57486 4622 57538
rect 4622 57486 4674 57538
rect 4674 57486 4676 57538
rect 4620 57484 4676 57486
rect 4508 57372 4564 57428
rect 4476 57258 4532 57260
rect 4476 57206 4478 57258
rect 4478 57206 4530 57258
rect 4530 57206 4532 57258
rect 4476 57204 4532 57206
rect 4580 57258 4636 57260
rect 4580 57206 4582 57258
rect 4582 57206 4634 57258
rect 4634 57206 4636 57258
rect 4580 57204 4636 57206
rect 4684 57258 4740 57260
rect 4684 57206 4686 57258
rect 4686 57206 4738 57258
rect 4738 57206 4740 57258
rect 4684 57204 4740 57206
rect 9772 60002 9828 60004
rect 9772 59950 9774 60002
rect 9774 59950 9826 60002
rect 9826 59950 9828 60002
rect 9772 59948 9828 59950
rect 5068 59890 5124 59892
rect 5068 59838 5070 59890
rect 5070 59838 5122 59890
rect 5122 59838 5124 59890
rect 5068 59836 5124 59838
rect 5852 59836 5908 59892
rect 6300 59890 6356 59892
rect 6300 59838 6302 59890
rect 6302 59838 6354 59890
rect 6354 59838 6356 59890
rect 6300 59836 6356 59838
rect 7644 59836 7700 59892
rect 5740 59388 5796 59444
rect 5068 59330 5124 59332
rect 5068 59278 5070 59330
rect 5070 59278 5122 59330
rect 5122 59278 5124 59330
rect 5068 59276 5124 59278
rect 4956 57820 5012 57876
rect 5068 57538 5124 57540
rect 5068 57486 5070 57538
rect 5070 57486 5122 57538
rect 5122 57486 5124 57538
rect 5068 57484 5124 57486
rect 4284 56642 4340 56644
rect 4284 56590 4286 56642
rect 4286 56590 4338 56642
rect 4338 56590 4340 56642
rect 4284 56588 4340 56590
rect 4620 55970 4676 55972
rect 4620 55918 4622 55970
rect 4622 55918 4674 55970
rect 4674 55918 4676 55970
rect 4620 55916 4676 55918
rect 4732 55804 4788 55860
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 5180 56588 5236 56644
rect 5068 55804 5124 55860
rect 5068 55468 5124 55524
rect 4844 55244 4900 55300
rect 4172 54908 4228 54964
rect 4844 55074 4900 55076
rect 4844 55022 4846 55074
rect 4846 55022 4898 55074
rect 4898 55022 4900 55074
rect 4844 55020 4900 55022
rect 4396 54908 4452 54964
rect 4396 54514 4452 54516
rect 4396 54462 4398 54514
rect 4398 54462 4450 54514
rect 4450 54462 4452 54514
rect 4396 54460 4452 54462
rect 4956 54514 5012 54516
rect 4956 54462 4958 54514
rect 4958 54462 5010 54514
rect 5010 54462 5012 54514
rect 4956 54460 5012 54462
rect 3948 54402 4004 54404
rect 3948 54350 3950 54402
rect 3950 54350 4002 54402
rect 4002 54350 4004 54402
rect 3948 54348 4004 54350
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 4508 53900 4564 53956
rect 4284 53788 4340 53844
rect 3724 53228 3780 53284
rect 3836 53676 3892 53732
rect 3500 52834 3556 52836
rect 3500 52782 3502 52834
rect 3502 52782 3554 52834
rect 3554 52782 3556 52834
rect 3500 52780 3556 52782
rect 3612 51378 3668 51380
rect 3612 51326 3614 51378
rect 3614 51326 3666 51378
rect 3666 51326 3668 51378
rect 3612 51324 3668 51326
rect 4172 53730 4228 53732
rect 4172 53678 4174 53730
rect 4174 53678 4226 53730
rect 4226 53678 4228 53730
rect 4172 53676 4228 53678
rect 3836 51100 3892 51156
rect 3836 50652 3892 50708
rect 3388 50540 3444 50596
rect 3724 50540 3780 50596
rect 3388 50204 3444 50260
rect 3500 50370 3556 50372
rect 3500 50318 3502 50370
rect 3502 50318 3554 50370
rect 3554 50318 3556 50370
rect 3500 50316 3556 50318
rect 3500 49980 3556 50036
rect 3612 50092 3668 50148
rect 3276 49756 3332 49812
rect 2604 47458 2660 47460
rect 2604 47406 2606 47458
rect 2606 47406 2658 47458
rect 2658 47406 2660 47458
rect 2604 47404 2660 47406
rect 2044 45948 2100 46004
rect 2604 46396 2660 46452
rect 2156 45218 2212 45220
rect 2156 45166 2158 45218
rect 2158 45166 2210 45218
rect 2210 45166 2212 45218
rect 2156 45164 2212 45166
rect 1820 45052 1876 45108
rect 1596 40236 1652 40292
rect 1708 41580 1764 41636
rect 1484 38108 1540 38164
rect 1596 40012 1652 40068
rect 1596 37436 1652 37492
rect 1932 43932 1988 43988
rect 2156 44156 2212 44212
rect 1932 41804 1988 41860
rect 1820 38892 1876 38948
rect 2044 40124 2100 40180
rect 2156 39452 2212 39508
rect 2492 45388 2548 45444
rect 2492 45106 2548 45108
rect 2492 45054 2494 45106
rect 2494 45054 2546 45106
rect 2546 45054 2548 45106
rect 2492 45052 2548 45054
rect 2380 44994 2436 44996
rect 2380 44942 2382 44994
rect 2382 44942 2434 44994
rect 2434 44942 2436 44994
rect 2380 44940 2436 44942
rect 2828 47964 2884 48020
rect 2828 47628 2884 47684
rect 2940 46732 2996 46788
rect 2828 46674 2884 46676
rect 2828 46622 2830 46674
rect 2830 46622 2882 46674
rect 2882 46622 2884 46674
rect 2828 46620 2884 46622
rect 2828 45164 2884 45220
rect 2940 45052 2996 45108
rect 3276 48972 3332 49028
rect 3500 48076 3556 48132
rect 4956 53730 5012 53732
rect 4956 53678 4958 53730
rect 4958 53678 5010 53730
rect 5010 53678 5012 53730
rect 4956 53676 5012 53678
rect 5068 53340 5124 53396
rect 5404 56306 5460 56308
rect 5404 56254 5406 56306
rect 5406 56254 5458 56306
rect 5458 56254 5460 56306
rect 5404 56252 5460 56254
rect 5292 54012 5348 54068
rect 5404 53676 5460 53732
rect 5404 53452 5460 53508
rect 6748 59388 6804 59444
rect 6412 59330 6468 59332
rect 6412 59278 6414 59330
rect 6414 59278 6466 59330
rect 6466 59278 6468 59330
rect 6412 59276 6468 59278
rect 5852 59164 5908 59220
rect 7196 59164 7252 59220
rect 5964 59106 6020 59108
rect 5964 59054 5966 59106
rect 5966 59054 6018 59106
rect 6018 59054 6020 59106
rect 5964 59052 6020 59054
rect 8092 59388 8148 59444
rect 10668 59724 10724 59780
rect 8988 59612 9044 59668
rect 10108 59612 10164 59668
rect 9884 59500 9940 59556
rect 8652 59330 8708 59332
rect 8652 59278 8654 59330
rect 8654 59278 8706 59330
rect 8706 59278 8708 59330
rect 8652 59276 8708 59278
rect 5852 58940 5908 58996
rect 6300 58716 6356 58772
rect 5964 58210 6020 58212
rect 5964 58158 5966 58210
rect 5966 58158 6018 58210
rect 6018 58158 6020 58210
rect 5964 58156 6020 58158
rect 5852 56700 5908 56756
rect 5740 54402 5796 54404
rect 5740 54350 5742 54402
rect 5742 54350 5794 54402
rect 5794 54350 5796 54402
rect 5740 54348 5796 54350
rect 6748 58210 6804 58212
rect 6748 58158 6750 58210
rect 6750 58158 6802 58210
rect 6802 58158 6804 58210
rect 6748 58156 6804 58158
rect 6412 56642 6468 56644
rect 6412 56590 6414 56642
rect 6414 56590 6466 56642
rect 6466 56590 6468 56642
rect 6412 56588 6468 56590
rect 6188 54684 6244 54740
rect 6076 54572 6132 54628
rect 5628 53676 5684 53732
rect 6412 54572 6468 54628
rect 6300 54348 6356 54404
rect 6076 53506 6132 53508
rect 6076 53454 6078 53506
rect 6078 53454 6130 53506
rect 6130 53454 6132 53506
rect 6076 53452 6132 53454
rect 6188 53676 6244 53732
rect 5404 53058 5460 53060
rect 5404 53006 5406 53058
rect 5406 53006 5458 53058
rect 5458 53006 5460 53058
rect 5404 53004 5460 53006
rect 5516 52892 5572 52948
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 4284 52332 4340 52388
rect 4396 52220 4452 52276
rect 4172 51548 4228 51604
rect 4060 51100 4116 51156
rect 4060 50594 4116 50596
rect 4060 50542 4062 50594
rect 4062 50542 4114 50594
rect 4114 50542 4116 50594
rect 4060 50540 4116 50542
rect 3948 50428 4004 50484
rect 3948 49810 4004 49812
rect 3948 49758 3950 49810
rect 3950 49758 4002 49810
rect 4002 49758 4004 49810
rect 3948 49756 4004 49758
rect 5292 52220 5348 52276
rect 4844 52162 4900 52164
rect 4844 52110 4846 52162
rect 4846 52110 4898 52162
rect 4898 52110 4900 52162
rect 4844 52108 4900 52110
rect 4844 51602 4900 51604
rect 4844 51550 4846 51602
rect 4846 51550 4898 51602
rect 4898 51550 4900 51602
rect 4844 51548 4900 51550
rect 6860 57538 6916 57540
rect 6860 57486 6862 57538
rect 6862 57486 6914 57538
rect 6914 57486 6916 57538
rect 6860 57484 6916 57486
rect 7308 58322 7364 58324
rect 7308 58270 7310 58322
rect 7310 58270 7362 58322
rect 7362 58270 7364 58322
rect 7308 58268 7364 58270
rect 6860 56306 6916 56308
rect 6860 56254 6862 56306
rect 6862 56254 6914 56306
rect 6914 56254 6916 56306
rect 6860 56252 6916 56254
rect 6524 54012 6580 54068
rect 6636 55916 6692 55972
rect 6412 53900 6468 53956
rect 6524 53730 6580 53732
rect 6524 53678 6526 53730
rect 6526 53678 6578 53730
rect 6578 53678 6580 53730
rect 6524 53676 6580 53678
rect 6300 53170 6356 53172
rect 6300 53118 6302 53170
rect 6302 53118 6354 53170
rect 6354 53118 6356 53170
rect 6300 53116 6356 53118
rect 6076 52274 6132 52276
rect 6076 52222 6078 52274
rect 6078 52222 6130 52274
rect 6130 52222 6132 52274
rect 6076 52220 6132 52222
rect 5404 51548 5460 51604
rect 4396 51100 4452 51156
rect 5404 51212 5460 51268
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 4508 50706 4564 50708
rect 4508 50654 4510 50706
rect 4510 50654 4562 50706
rect 4562 50654 4564 50706
rect 4508 50652 4564 50654
rect 4844 50540 4900 50596
rect 4732 49922 4788 49924
rect 4732 49870 4734 49922
rect 4734 49870 4786 49922
rect 4786 49870 4788 49922
rect 4732 49868 4788 49870
rect 4956 50204 5012 50260
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 4172 48860 4228 48916
rect 5180 49644 5236 49700
rect 5068 49586 5124 49588
rect 5068 49534 5070 49586
rect 5070 49534 5122 49586
rect 5122 49534 5124 49586
rect 5068 49532 5124 49534
rect 4620 48802 4676 48804
rect 4620 48750 4622 48802
rect 4622 48750 4674 48802
rect 4674 48750 4676 48802
rect 4620 48748 4676 48750
rect 3724 47964 3780 48020
rect 3612 47346 3668 47348
rect 3612 47294 3614 47346
rect 3614 47294 3666 47346
rect 3666 47294 3668 47346
rect 3612 47292 3668 47294
rect 3948 46956 4004 47012
rect 3276 45612 3332 45668
rect 2716 44322 2772 44324
rect 2716 44270 2718 44322
rect 2718 44270 2770 44322
rect 2770 44270 2772 44322
rect 2716 44268 2772 44270
rect 3164 45276 3220 45332
rect 3500 46786 3556 46788
rect 3500 46734 3502 46786
rect 3502 46734 3554 46786
rect 3554 46734 3556 46786
rect 3500 46732 3556 46734
rect 3612 46172 3668 46228
rect 3612 45388 3668 45444
rect 3612 45164 3668 45220
rect 3388 44492 3444 44548
rect 3052 44268 3108 44324
rect 2492 43148 2548 43204
rect 2604 42866 2660 42868
rect 2604 42814 2606 42866
rect 2606 42814 2658 42866
rect 2658 42814 2660 42866
rect 2604 42812 2660 42814
rect 2492 42082 2548 42084
rect 2492 42030 2494 42082
rect 2494 42030 2546 42082
rect 2546 42030 2548 42082
rect 2492 42028 2548 42030
rect 2044 39394 2100 39396
rect 2044 39342 2046 39394
rect 2046 39342 2098 39394
rect 2098 39342 2100 39394
rect 2044 39340 2100 39342
rect 2380 40124 2436 40180
rect 2940 44044 2996 44100
rect 3724 44044 3780 44100
rect 3500 43932 3556 43988
rect 3388 43708 3444 43764
rect 3052 43596 3108 43652
rect 2940 42866 2996 42868
rect 2940 42814 2942 42866
rect 2942 42814 2994 42866
rect 2994 42814 2996 42866
rect 2940 42812 2996 42814
rect 2044 38834 2100 38836
rect 2044 38782 2046 38834
rect 2046 38782 2098 38834
rect 2098 38782 2100 38834
rect 2044 38780 2100 38782
rect 2380 39900 2436 39956
rect 1932 38668 1988 38724
rect 1708 36428 1764 36484
rect 1484 36316 1540 36372
rect 2268 38612 2324 38668
rect 2604 41074 2660 41076
rect 2604 41022 2606 41074
rect 2606 41022 2658 41074
rect 2658 41022 2660 41074
rect 2604 41020 2660 41022
rect 3164 41132 3220 41188
rect 3276 43148 3332 43204
rect 2828 40460 2884 40516
rect 2716 40348 2772 40404
rect 2604 40124 2660 40180
rect 3500 42364 3556 42420
rect 3724 42530 3780 42532
rect 3724 42478 3726 42530
rect 3726 42478 3778 42530
rect 3778 42478 3780 42530
rect 3724 42476 3780 42478
rect 4060 47852 4116 47908
rect 4172 47740 4228 47796
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 4844 47852 4900 47908
rect 4284 47516 4340 47572
rect 4172 46562 4228 46564
rect 4172 46510 4174 46562
rect 4174 46510 4226 46562
rect 4226 46510 4228 46562
rect 4172 46508 4228 46510
rect 5740 51602 5796 51604
rect 5740 51550 5742 51602
rect 5742 51550 5794 51602
rect 5794 51550 5796 51602
rect 5740 51548 5796 51550
rect 6748 54124 6804 54180
rect 6860 53564 6916 53620
rect 6300 51884 6356 51940
rect 6188 51100 6244 51156
rect 6188 50652 6244 50708
rect 6076 50540 6132 50596
rect 5852 50428 5908 50484
rect 5740 50370 5796 50372
rect 5740 50318 5742 50370
rect 5742 50318 5794 50370
rect 5794 50318 5796 50370
rect 5740 50316 5796 50318
rect 5628 50034 5684 50036
rect 5628 49982 5630 50034
rect 5630 49982 5682 50034
rect 5682 49982 5684 50034
rect 5628 49980 5684 49982
rect 5628 49308 5684 49364
rect 5516 49084 5572 49140
rect 4396 47068 4452 47124
rect 4620 46956 4676 47012
rect 4844 47012 4900 47068
rect 4844 46898 4900 46900
rect 4844 46846 4846 46898
rect 4846 46846 4898 46898
rect 4898 46846 4900 46898
rect 4844 46844 4900 46846
rect 4732 46786 4788 46788
rect 4732 46734 4734 46786
rect 4734 46734 4786 46786
rect 4786 46734 4788 46786
rect 4732 46732 4788 46734
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 4956 45836 5012 45892
rect 4508 45778 4564 45780
rect 4508 45726 4510 45778
rect 4510 45726 4562 45778
rect 4562 45726 4564 45778
rect 4508 45724 4564 45726
rect 4284 45276 4340 45332
rect 4396 45500 4452 45556
rect 4844 45276 4900 45332
rect 4508 44994 4564 44996
rect 4508 44942 4510 44994
rect 4510 44942 4562 44994
rect 4562 44942 4564 44994
rect 4508 44940 4564 44942
rect 4060 44828 4116 44884
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4396 44492 4452 44548
rect 4284 44380 4340 44436
rect 5068 44940 5124 44996
rect 4956 44210 5012 44212
rect 4956 44158 4958 44210
rect 4958 44158 5010 44210
rect 5010 44158 5012 44210
rect 4956 44156 5012 44158
rect 4844 43596 4900 43652
rect 5404 46844 5460 46900
rect 5292 43596 5348 43652
rect 5180 43484 5236 43540
rect 6748 53228 6804 53284
rect 7084 55468 7140 55524
rect 7644 59052 7700 59108
rect 7644 56700 7700 56756
rect 7420 56642 7476 56644
rect 7420 56590 7422 56642
rect 7422 56590 7474 56642
rect 7474 56590 7476 56642
rect 7420 56588 7476 56590
rect 7308 55970 7364 55972
rect 7308 55918 7310 55970
rect 7310 55918 7362 55970
rect 7362 55918 7364 55970
rect 7308 55916 7364 55918
rect 7196 55244 7252 55300
rect 7196 55074 7252 55076
rect 7196 55022 7198 55074
rect 7198 55022 7250 55074
rect 7250 55022 7252 55074
rect 7196 55020 7252 55022
rect 7420 54796 7476 54852
rect 7532 55132 7588 55188
rect 7308 54402 7364 54404
rect 7308 54350 7310 54402
rect 7310 54350 7362 54402
rect 7362 54350 7364 54402
rect 7308 54348 7364 54350
rect 7084 53676 7140 53732
rect 7532 53730 7588 53732
rect 7532 53678 7534 53730
rect 7534 53678 7586 53730
rect 7586 53678 7588 53730
rect 7532 53676 7588 53678
rect 7196 53564 7252 53620
rect 6972 53228 7028 53284
rect 5852 49532 5908 49588
rect 6300 49644 6356 49700
rect 6076 49084 6132 49140
rect 6076 48748 6132 48804
rect 5964 48636 6020 48692
rect 5964 48412 6020 48468
rect 5852 48188 5908 48244
rect 6188 47964 6244 48020
rect 5628 47516 5684 47572
rect 6076 47516 6132 47572
rect 5964 47292 6020 47348
rect 5628 46284 5684 46340
rect 4060 43314 4116 43316
rect 4060 43262 4062 43314
rect 4062 43262 4114 43314
rect 4114 43262 4116 43314
rect 4060 43260 4116 43262
rect 4060 42754 4116 42756
rect 4060 42702 4062 42754
rect 4062 42702 4114 42754
rect 4114 42702 4116 42754
rect 4060 42700 4116 42702
rect 3948 42364 4004 42420
rect 3724 42194 3780 42196
rect 3724 42142 3726 42194
rect 3726 42142 3778 42194
rect 3778 42142 3780 42194
rect 3724 42140 3780 42142
rect 3612 41410 3668 41412
rect 3612 41358 3614 41410
rect 3614 41358 3666 41410
rect 3666 41358 3668 41410
rect 3612 41356 3668 41358
rect 3836 41298 3892 41300
rect 3836 41246 3838 41298
rect 3838 41246 3890 41298
rect 3890 41246 3892 41298
rect 3836 41244 3892 41246
rect 3388 39900 3444 39956
rect 3500 40460 3556 40516
rect 3612 39788 3668 39844
rect 3388 39676 3444 39732
rect 2604 39228 2660 39284
rect 2492 38722 2548 38724
rect 2492 38670 2494 38722
rect 2494 38670 2546 38722
rect 2546 38670 2548 38722
rect 2492 38668 2548 38670
rect 2380 38162 2436 38164
rect 2380 38110 2382 38162
rect 2382 38110 2434 38162
rect 2434 38110 2436 38162
rect 2380 38108 2436 38110
rect 2604 38108 2660 38164
rect 3276 39340 3332 39396
rect 2940 38668 2996 38724
rect 3388 38722 3444 38724
rect 3388 38670 3390 38722
rect 3390 38670 3442 38722
rect 3442 38670 3444 38722
rect 3388 38668 3444 38670
rect 3612 39228 3668 39284
rect 4172 41970 4228 41972
rect 4172 41918 4174 41970
rect 4174 41918 4226 41970
rect 4226 41918 4228 41970
rect 4172 41916 4228 41918
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 4620 42028 4676 42084
rect 4956 41858 5012 41860
rect 4956 41806 4958 41858
rect 4958 41806 5010 41858
rect 5010 41806 5012 41858
rect 4956 41804 5012 41806
rect 4060 41132 4116 41188
rect 3836 39228 3892 39284
rect 3724 39116 3780 39172
rect 3836 39058 3892 39060
rect 3836 39006 3838 39058
rect 3838 39006 3890 39058
rect 3890 39006 3892 39058
rect 3836 39004 3892 39006
rect 3276 37826 3332 37828
rect 3276 37774 3278 37826
rect 3278 37774 3330 37826
rect 3330 37774 3332 37826
rect 3276 37772 3332 37774
rect 4060 39730 4116 39732
rect 4060 39678 4062 39730
rect 4062 39678 4114 39730
rect 4114 39678 4116 39730
rect 4060 39676 4116 39678
rect 3612 37660 3668 37716
rect 4060 39116 4116 39172
rect 3836 38444 3892 38500
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 5068 41580 5124 41636
rect 5180 42140 5236 42196
rect 4684 41524 4740 41526
rect 4844 41356 4900 41412
rect 4508 41186 4564 41188
rect 4508 41134 4510 41186
rect 4510 41134 4562 41186
rect 4562 41134 4564 41186
rect 4508 41132 4564 41134
rect 4732 40684 4788 40740
rect 4284 40626 4340 40628
rect 4284 40574 4286 40626
rect 4286 40574 4338 40626
rect 4338 40574 4340 40626
rect 4284 40572 4340 40574
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 4620 39506 4676 39508
rect 4620 39454 4622 39506
rect 4622 39454 4674 39506
rect 4674 39454 4676 39506
rect 4620 39452 4676 39454
rect 4172 38444 4228 38500
rect 4284 38892 4340 38948
rect 4060 38220 4116 38276
rect 4620 38946 4676 38948
rect 4620 38894 4622 38946
rect 4622 38894 4674 38946
rect 4674 38894 4676 38946
rect 4620 38892 4676 38894
rect 5068 40962 5124 40964
rect 5068 40910 5070 40962
rect 5070 40910 5122 40962
rect 5122 40910 5124 40962
rect 5068 40908 5124 40910
rect 4956 40460 5012 40516
rect 5068 40402 5124 40404
rect 5068 40350 5070 40402
rect 5070 40350 5122 40402
rect 5122 40350 5124 40402
rect 5068 40348 5124 40350
rect 5180 39676 5236 39732
rect 6076 46898 6132 46900
rect 6076 46846 6078 46898
rect 6078 46846 6130 46898
rect 6130 46846 6132 46898
rect 6076 46844 6132 46846
rect 6076 45500 6132 45556
rect 5740 43932 5796 43988
rect 5628 41916 5684 41972
rect 5740 42364 5796 42420
rect 5516 41858 5572 41860
rect 5516 41806 5518 41858
rect 5518 41806 5570 41858
rect 5570 41806 5572 41858
rect 5516 41804 5572 41806
rect 5964 45052 6020 45108
rect 6076 44716 6132 44772
rect 5964 44322 6020 44324
rect 5964 44270 5966 44322
rect 5966 44270 6018 44322
rect 6018 44270 6020 44322
rect 5964 44268 6020 44270
rect 6636 51772 6692 51828
rect 6860 52668 6916 52724
rect 6972 52332 7028 52388
rect 7196 52892 7252 52948
rect 6860 51548 6916 51604
rect 6748 51436 6804 51492
rect 7084 51436 7140 51492
rect 6860 51378 6916 51380
rect 6860 51326 6862 51378
rect 6862 51326 6914 51378
rect 6914 51326 6916 51378
rect 6860 51324 6916 51326
rect 6524 50204 6580 50260
rect 6972 50876 7028 50932
rect 6860 50706 6916 50708
rect 6860 50654 6862 50706
rect 6862 50654 6914 50706
rect 6914 50654 6916 50706
rect 6860 50652 6916 50654
rect 6748 50370 6804 50372
rect 6748 50318 6750 50370
rect 6750 50318 6802 50370
rect 6802 50318 6804 50370
rect 6748 50316 6804 50318
rect 6748 49532 6804 49588
rect 6748 48300 6804 48356
rect 6748 47516 6804 47572
rect 6860 49420 6916 49476
rect 6972 49084 7028 49140
rect 7308 52780 7364 52836
rect 7868 56476 7924 56532
rect 7756 52780 7812 52836
rect 8092 58716 8148 58772
rect 8652 57708 8708 57764
rect 8764 57820 8820 57876
rect 8204 57260 8260 57316
rect 8428 57484 8484 57540
rect 8092 56812 8148 56868
rect 8204 57036 8260 57092
rect 7980 55468 8036 55524
rect 8092 56588 8148 56644
rect 8092 56082 8148 56084
rect 8092 56030 8094 56082
rect 8094 56030 8146 56082
rect 8146 56030 8148 56082
rect 8092 56028 8148 56030
rect 8092 55244 8148 55300
rect 7868 55020 7924 55076
rect 7644 52668 7700 52724
rect 8092 55074 8148 55076
rect 8092 55022 8094 55074
rect 8094 55022 8146 55074
rect 8146 55022 8148 55074
rect 8092 55020 8148 55022
rect 8092 54796 8148 54852
rect 7980 53506 8036 53508
rect 7980 53454 7982 53506
rect 7982 53454 8034 53506
rect 8034 53454 8036 53506
rect 7980 53452 8036 53454
rect 8540 57426 8596 57428
rect 8540 57374 8542 57426
rect 8542 57374 8594 57426
rect 8594 57374 8596 57426
rect 8540 57372 8596 57374
rect 8764 56700 8820 56756
rect 8540 56364 8596 56420
rect 9772 59276 9828 59332
rect 9324 59052 9380 59108
rect 9100 58322 9156 58324
rect 9100 58270 9102 58322
rect 9102 58270 9154 58322
rect 9154 58270 9156 58322
rect 9100 58268 9156 58270
rect 8876 56364 8932 56420
rect 8988 58044 9044 58100
rect 8988 56252 9044 56308
rect 9212 56140 9268 56196
rect 8540 56028 8596 56084
rect 8764 55244 8820 55300
rect 8092 52834 8148 52836
rect 8092 52782 8094 52834
rect 8094 52782 8146 52834
rect 8146 52782 8148 52834
rect 8092 52780 8148 52782
rect 7644 51772 7700 51828
rect 7308 49698 7364 49700
rect 7308 49646 7310 49698
rect 7310 49646 7362 49698
rect 7362 49646 7364 49698
rect 7308 49644 7364 49646
rect 7308 49138 7364 49140
rect 7308 49086 7310 49138
rect 7310 49086 7362 49138
rect 7362 49086 7364 49138
rect 7308 49084 7364 49086
rect 6972 47740 7028 47796
rect 6860 47292 6916 47348
rect 7420 48636 7476 48692
rect 7756 51212 7812 51268
rect 7644 50876 7700 50932
rect 7868 50876 7924 50932
rect 7980 50652 8036 50708
rect 7868 50540 7924 50596
rect 7644 50482 7700 50484
rect 7644 50430 7646 50482
rect 7646 50430 7698 50482
rect 7698 50430 7700 50482
rect 7644 50428 7700 50430
rect 7980 50316 8036 50372
rect 7868 48802 7924 48804
rect 7868 48750 7870 48802
rect 7870 48750 7922 48802
rect 7922 48750 7924 48802
rect 7868 48748 7924 48750
rect 6636 46786 6692 46788
rect 6636 46734 6638 46786
rect 6638 46734 6690 46786
rect 6690 46734 6692 46786
rect 6636 46732 6692 46734
rect 6412 44940 6468 44996
rect 6412 43932 6468 43988
rect 6636 45890 6692 45892
rect 6636 45838 6638 45890
rect 6638 45838 6690 45890
rect 6690 45838 6692 45890
rect 6636 45836 6692 45838
rect 6972 46396 7028 46452
rect 7196 46674 7252 46676
rect 7196 46622 7198 46674
rect 7198 46622 7250 46674
rect 7250 46622 7252 46674
rect 7196 46620 7252 46622
rect 7868 47964 7924 48020
rect 7756 47516 7812 47572
rect 7644 47458 7700 47460
rect 7644 47406 7646 47458
rect 7646 47406 7698 47458
rect 7698 47406 7700 47458
rect 7644 47404 7700 47406
rect 7084 46060 7140 46116
rect 7532 46956 7588 47012
rect 6748 45724 6804 45780
rect 6636 45106 6692 45108
rect 6636 45054 6638 45106
rect 6638 45054 6690 45106
rect 6690 45054 6692 45106
rect 6636 45052 6692 45054
rect 6860 45666 6916 45668
rect 6860 45614 6862 45666
rect 6862 45614 6914 45666
rect 6914 45614 6916 45666
rect 6860 45612 6916 45614
rect 7084 45500 7140 45556
rect 7644 46786 7700 46788
rect 7644 46734 7646 46786
rect 7646 46734 7698 46786
rect 7698 46734 7700 46786
rect 7644 46732 7700 46734
rect 7308 45948 7364 46004
rect 8316 52780 8372 52836
rect 8204 51772 8260 51828
rect 8204 51324 8260 51380
rect 8540 52274 8596 52276
rect 8540 52222 8542 52274
rect 8542 52222 8594 52274
rect 8594 52222 8596 52274
rect 8540 52220 8596 52222
rect 9100 55132 9156 55188
rect 8988 55074 9044 55076
rect 8988 55022 8990 55074
rect 8990 55022 9042 55074
rect 9042 55022 9044 55074
rect 8988 55020 9044 55022
rect 8876 53676 8932 53732
rect 8988 53564 9044 53620
rect 9212 53730 9268 53732
rect 9212 53678 9214 53730
rect 9214 53678 9266 53730
rect 9266 53678 9268 53730
rect 9212 53676 9268 53678
rect 9100 53116 9156 53172
rect 9100 52162 9156 52164
rect 9100 52110 9102 52162
rect 9102 52110 9154 52162
rect 9154 52110 9156 52162
rect 9100 52108 9156 52110
rect 8652 51378 8708 51380
rect 8652 51326 8654 51378
rect 8654 51326 8706 51378
rect 8706 51326 8708 51378
rect 8652 51324 8708 51326
rect 8428 50316 8484 50372
rect 8652 50540 8708 50596
rect 8316 50034 8372 50036
rect 8316 49982 8318 50034
rect 8318 49982 8370 50034
rect 8370 49982 8372 50034
rect 8316 49980 8372 49982
rect 8876 51212 8932 51268
rect 9436 58268 9492 58324
rect 9436 57372 9492 57428
rect 14364 59836 14420 59892
rect 12348 59778 12404 59780
rect 12348 59726 12350 59778
rect 12350 59726 12402 59778
rect 12402 59726 12404 59778
rect 12348 59724 12404 59726
rect 12460 59612 12516 59668
rect 11564 59388 11620 59444
rect 10668 59330 10724 59332
rect 10668 59278 10670 59330
rect 10670 59278 10722 59330
rect 10722 59278 10724 59330
rect 10668 59276 10724 59278
rect 11004 59164 11060 59220
rect 9884 58322 9940 58324
rect 9884 58270 9886 58322
rect 9886 58270 9938 58322
rect 9938 58270 9940 58322
rect 9884 58268 9940 58270
rect 10780 59052 10836 59108
rect 9996 57650 10052 57652
rect 9996 57598 9998 57650
rect 9998 57598 10050 57650
rect 10050 57598 10052 57650
rect 9996 57596 10052 57598
rect 10444 57650 10500 57652
rect 10444 57598 10446 57650
rect 10446 57598 10498 57650
rect 10498 57598 10500 57650
rect 10444 57596 10500 57598
rect 10332 57260 10388 57316
rect 9772 55132 9828 55188
rect 9660 55020 9716 55076
rect 9772 54236 9828 54292
rect 9548 53788 9604 53844
rect 9660 54124 9716 54180
rect 9996 56194 10052 56196
rect 9996 56142 9998 56194
rect 9998 56142 10050 56194
rect 10050 56142 10052 56194
rect 9996 56140 10052 56142
rect 10108 55244 10164 55300
rect 9996 55186 10052 55188
rect 9996 55134 9998 55186
rect 9998 55134 10050 55186
rect 10050 55134 10052 55186
rect 9996 55132 10052 55134
rect 10220 55020 10276 55076
rect 10108 54908 10164 54964
rect 10780 58044 10836 58100
rect 10556 57148 10612 57204
rect 10780 56140 10836 56196
rect 10668 55356 10724 55412
rect 11340 57708 11396 57764
rect 11116 56866 11172 56868
rect 11116 56814 11118 56866
rect 11118 56814 11170 56866
rect 11170 56814 11172 56866
rect 11116 56812 11172 56814
rect 11788 58716 11844 58772
rect 11564 57372 11620 57428
rect 11676 58210 11732 58212
rect 11676 58158 11678 58210
rect 11678 58158 11730 58210
rect 11730 58158 11732 58210
rect 11676 58156 11732 58158
rect 11676 57260 11732 57316
rect 11564 56642 11620 56644
rect 11564 56590 11566 56642
rect 11566 56590 11618 56642
rect 11618 56590 11620 56642
rect 11564 56588 11620 56590
rect 11228 56476 11284 56532
rect 11116 56306 11172 56308
rect 11116 56254 11118 56306
rect 11118 56254 11170 56306
rect 11170 56254 11172 56306
rect 11116 56252 11172 56254
rect 11340 56082 11396 56084
rect 11340 56030 11342 56082
rect 11342 56030 11394 56082
rect 11394 56030 11396 56082
rect 11340 56028 11396 56030
rect 12348 59106 12404 59108
rect 12348 59054 12350 59106
rect 12350 59054 12402 59106
rect 12402 59054 12404 59106
rect 12348 59052 12404 59054
rect 12124 58940 12180 58996
rect 12348 57148 12404 57204
rect 12012 57036 12068 57092
rect 11900 56140 11956 56196
rect 11788 55916 11844 55972
rect 12124 56082 12180 56084
rect 12124 56030 12126 56082
rect 12126 56030 12178 56082
rect 12178 56030 12180 56082
rect 12124 56028 12180 56030
rect 11004 55356 11060 55412
rect 11452 55804 11508 55860
rect 10444 55244 10500 55300
rect 11228 55132 11284 55188
rect 10332 54684 10388 54740
rect 10108 54572 10164 54628
rect 9884 53170 9940 53172
rect 9884 53118 9886 53170
rect 9886 53118 9938 53170
rect 9938 53118 9940 53170
rect 9884 53116 9940 53118
rect 9436 52668 9492 52724
rect 10220 54402 10276 54404
rect 10220 54350 10222 54402
rect 10222 54350 10274 54402
rect 10274 54350 10276 54402
rect 10220 54348 10276 54350
rect 10556 54236 10612 54292
rect 10444 54012 10500 54068
rect 10108 53116 10164 53172
rect 10332 53676 10388 53732
rect 9996 52220 10052 52276
rect 9324 51212 9380 51268
rect 8988 50652 9044 50708
rect 9772 51100 9828 51156
rect 9100 50594 9156 50596
rect 9100 50542 9102 50594
rect 9102 50542 9154 50594
rect 9154 50542 9156 50594
rect 9100 50540 9156 50542
rect 8316 49644 8372 49700
rect 8092 46956 8148 47012
rect 8540 49084 8596 49140
rect 7868 46620 7924 46676
rect 6524 43708 6580 43764
rect 6076 42754 6132 42756
rect 6076 42702 6078 42754
rect 6078 42702 6130 42754
rect 6130 42702 6132 42754
rect 6076 42700 6132 42702
rect 5964 41692 6020 41748
rect 5852 41356 5908 41412
rect 5852 40236 5908 40292
rect 6076 41074 6132 41076
rect 6076 41022 6078 41074
rect 6078 41022 6130 41074
rect 6130 41022 6132 41074
rect 6076 41020 6132 41022
rect 5740 39900 5796 39956
rect 4956 39564 5012 39620
rect 4844 38946 4900 38948
rect 4844 38894 4846 38946
rect 4846 38894 4898 38946
rect 4898 38894 4900 38946
rect 4844 38892 4900 38894
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4620 38220 4676 38276
rect 4060 38050 4116 38052
rect 4060 37998 4062 38050
rect 4062 37998 4114 38050
rect 4114 37998 4116 38050
rect 4060 37996 4116 37998
rect 2268 37100 2324 37156
rect 2268 36258 2324 36260
rect 2268 36206 2270 36258
rect 2270 36206 2322 36258
rect 2322 36206 2324 36258
rect 2268 36204 2324 36206
rect 2044 35756 2100 35812
rect 1820 35084 1876 35140
rect 1484 32844 1540 32900
rect 1596 34748 1652 34804
rect 1484 30716 1540 30772
rect 2044 34412 2100 34468
rect 1932 34018 1988 34020
rect 1932 33966 1934 34018
rect 1934 33966 1986 34018
rect 1986 33966 1988 34018
rect 1932 33964 1988 33966
rect 2380 35196 2436 35252
rect 2492 36988 2548 37044
rect 2380 34636 2436 34692
rect 2156 33964 2212 34020
rect 2268 34188 2324 34244
rect 1932 32844 1988 32900
rect 2492 32732 2548 32788
rect 3052 37154 3108 37156
rect 3052 37102 3054 37154
rect 3054 37102 3106 37154
rect 3106 37102 3108 37154
rect 3052 37100 3108 37102
rect 2940 36540 2996 36596
rect 2828 36482 2884 36484
rect 2828 36430 2830 36482
rect 2830 36430 2882 36482
rect 2882 36430 2884 36482
rect 2828 36428 2884 36430
rect 2828 34690 2884 34692
rect 2828 34638 2830 34690
rect 2830 34638 2882 34690
rect 2882 34638 2884 34690
rect 2828 34636 2884 34638
rect 3276 36428 3332 36484
rect 3276 35868 3332 35924
rect 2828 33122 2884 33124
rect 2828 33070 2830 33122
rect 2830 33070 2882 33122
rect 2882 33070 2884 33122
rect 2828 33068 2884 33070
rect 3388 36092 3444 36148
rect 3836 37378 3892 37380
rect 3836 37326 3838 37378
rect 3838 37326 3890 37378
rect 3890 37326 3892 37378
rect 3836 37324 3892 37326
rect 4284 37938 4340 37940
rect 4284 37886 4286 37938
rect 4286 37886 4338 37938
rect 4338 37886 4340 37938
rect 4284 37884 4340 37886
rect 4172 37772 4228 37828
rect 3948 37212 4004 37268
rect 4060 37660 4116 37716
rect 3724 36988 3780 37044
rect 3948 36370 4004 36372
rect 3948 36318 3950 36370
rect 3950 36318 4002 36370
rect 4002 36318 4004 36370
rect 3948 36316 4004 36318
rect 3836 36092 3892 36148
rect 3724 35474 3780 35476
rect 3724 35422 3726 35474
rect 3726 35422 3778 35474
rect 3778 35422 3780 35474
rect 3724 35420 3780 35422
rect 3500 35196 3556 35252
rect 3388 34914 3444 34916
rect 3388 34862 3390 34914
rect 3390 34862 3442 34914
rect 3442 34862 3444 34914
rect 3388 34860 3444 34862
rect 4508 37660 4564 37716
rect 5180 39340 5236 39396
rect 5516 39116 5572 39172
rect 5068 38332 5124 38388
rect 5628 38722 5684 38724
rect 5628 38670 5630 38722
rect 5630 38670 5682 38722
rect 5682 38670 5684 38722
rect 5628 38668 5684 38670
rect 5068 38162 5124 38164
rect 5068 38110 5070 38162
rect 5070 38110 5122 38162
rect 5122 38110 5124 38162
rect 5068 38108 5124 38110
rect 4620 37100 4676 37156
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4732 35698 4788 35700
rect 4732 35646 4734 35698
rect 4734 35646 4786 35698
rect 4786 35646 4788 35698
rect 4732 35644 4788 35646
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 3388 33516 3444 33572
rect 3724 34076 3780 34132
rect 3500 33292 3556 33348
rect 3612 33628 3668 33684
rect 2940 32450 2996 32452
rect 2940 32398 2942 32450
rect 2942 32398 2994 32450
rect 2994 32398 2996 32450
rect 2940 32396 2996 32398
rect 3388 32284 3444 32340
rect 2268 31836 2324 31892
rect 2044 31500 2100 31556
rect 1708 26460 1764 26516
rect 1596 23996 1652 24052
rect 1932 29820 1988 29876
rect 2380 31948 2436 32004
rect 3836 33628 3892 33684
rect 4396 35026 4452 35028
rect 4396 34974 4398 35026
rect 4398 34974 4450 35026
rect 4450 34974 4452 35026
rect 4396 34972 4452 34974
rect 5068 37884 5124 37940
rect 5404 37100 5460 37156
rect 4956 35308 5012 35364
rect 5068 36204 5124 36260
rect 4844 34748 4900 34804
rect 4284 34412 4340 34468
rect 4508 34636 4564 34692
rect 4172 34354 4228 34356
rect 4172 34302 4174 34354
rect 4174 34302 4226 34354
rect 4226 34302 4228 34354
rect 4172 34300 4228 34302
rect 3948 33404 4004 33460
rect 4172 33964 4228 34020
rect 4284 33852 4340 33908
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4060 33516 4116 33572
rect 3500 31948 3556 32004
rect 3836 32508 3892 32564
rect 2828 31666 2884 31668
rect 2828 31614 2830 31666
rect 2830 31614 2882 31666
rect 2882 31614 2884 31666
rect 2828 31612 2884 31614
rect 3388 31276 3444 31332
rect 2380 29820 2436 29876
rect 3388 30380 3444 30436
rect 2716 30156 2772 30212
rect 2044 27916 2100 27972
rect 1932 27746 1988 27748
rect 1932 27694 1934 27746
rect 1934 27694 1986 27746
rect 1986 27694 1988 27746
rect 1932 27692 1988 27694
rect 1932 26850 1988 26852
rect 1932 26798 1934 26850
rect 1934 26798 1986 26850
rect 1986 26798 1988 26850
rect 1932 26796 1988 26798
rect 1932 26514 1988 26516
rect 1932 26462 1934 26514
rect 1934 26462 1986 26514
rect 1986 26462 1988 26514
rect 1932 26460 1988 26462
rect 1820 25564 1876 25620
rect 3276 30210 3332 30212
rect 3276 30158 3278 30210
rect 3278 30158 3330 30210
rect 3330 30158 3332 30210
rect 3276 30156 3332 30158
rect 3500 29650 3556 29652
rect 3500 29598 3502 29650
rect 3502 29598 3554 29650
rect 3554 29598 3556 29650
rect 3500 29596 3556 29598
rect 2492 26908 2548 26964
rect 2604 27132 2660 27188
rect 2380 26796 2436 26852
rect 2268 26460 2324 26516
rect 2492 26124 2548 26180
rect 2268 25452 2324 25508
rect 2380 25282 2436 25284
rect 2380 25230 2382 25282
rect 2382 25230 2434 25282
rect 2434 25230 2436 25282
rect 2380 25228 2436 25230
rect 1484 23436 1540 23492
rect 1820 21980 1876 22036
rect 3052 27074 3108 27076
rect 3052 27022 3054 27074
rect 3054 27022 3106 27074
rect 3106 27022 3108 27074
rect 3052 27020 3108 27022
rect 3500 27692 3556 27748
rect 2940 26514 2996 26516
rect 2940 26462 2942 26514
rect 2942 26462 2994 26514
rect 2994 26462 2996 26514
rect 2940 26460 2996 26462
rect 3388 26236 3444 26292
rect 3500 27132 3556 27188
rect 2828 26124 2884 26180
rect 2716 25116 2772 25172
rect 2268 23212 2324 23268
rect 2156 22482 2212 22484
rect 2156 22430 2158 22482
rect 2158 22430 2210 22482
rect 2210 22430 2212 22482
rect 2156 22428 2212 22430
rect 3276 26178 3332 26180
rect 3276 26126 3278 26178
rect 3278 26126 3330 26178
rect 3330 26126 3332 26178
rect 3276 26124 3332 26126
rect 2940 25788 2996 25844
rect 3164 25228 3220 25284
rect 3500 25788 3556 25844
rect 2828 22428 2884 22484
rect 2716 21868 2772 21924
rect 1820 21698 1876 21700
rect 1820 21646 1822 21698
rect 1822 21646 1874 21698
rect 1874 21646 1876 21698
rect 1820 21644 1876 21646
rect 2156 21532 2212 21588
rect 2268 21756 2324 21812
rect 1932 20300 1988 20356
rect 3052 21756 3108 21812
rect 3724 31836 3780 31892
rect 3836 30828 3892 30884
rect 3724 28812 3780 28868
rect 3948 29036 4004 29092
rect 3836 27692 3892 27748
rect 4284 33234 4340 33236
rect 4284 33182 4286 33234
rect 4286 33182 4338 33234
rect 4338 33182 4340 33234
rect 4284 33180 4340 33182
rect 5740 38332 5796 38388
rect 5628 37154 5684 37156
rect 5628 37102 5630 37154
rect 5630 37102 5682 37154
rect 5682 37102 5684 37154
rect 5628 37100 5684 37102
rect 5516 36988 5572 37044
rect 5740 36764 5796 36820
rect 6300 43426 6356 43428
rect 6300 43374 6302 43426
rect 6302 43374 6354 43426
rect 6354 43374 6356 43426
rect 6300 43372 6356 43374
rect 7532 45948 7588 46004
rect 7532 45276 7588 45332
rect 7980 45890 8036 45892
rect 7980 45838 7982 45890
rect 7982 45838 8034 45890
rect 8034 45838 8036 45890
rect 7980 45836 8036 45838
rect 8204 46508 8260 46564
rect 8316 48860 8372 48916
rect 8204 45778 8260 45780
rect 8204 45726 8206 45778
rect 8206 45726 8258 45778
rect 8258 45726 8260 45778
rect 8204 45724 8260 45726
rect 8092 45612 8148 45668
rect 7084 44604 7140 44660
rect 7196 44044 7252 44100
rect 7084 43596 7140 43652
rect 6748 43538 6804 43540
rect 6748 43486 6750 43538
rect 6750 43486 6802 43538
rect 6802 43486 6804 43538
rect 6748 43484 6804 43486
rect 6412 42812 6468 42868
rect 6860 42812 6916 42868
rect 6636 42476 6692 42532
rect 6524 42252 6580 42308
rect 6300 42140 6356 42196
rect 6636 41916 6692 41972
rect 6524 41804 6580 41860
rect 7868 43820 7924 43876
rect 7868 43596 7924 43652
rect 7420 43484 7476 43540
rect 7420 41970 7476 41972
rect 7420 41918 7422 41970
rect 7422 41918 7474 41970
rect 7474 41918 7476 41970
rect 7420 41916 7476 41918
rect 6748 40796 6804 40852
rect 6412 40626 6468 40628
rect 6412 40574 6414 40626
rect 6414 40574 6466 40626
rect 6466 40574 6468 40626
rect 6412 40572 6468 40574
rect 6972 40626 7028 40628
rect 6972 40574 6974 40626
rect 6974 40574 7026 40626
rect 7026 40574 7028 40626
rect 6972 40572 7028 40574
rect 7420 41132 7476 41188
rect 7644 43538 7700 43540
rect 7644 43486 7646 43538
rect 7646 43486 7698 43538
rect 7698 43486 7700 43538
rect 7644 43484 7700 43486
rect 7756 42812 7812 42868
rect 7532 40908 7588 40964
rect 7196 40572 7252 40628
rect 7756 40796 7812 40852
rect 7868 40460 7924 40516
rect 10332 52556 10388 52612
rect 9772 50482 9828 50484
rect 9772 50430 9774 50482
rect 9774 50430 9826 50482
rect 9826 50430 9828 50482
rect 9772 50428 9828 50430
rect 8988 50316 9044 50372
rect 10220 50652 10276 50708
rect 11116 54012 11172 54068
rect 10892 52556 10948 52612
rect 11228 52556 11284 52612
rect 11340 52220 11396 52276
rect 10444 52050 10500 52052
rect 10444 51998 10446 52050
rect 10446 51998 10498 52050
rect 10498 51998 10500 52050
rect 10444 51996 10500 51998
rect 10444 51212 10500 51268
rect 10556 50316 10612 50372
rect 9996 49868 10052 49924
rect 8876 48802 8932 48804
rect 8876 48750 8878 48802
rect 8878 48750 8930 48802
rect 8930 48750 8932 48802
rect 8876 48748 8932 48750
rect 8428 48636 8484 48692
rect 8428 48242 8484 48244
rect 8428 48190 8430 48242
rect 8430 48190 8482 48242
rect 8482 48190 8484 48242
rect 8428 48188 8484 48190
rect 8428 44380 8484 44436
rect 8652 48188 8708 48244
rect 9548 49756 9604 49812
rect 9212 49420 9268 49476
rect 8988 48412 9044 48468
rect 8764 47852 8820 47908
rect 8764 46956 8820 47012
rect 9436 47516 9492 47572
rect 9212 47346 9268 47348
rect 9212 47294 9214 47346
rect 9214 47294 9266 47346
rect 9266 47294 9268 47346
rect 9212 47292 9268 47294
rect 10108 49308 10164 49364
rect 11116 51884 11172 51940
rect 11788 54460 11844 54516
rect 12796 59500 12852 59556
rect 13468 59612 13524 59668
rect 12908 58828 12964 58884
rect 13020 59164 13076 59220
rect 12684 58380 12740 58436
rect 13244 59106 13300 59108
rect 13244 59054 13246 59106
rect 13246 59054 13298 59106
rect 13298 59054 13300 59106
rect 13244 59052 13300 59054
rect 13468 58940 13524 58996
rect 12124 55410 12180 55412
rect 12124 55358 12126 55410
rect 12126 55358 12178 55410
rect 12178 55358 12180 55410
rect 12124 55356 12180 55358
rect 12012 55244 12068 55300
rect 12124 55132 12180 55188
rect 11900 53116 11956 53172
rect 11676 52332 11732 52388
rect 11564 51772 11620 51828
rect 10892 50594 10948 50596
rect 10892 50542 10894 50594
rect 10894 50542 10946 50594
rect 10946 50542 10948 50594
rect 10892 50540 10948 50542
rect 10668 49980 10724 50036
rect 11116 51378 11172 51380
rect 11116 51326 11118 51378
rect 11118 51326 11170 51378
rect 11170 51326 11172 51378
rect 11116 51324 11172 51326
rect 11564 51154 11620 51156
rect 11564 51102 11566 51154
rect 11566 51102 11618 51154
rect 11618 51102 11620 51154
rect 11564 51100 11620 51102
rect 11676 50652 11732 50708
rect 10892 49980 10948 50036
rect 9884 48748 9940 48804
rect 9996 48412 10052 48468
rect 9772 47964 9828 48020
rect 10332 49026 10388 49028
rect 10332 48974 10334 49026
rect 10334 48974 10386 49026
rect 10386 48974 10388 49026
rect 10332 48972 10388 48974
rect 10668 48972 10724 49028
rect 10220 48636 10276 48692
rect 10220 48412 10276 48468
rect 10332 48748 10388 48804
rect 10220 48242 10276 48244
rect 10220 48190 10222 48242
rect 10222 48190 10274 48242
rect 10274 48190 10276 48242
rect 10220 48188 10276 48190
rect 9100 46620 9156 46676
rect 8652 45948 8708 46004
rect 8764 46508 8820 46564
rect 8876 46396 8932 46452
rect 8652 44380 8708 44436
rect 8540 44098 8596 44100
rect 8540 44046 8542 44098
rect 8542 44046 8594 44098
rect 8594 44046 8596 44098
rect 8540 44044 8596 44046
rect 8540 43820 8596 43876
rect 8876 45948 8932 46004
rect 9100 45890 9156 45892
rect 9100 45838 9102 45890
rect 9102 45838 9154 45890
rect 9154 45838 9156 45890
rect 9100 45836 9156 45838
rect 9772 46562 9828 46564
rect 9772 46510 9774 46562
rect 9774 46510 9826 46562
rect 9826 46510 9828 46562
rect 9772 46508 9828 46510
rect 9772 46172 9828 46228
rect 9660 44994 9716 44996
rect 9660 44942 9662 44994
rect 9662 44942 9714 44994
rect 9714 44942 9716 44994
rect 9660 44940 9716 44942
rect 9212 44828 9268 44884
rect 9436 44156 9492 44212
rect 8764 43596 8820 43652
rect 8876 43820 8932 43876
rect 8092 43036 8148 43092
rect 8428 42812 8484 42868
rect 8540 42754 8596 42756
rect 8540 42702 8542 42754
rect 8542 42702 8594 42754
rect 8594 42702 8596 42754
rect 8540 42700 8596 42702
rect 8428 42252 8484 42308
rect 8204 42028 8260 42084
rect 7980 40572 8036 40628
rect 6300 39564 6356 39620
rect 6188 39340 6244 39396
rect 6076 38834 6132 38836
rect 6076 38782 6078 38834
rect 6078 38782 6130 38834
rect 6130 38782 6132 38834
rect 6076 38780 6132 38782
rect 5964 37212 6020 37268
rect 6076 37154 6132 37156
rect 6076 37102 6078 37154
rect 6078 37102 6130 37154
rect 6130 37102 6132 37154
rect 6076 37100 6132 37102
rect 6300 38892 6356 38948
rect 6636 39564 6692 39620
rect 7084 39788 7140 39844
rect 6300 38722 6356 38724
rect 6300 38670 6302 38722
rect 6302 38670 6354 38722
rect 6354 38670 6356 38722
rect 6300 38668 6356 38670
rect 6860 39116 6916 39172
rect 6748 38332 6804 38388
rect 6636 37884 6692 37940
rect 6748 38050 6804 38052
rect 6748 37998 6750 38050
rect 6750 37998 6802 38050
rect 6802 37998 6804 38050
rect 6748 37996 6804 37998
rect 7084 38668 7140 38724
rect 7308 40178 7364 40180
rect 7308 40126 7310 40178
rect 7310 40126 7362 40178
rect 7362 40126 7364 40178
rect 7308 40124 7364 40126
rect 7308 38946 7364 38948
rect 7308 38894 7310 38946
rect 7310 38894 7362 38946
rect 7362 38894 7364 38946
rect 7308 38892 7364 38894
rect 7084 37996 7140 38052
rect 6748 37436 6804 37492
rect 6860 37212 6916 37268
rect 5852 36092 5908 36148
rect 5740 35698 5796 35700
rect 5740 35646 5742 35698
rect 5742 35646 5794 35698
rect 5794 35646 5796 35698
rect 5740 35644 5796 35646
rect 5516 35532 5572 35588
rect 5404 34972 5460 35028
rect 5516 35308 5572 35364
rect 5516 34860 5572 34916
rect 5292 34524 5348 34580
rect 5516 34524 5572 34580
rect 5404 34412 5460 34468
rect 5180 34188 5236 34244
rect 5292 33852 5348 33908
rect 5068 33628 5124 33684
rect 4844 33180 4900 33236
rect 5180 33292 5236 33348
rect 4284 32508 4340 32564
rect 4508 32562 4564 32564
rect 4508 32510 4510 32562
rect 4510 32510 4562 32562
rect 4562 32510 4564 32562
rect 4508 32508 4564 32510
rect 4172 31276 4228 31332
rect 4284 32284 4340 32340
rect 4172 30940 4228 30996
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4844 32172 4900 32228
rect 4684 32116 4740 32118
rect 5068 31890 5124 31892
rect 5068 31838 5070 31890
rect 5070 31838 5122 31890
rect 5122 31838 5124 31890
rect 5068 31836 5124 31838
rect 5180 30994 5236 30996
rect 5180 30942 5182 30994
rect 5182 30942 5234 30994
rect 5234 30942 5236 30994
rect 5180 30940 5236 30942
rect 5292 33068 5348 33124
rect 4844 30828 4900 30884
rect 4620 30716 4676 30772
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 5068 30268 5124 30324
rect 6188 36652 6244 36708
rect 5964 35308 6020 35364
rect 6076 34748 6132 34804
rect 5964 34690 6020 34692
rect 5964 34638 5966 34690
rect 5966 34638 6018 34690
rect 6018 34638 6020 34690
rect 5964 34636 6020 34638
rect 5964 34242 6020 34244
rect 5964 34190 5966 34242
rect 5966 34190 6018 34242
rect 6018 34190 6020 34242
rect 5964 34188 6020 34190
rect 6524 36764 6580 36820
rect 6636 37100 6692 37156
rect 6412 36204 6468 36260
rect 6300 34860 6356 34916
rect 5628 33346 5684 33348
rect 5628 33294 5630 33346
rect 5630 33294 5682 33346
rect 5682 33294 5684 33346
rect 5628 33292 5684 33294
rect 5516 32786 5572 32788
rect 5516 32734 5518 32786
rect 5518 32734 5570 32786
rect 5570 32734 5572 32786
rect 5516 32732 5572 32734
rect 5516 32172 5572 32228
rect 4620 29820 4676 29876
rect 4284 29650 4340 29652
rect 4284 29598 4286 29650
rect 4286 29598 4338 29650
rect 4338 29598 4340 29650
rect 4284 29596 4340 29598
rect 4620 29484 4676 29540
rect 4172 28812 4228 28868
rect 4172 27580 4228 27636
rect 4172 27186 4228 27188
rect 4172 27134 4174 27186
rect 4174 27134 4226 27186
rect 4226 27134 4228 27186
rect 4172 27132 4228 27134
rect 3612 25228 3668 25284
rect 3724 24946 3780 24948
rect 3724 24894 3726 24946
rect 3726 24894 3778 24946
rect 3778 24894 3780 24946
rect 3724 24892 3780 24894
rect 4060 26572 4116 26628
rect 4844 29484 4900 29540
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4508 28754 4564 28756
rect 4508 28702 4510 28754
rect 4510 28702 4562 28754
rect 4562 28702 4564 28754
rect 4508 28700 4564 28702
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4284 26572 4340 26628
rect 4732 26908 4788 26964
rect 4172 26460 4228 26516
rect 4284 26236 4340 26292
rect 4060 25788 4116 25844
rect 5404 30940 5460 30996
rect 5404 30268 5460 30324
rect 5628 30380 5684 30436
rect 5516 29596 5572 29652
rect 5180 28700 5236 28756
rect 4956 27132 5012 27188
rect 4956 26962 5012 26964
rect 4956 26910 4958 26962
rect 4958 26910 5010 26962
rect 5010 26910 5012 26962
rect 4956 26908 5012 26910
rect 4844 26684 4900 26740
rect 5068 26796 5124 26852
rect 4844 26402 4900 26404
rect 4844 26350 4846 26402
rect 4846 26350 4898 26402
rect 4898 26350 4900 26402
rect 4844 26348 4900 26350
rect 4956 26124 5012 26180
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4060 25394 4116 25396
rect 4060 25342 4062 25394
rect 4062 25342 4114 25394
rect 4114 25342 4116 25394
rect 4060 25340 4116 25342
rect 3500 24108 3556 24164
rect 3724 24050 3780 24052
rect 3724 23998 3726 24050
rect 3726 23998 3778 24050
rect 3778 23998 3780 24050
rect 3724 23996 3780 23998
rect 3612 23548 3668 23604
rect 3052 21586 3108 21588
rect 3052 21534 3054 21586
rect 3054 21534 3106 21586
rect 3106 21534 3108 21586
rect 3052 21532 3108 21534
rect 2716 20914 2772 20916
rect 2716 20862 2718 20914
rect 2718 20862 2770 20914
rect 2770 20862 2772 20914
rect 2716 20860 2772 20862
rect 3164 21420 3220 21476
rect 3948 24668 4004 24724
rect 4060 22482 4116 22484
rect 4060 22430 4062 22482
rect 4062 22430 4114 22482
rect 4114 22430 4116 22482
rect 4060 22428 4116 22430
rect 3724 21420 3780 21476
rect 3948 21644 4004 21700
rect 2380 20076 2436 20132
rect 1820 19906 1876 19908
rect 1820 19854 1822 19906
rect 1822 19854 1874 19906
rect 1874 19854 1876 19906
rect 1820 19852 1876 19854
rect 1148 19740 1204 19796
rect 3052 20018 3108 20020
rect 3052 19966 3054 20018
rect 3054 19966 3106 20018
rect 3106 19966 3108 20018
rect 3052 19964 3108 19966
rect 3500 20018 3556 20020
rect 3500 19966 3502 20018
rect 3502 19966 3554 20018
rect 3554 19966 3556 20018
rect 3500 19964 3556 19966
rect 3612 19852 3668 19908
rect 4060 22204 4116 22260
rect 3948 21474 4004 21476
rect 3948 21422 3950 21474
rect 3950 21422 4002 21474
rect 4002 21422 4004 21474
rect 3948 21420 4004 21422
rect 4172 22092 4228 22148
rect 4060 20914 4116 20916
rect 4060 20862 4062 20914
rect 4062 20862 4114 20914
rect 4114 20862 4116 20914
rect 4060 20860 4116 20862
rect 3612 19180 3668 19236
rect 3724 18562 3780 18564
rect 3724 18510 3726 18562
rect 3726 18510 3778 18562
rect 3778 18510 3780 18562
rect 3724 18508 3780 18510
rect 4172 19404 4228 19460
rect 4956 25340 5012 25396
rect 4844 25282 4900 25284
rect 4844 25230 4846 25282
rect 4846 25230 4898 25282
rect 4898 25230 4900 25282
rect 4844 25228 4900 25230
rect 4732 24722 4788 24724
rect 4732 24670 4734 24722
rect 4734 24670 4786 24722
rect 4786 24670 4788 24722
rect 4732 24668 4788 24670
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4956 23826 5012 23828
rect 4956 23774 4958 23826
rect 4958 23774 5010 23826
rect 5010 23774 5012 23826
rect 4956 23772 5012 23774
rect 4620 23266 4676 23268
rect 4620 23214 4622 23266
rect 4622 23214 4674 23266
rect 4674 23214 4676 23266
rect 4620 23212 4676 23214
rect 5068 23266 5124 23268
rect 5068 23214 5070 23266
rect 5070 23214 5122 23266
rect 5122 23214 5124 23266
rect 5068 23212 5124 23214
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4844 22370 4900 22372
rect 4844 22318 4846 22370
rect 4846 22318 4898 22370
rect 4898 22318 4900 22370
rect 4844 22316 4900 22318
rect 5068 22204 5124 22260
rect 4844 21586 4900 21588
rect 4844 21534 4846 21586
rect 4846 21534 4898 21586
rect 4898 21534 4900 21586
rect 4844 21532 4900 21534
rect 4396 21474 4452 21476
rect 4396 21422 4398 21474
rect 4398 21422 4450 21474
rect 4450 21422 4452 21474
rect 4396 21420 4452 21422
rect 5852 29148 5908 29204
rect 5404 28476 5460 28532
rect 5740 28476 5796 28532
rect 5292 27244 5348 27300
rect 5292 26908 5348 26964
rect 6636 35084 6692 35140
rect 6412 34130 6468 34132
rect 6412 34078 6414 34130
rect 6414 34078 6466 34130
rect 6466 34078 6468 34130
rect 6412 34076 6468 34078
rect 6524 34188 6580 34244
rect 6412 33852 6468 33908
rect 6076 33516 6132 33572
rect 6076 33068 6132 33124
rect 6188 32674 6244 32676
rect 6188 32622 6190 32674
rect 6190 32622 6242 32674
rect 6242 32622 6244 32674
rect 6188 32620 6244 32622
rect 6076 31948 6132 32004
rect 6412 33180 6468 33236
rect 7084 36988 7140 37044
rect 7196 36876 7252 36932
rect 7644 39900 7700 39956
rect 7756 39788 7812 39844
rect 7644 39340 7700 39396
rect 7868 39618 7924 39620
rect 7868 39566 7870 39618
rect 7870 39566 7922 39618
rect 7922 39566 7924 39618
rect 7868 39564 7924 39566
rect 7756 39004 7812 39060
rect 7420 38444 7476 38500
rect 7644 38834 7700 38836
rect 7644 38782 7646 38834
rect 7646 38782 7698 38834
rect 7698 38782 7700 38834
rect 7644 38780 7700 38782
rect 7756 38556 7812 38612
rect 7532 37938 7588 37940
rect 7532 37886 7534 37938
rect 7534 37886 7586 37938
rect 7586 37886 7588 37938
rect 7532 37884 7588 37886
rect 7980 39004 8036 39060
rect 8092 40908 8148 40964
rect 8316 40572 8372 40628
rect 8988 43426 9044 43428
rect 8988 43374 8990 43426
rect 8990 43374 9042 43426
rect 9042 43374 9044 43426
rect 8988 43372 9044 43374
rect 9100 43148 9156 43204
rect 8764 43036 8820 43092
rect 8988 42754 9044 42756
rect 8988 42702 8990 42754
rect 8990 42702 9042 42754
rect 9042 42702 9044 42754
rect 8988 42700 9044 42702
rect 8652 41020 8708 41076
rect 8764 42252 8820 42308
rect 8316 39116 8372 39172
rect 8316 38892 8372 38948
rect 7980 38722 8036 38724
rect 7980 38670 7982 38722
rect 7982 38670 8034 38722
rect 8034 38670 8036 38722
rect 7980 38668 8036 38670
rect 8428 38780 8484 38836
rect 8092 38220 8148 38276
rect 8204 38444 8260 38500
rect 7756 36988 7812 37044
rect 7980 37154 8036 37156
rect 7980 37102 7982 37154
rect 7982 37102 8034 37154
rect 8034 37102 8036 37154
rect 7980 37100 8036 37102
rect 7308 36540 7364 36596
rect 7868 36594 7924 36596
rect 7868 36542 7870 36594
rect 7870 36542 7922 36594
rect 7922 36542 7924 36594
rect 7868 36540 7924 36542
rect 7308 35868 7364 35924
rect 7420 36316 7476 36372
rect 6860 34188 6916 34244
rect 6972 35196 7028 35252
rect 7196 35084 7252 35140
rect 7308 34914 7364 34916
rect 7308 34862 7310 34914
rect 7310 34862 7362 34914
rect 7362 34862 7364 34914
rect 7308 34860 7364 34862
rect 6748 34076 6804 34132
rect 7196 34690 7252 34692
rect 7196 34638 7198 34690
rect 7198 34638 7250 34690
rect 7250 34638 7252 34690
rect 7196 34636 7252 34638
rect 7644 36092 7700 36148
rect 7644 35586 7700 35588
rect 7644 35534 7646 35586
rect 7646 35534 7698 35586
rect 7698 35534 7700 35586
rect 7644 35532 7700 35534
rect 6972 33404 7028 33460
rect 6188 31724 6244 31780
rect 6300 31500 6356 31556
rect 6188 31388 6244 31444
rect 6076 29650 6132 29652
rect 6076 29598 6078 29650
rect 6078 29598 6130 29650
rect 6130 29598 6132 29650
rect 6076 29596 6132 29598
rect 6300 31276 6356 31332
rect 7084 34188 7140 34244
rect 6972 32732 7028 32788
rect 6972 32172 7028 32228
rect 7532 33292 7588 33348
rect 8652 40348 8708 40404
rect 8876 42028 8932 42084
rect 8876 41858 8932 41860
rect 8876 41806 8878 41858
rect 8878 41806 8930 41858
rect 8930 41806 8932 41858
rect 8876 41804 8932 41806
rect 9212 42754 9268 42756
rect 9212 42702 9214 42754
rect 9214 42702 9266 42754
rect 9266 42702 9268 42754
rect 9212 42700 9268 42702
rect 9324 42252 9380 42308
rect 9212 41074 9268 41076
rect 9212 41022 9214 41074
rect 9214 41022 9266 41074
rect 9266 41022 9268 41074
rect 9212 41020 9268 41022
rect 9660 44044 9716 44100
rect 10220 47628 10276 47684
rect 10444 48412 10500 48468
rect 10556 47628 10612 47684
rect 10556 47292 10612 47348
rect 10556 46786 10612 46788
rect 10556 46734 10558 46786
rect 10558 46734 10610 46786
rect 10610 46734 10612 46786
rect 10556 46732 10612 46734
rect 10892 49586 10948 49588
rect 10892 49534 10894 49586
rect 10894 49534 10946 49586
rect 10946 49534 10948 49586
rect 10892 49532 10948 49534
rect 11004 48972 11060 49028
rect 11116 49084 11172 49140
rect 11004 48802 11060 48804
rect 11004 48750 11006 48802
rect 11006 48750 11058 48802
rect 11058 48750 11060 48802
rect 11004 48748 11060 48750
rect 11004 48412 11060 48468
rect 10892 48076 10948 48132
rect 11452 50034 11508 50036
rect 11452 49982 11454 50034
rect 11454 49982 11506 50034
rect 11506 49982 11508 50034
rect 11452 49980 11508 49982
rect 11676 50034 11732 50036
rect 11676 49982 11678 50034
rect 11678 49982 11730 50034
rect 11730 49982 11732 50034
rect 11676 49980 11732 49982
rect 11452 49756 11508 49812
rect 11788 49420 11844 49476
rect 11452 49308 11508 49364
rect 11676 49196 11732 49252
rect 11340 48242 11396 48244
rect 11340 48190 11342 48242
rect 11342 48190 11394 48242
rect 11394 48190 11396 48242
rect 11340 48188 11396 48190
rect 11452 47628 11508 47684
rect 11116 47180 11172 47236
rect 11004 47068 11060 47124
rect 10108 44604 10164 44660
rect 10444 45052 10500 45108
rect 10332 44940 10388 44996
rect 10220 44380 10276 44436
rect 10332 44322 10388 44324
rect 10332 44270 10334 44322
rect 10334 44270 10386 44322
rect 10386 44270 10388 44322
rect 10332 44268 10388 44270
rect 10220 44156 10276 44212
rect 9772 43650 9828 43652
rect 9772 43598 9774 43650
rect 9774 43598 9826 43650
rect 9826 43598 9828 43650
rect 9772 43596 9828 43598
rect 10444 44210 10500 44212
rect 10444 44158 10446 44210
rect 10446 44158 10498 44210
rect 10498 44158 10500 44210
rect 10444 44156 10500 44158
rect 10332 43708 10388 43764
rect 10444 43650 10500 43652
rect 10444 43598 10446 43650
rect 10446 43598 10498 43650
rect 10498 43598 10500 43650
rect 10444 43596 10500 43598
rect 10220 43314 10276 43316
rect 10220 43262 10222 43314
rect 10222 43262 10274 43314
rect 10274 43262 10276 43314
rect 10220 43260 10276 43262
rect 9660 42812 9716 42868
rect 9884 42642 9940 42644
rect 9884 42590 9886 42642
rect 9886 42590 9938 42642
rect 9938 42590 9940 42642
rect 9884 42588 9940 42590
rect 10332 42476 10388 42532
rect 10780 46284 10836 46340
rect 11004 46844 11060 46900
rect 11564 46956 11620 47012
rect 11340 46732 11396 46788
rect 10780 45330 10836 45332
rect 10780 45278 10782 45330
rect 10782 45278 10834 45330
rect 10834 45278 10836 45330
rect 10780 45276 10836 45278
rect 10780 45106 10836 45108
rect 10780 45054 10782 45106
rect 10782 45054 10834 45106
rect 10834 45054 10836 45106
rect 10780 45052 10836 45054
rect 10668 42700 10724 42756
rect 10668 42364 10724 42420
rect 10108 41468 10164 41524
rect 9548 41244 9604 41300
rect 9436 41020 9492 41076
rect 8652 38332 8708 38388
rect 8988 39058 9044 39060
rect 8988 39006 8990 39058
rect 8990 39006 9042 39058
rect 9042 39006 9044 39058
rect 8988 39004 9044 39006
rect 8764 38108 8820 38164
rect 9212 38668 9268 38724
rect 9772 40908 9828 40964
rect 7756 33292 7812 33348
rect 7980 34802 8036 34804
rect 7980 34750 7982 34802
rect 7982 34750 8034 34802
rect 8034 34750 8036 34802
rect 7980 34748 8036 34750
rect 8428 36540 8484 36596
rect 8764 37212 8820 37268
rect 8652 36876 8708 36932
rect 8652 36652 8708 36708
rect 8540 36092 8596 36148
rect 8540 35922 8596 35924
rect 8540 35870 8542 35922
rect 8542 35870 8594 35922
rect 8594 35870 8596 35922
rect 8540 35868 8596 35870
rect 8092 34690 8148 34692
rect 8092 34638 8094 34690
rect 8094 34638 8146 34690
rect 8146 34638 8148 34690
rect 8092 34636 8148 34638
rect 7868 33180 7924 33236
rect 7868 32844 7924 32900
rect 7644 32620 7700 32676
rect 7196 31948 7252 32004
rect 6636 31276 6692 31332
rect 6636 30492 6692 30548
rect 6412 28754 6468 28756
rect 6412 28702 6414 28754
rect 6414 28702 6466 28754
rect 6466 28702 6468 28754
rect 6412 28700 6468 28702
rect 6524 27916 6580 27972
rect 6300 27132 6356 27188
rect 6748 30828 6804 30884
rect 7084 30994 7140 30996
rect 7084 30942 7086 30994
rect 7086 30942 7138 30994
rect 7138 30942 7140 30994
rect 7084 30940 7140 30942
rect 7756 31778 7812 31780
rect 7756 31726 7758 31778
rect 7758 31726 7810 31778
rect 7810 31726 7812 31778
rect 7756 31724 7812 31726
rect 7644 31554 7700 31556
rect 7644 31502 7646 31554
rect 7646 31502 7698 31554
rect 7698 31502 7700 31554
rect 7644 31500 7700 31502
rect 7308 30882 7364 30884
rect 7308 30830 7310 30882
rect 7310 30830 7362 30882
rect 7362 30830 7364 30882
rect 7308 30828 7364 30830
rect 6860 29484 6916 29540
rect 7196 30210 7252 30212
rect 7196 30158 7198 30210
rect 7198 30158 7250 30210
rect 7250 30158 7252 30210
rect 7196 30156 7252 30158
rect 8092 34188 8148 34244
rect 8764 34972 8820 35028
rect 7980 33852 8036 33908
rect 8540 34412 8596 34468
rect 8428 33740 8484 33796
rect 8092 33458 8148 33460
rect 8092 33406 8094 33458
rect 8094 33406 8146 33458
rect 8146 33406 8148 33458
rect 8092 33404 8148 33406
rect 8540 32844 8596 32900
rect 8428 32732 8484 32788
rect 8092 32450 8148 32452
rect 8092 32398 8094 32450
rect 8094 32398 8146 32450
rect 8146 32398 8148 32450
rect 8092 32396 8148 32398
rect 7980 31612 8036 31668
rect 8092 31276 8148 31332
rect 7980 30210 8036 30212
rect 7980 30158 7982 30210
rect 7982 30158 8034 30210
rect 8034 30158 8036 30210
rect 7980 30156 8036 30158
rect 7084 28530 7140 28532
rect 7084 28478 7086 28530
rect 7086 28478 7138 28530
rect 7138 28478 7140 28530
rect 7084 28476 7140 28478
rect 6972 27580 7028 27636
rect 7532 27916 7588 27972
rect 6748 27074 6804 27076
rect 6748 27022 6750 27074
rect 6750 27022 6802 27074
rect 6802 27022 6804 27074
rect 6748 27020 6804 27022
rect 7084 27020 7140 27076
rect 6524 26908 6580 26964
rect 5292 26684 5348 26740
rect 5404 26290 5460 26292
rect 5404 26238 5406 26290
rect 5406 26238 5458 26290
rect 5458 26238 5460 26290
rect 5404 26236 5460 26238
rect 5964 26124 6020 26180
rect 5740 25116 5796 25172
rect 5740 23996 5796 24052
rect 5628 23378 5684 23380
rect 5628 23326 5630 23378
rect 5630 23326 5682 23378
rect 5682 23326 5684 23378
rect 5628 23324 5684 23326
rect 5292 22204 5348 22260
rect 5516 23212 5572 23268
rect 5740 22428 5796 22484
rect 6300 25676 6356 25732
rect 6748 26012 6804 26068
rect 6972 24722 7028 24724
rect 6972 24670 6974 24722
rect 6974 24670 7026 24722
rect 7026 24670 7028 24722
rect 6972 24668 7028 24670
rect 7308 26124 7364 26180
rect 7868 28924 7924 28980
rect 7980 28476 8036 28532
rect 8092 28252 8148 28308
rect 8092 27804 8148 27860
rect 7980 27468 8036 27524
rect 8652 31666 8708 31668
rect 8652 31614 8654 31666
rect 8654 31614 8706 31666
rect 8706 31614 8708 31666
rect 8652 31612 8708 31614
rect 8540 31164 8596 31220
rect 8428 30940 8484 30996
rect 9324 38556 9380 38612
rect 9436 40124 9492 40180
rect 8988 38274 9044 38276
rect 8988 38222 8990 38274
rect 8990 38222 9042 38274
rect 9042 38222 9044 38274
rect 8988 38220 9044 38222
rect 9100 38050 9156 38052
rect 9100 37998 9102 38050
rect 9102 37998 9154 38050
rect 9154 37998 9156 38050
rect 9100 37996 9156 37998
rect 9212 37884 9268 37940
rect 9212 37660 9268 37716
rect 9772 40124 9828 40180
rect 9884 39618 9940 39620
rect 9884 39566 9886 39618
rect 9886 39566 9938 39618
rect 9938 39566 9940 39618
rect 9884 39564 9940 39566
rect 10108 39676 10164 39732
rect 10220 39564 10276 39620
rect 10668 41186 10724 41188
rect 10668 41134 10670 41186
rect 10670 41134 10722 41186
rect 10722 41134 10724 41186
rect 10668 41132 10724 41134
rect 10556 40402 10612 40404
rect 10556 40350 10558 40402
rect 10558 40350 10610 40402
rect 10610 40350 10612 40402
rect 10556 40348 10612 40350
rect 10556 40178 10612 40180
rect 10556 40126 10558 40178
rect 10558 40126 10610 40178
rect 10610 40126 10612 40178
rect 10556 40124 10612 40126
rect 10444 40012 10500 40068
rect 11452 46284 11508 46340
rect 11788 48466 11844 48468
rect 11788 48414 11790 48466
rect 11790 48414 11842 48466
rect 11842 48414 11844 48466
rect 11788 48412 11844 48414
rect 11788 46732 11844 46788
rect 11452 45724 11508 45780
rect 11452 45052 11508 45108
rect 11676 46172 11732 46228
rect 11676 45164 11732 45220
rect 11564 44268 11620 44324
rect 11116 44156 11172 44212
rect 11564 43708 11620 43764
rect 11452 43650 11508 43652
rect 11452 43598 11454 43650
rect 11454 43598 11506 43650
rect 11506 43598 11508 43650
rect 11452 43596 11508 43598
rect 11228 42812 11284 42868
rect 12796 58210 12852 58212
rect 12796 58158 12798 58210
rect 12798 58158 12850 58210
rect 12850 58158 12852 58210
rect 12796 58156 12852 58158
rect 12796 57538 12852 57540
rect 12796 57486 12798 57538
rect 12798 57486 12850 57538
rect 12850 57486 12852 57538
rect 12796 57484 12852 57486
rect 13132 57372 13188 57428
rect 13020 56476 13076 56532
rect 12908 56252 12964 56308
rect 12796 56194 12852 56196
rect 12796 56142 12798 56194
rect 12798 56142 12850 56194
rect 12850 56142 12852 56194
rect 12796 56140 12852 56142
rect 12684 55580 12740 55636
rect 12236 54236 12292 54292
rect 13916 59052 13972 59108
rect 13804 58434 13860 58436
rect 13804 58382 13806 58434
rect 13806 58382 13858 58434
rect 13858 58382 13860 58434
rect 13804 58380 13860 58382
rect 13692 57484 13748 57540
rect 13692 57260 13748 57316
rect 13580 57036 13636 57092
rect 13468 56476 13524 56532
rect 13244 56364 13300 56420
rect 12348 52892 12404 52948
rect 12460 54012 12516 54068
rect 12236 52556 12292 52612
rect 12572 53730 12628 53732
rect 12572 53678 12574 53730
rect 12574 53678 12626 53730
rect 12626 53678 12628 53730
rect 12572 53676 12628 53678
rect 13356 55356 13412 55412
rect 13356 54460 13412 54516
rect 13244 53900 13300 53956
rect 14364 59218 14420 59220
rect 14364 59166 14366 59218
rect 14366 59166 14418 59218
rect 14418 59166 14420 59218
rect 14364 59164 14420 59166
rect 14700 59890 14756 59892
rect 14700 59838 14702 59890
rect 14702 59838 14754 59890
rect 14754 59838 14756 59890
rect 14700 59836 14756 59838
rect 14924 59778 14980 59780
rect 14924 59726 14926 59778
rect 14926 59726 14978 59778
rect 14978 59726 14980 59778
rect 14924 59724 14980 59726
rect 15708 59612 15764 59668
rect 15932 59724 15988 59780
rect 14028 58828 14084 58884
rect 14028 58156 14084 58212
rect 16044 59106 16100 59108
rect 16044 59054 16046 59106
rect 16046 59054 16098 59106
rect 16098 59054 16100 59106
rect 16044 59052 16100 59054
rect 15932 58828 15988 58884
rect 14700 58322 14756 58324
rect 14700 58270 14702 58322
rect 14702 58270 14754 58322
rect 14754 58270 14756 58322
rect 14700 58268 14756 58270
rect 15484 58322 15540 58324
rect 15484 58270 15486 58322
rect 15486 58270 15538 58322
rect 15538 58270 15540 58322
rect 15484 58268 15540 58270
rect 14924 57820 14980 57876
rect 14140 56866 14196 56868
rect 14140 56814 14142 56866
rect 14142 56814 14194 56866
rect 14194 56814 14196 56866
rect 14140 56812 14196 56814
rect 14028 55970 14084 55972
rect 14028 55918 14030 55970
rect 14030 55918 14082 55970
rect 14082 55918 14084 55970
rect 14028 55916 14084 55918
rect 14924 57538 14980 57540
rect 14924 57486 14926 57538
rect 14926 57486 14978 57538
rect 14978 57486 14980 57538
rect 14924 57484 14980 57486
rect 15260 57708 15316 57764
rect 14812 56924 14868 56980
rect 14364 56812 14420 56868
rect 14588 56642 14644 56644
rect 14588 56590 14590 56642
rect 14590 56590 14642 56642
rect 14642 56590 14644 56642
rect 14588 56588 14644 56590
rect 14252 56140 14308 56196
rect 13804 55132 13860 55188
rect 13692 53676 13748 53732
rect 12908 53340 12964 53396
rect 12684 53170 12740 53172
rect 12684 53118 12686 53170
rect 12686 53118 12738 53170
rect 12738 53118 12740 53170
rect 12684 53116 12740 53118
rect 12460 52162 12516 52164
rect 12460 52110 12462 52162
rect 12462 52110 12514 52162
rect 12514 52110 12516 52162
rect 12460 52108 12516 52110
rect 12460 51884 12516 51940
rect 12348 51772 12404 51828
rect 12236 50706 12292 50708
rect 12236 50654 12238 50706
rect 12238 50654 12290 50706
rect 12290 50654 12292 50706
rect 12236 50652 12292 50654
rect 13132 52834 13188 52836
rect 13132 52782 13134 52834
rect 13134 52782 13186 52834
rect 13186 52782 13188 52834
rect 13132 52780 13188 52782
rect 13468 52780 13524 52836
rect 13132 52444 13188 52500
rect 13020 52162 13076 52164
rect 13020 52110 13022 52162
rect 13022 52110 13074 52162
rect 13074 52110 13076 52162
rect 13020 52108 13076 52110
rect 12572 50988 12628 51044
rect 12684 50540 12740 50596
rect 12460 49922 12516 49924
rect 12460 49870 12462 49922
rect 12462 49870 12514 49922
rect 12514 49870 12516 49922
rect 12460 49868 12516 49870
rect 12348 49810 12404 49812
rect 12348 49758 12350 49810
rect 12350 49758 12402 49810
rect 12402 49758 12404 49810
rect 12348 49756 12404 49758
rect 12124 48748 12180 48804
rect 12348 49138 12404 49140
rect 12348 49086 12350 49138
rect 12350 49086 12402 49138
rect 12402 49086 12404 49138
rect 12348 49084 12404 49086
rect 12236 48636 12292 48692
rect 12012 48076 12068 48132
rect 12796 49532 12852 49588
rect 12572 48972 12628 49028
rect 12684 48802 12740 48804
rect 12684 48750 12686 48802
rect 12686 48750 12738 48802
rect 12738 48750 12740 48802
rect 12684 48748 12740 48750
rect 12572 48188 12628 48244
rect 12236 46956 12292 47012
rect 12124 46002 12180 46004
rect 12124 45950 12126 46002
rect 12126 45950 12178 46002
rect 12178 45950 12180 46002
rect 12124 45948 12180 45950
rect 12348 44828 12404 44884
rect 12012 44322 12068 44324
rect 12012 44270 12014 44322
rect 12014 44270 12066 44322
rect 12066 44270 12068 44322
rect 12012 44268 12068 44270
rect 12236 44268 12292 44324
rect 11788 43820 11844 43876
rect 12348 43932 12404 43988
rect 12908 48242 12964 48244
rect 12908 48190 12910 48242
rect 12910 48190 12962 48242
rect 12962 48190 12964 48242
rect 12908 48188 12964 48190
rect 13244 49698 13300 49700
rect 13244 49646 13246 49698
rect 13246 49646 13298 49698
rect 13298 49646 13300 49698
rect 13244 49644 13300 49646
rect 13132 49532 13188 49588
rect 13356 48972 13412 49028
rect 12684 46172 12740 46228
rect 12684 46002 12740 46004
rect 12684 45950 12686 46002
rect 12686 45950 12738 46002
rect 12738 45950 12740 46002
rect 12684 45948 12740 45950
rect 12796 45836 12852 45892
rect 12684 45276 12740 45332
rect 12572 44828 12628 44884
rect 12796 45218 12852 45220
rect 12796 45166 12798 45218
rect 12798 45166 12850 45218
rect 12850 45166 12852 45218
rect 12796 45164 12852 45166
rect 12684 44044 12740 44100
rect 13356 48076 13412 48132
rect 14140 54684 14196 54740
rect 14028 54626 14084 54628
rect 14028 54574 14030 54626
rect 14030 54574 14082 54626
rect 14082 54574 14084 54626
rect 14028 54572 14084 54574
rect 14252 54572 14308 54628
rect 14028 54124 14084 54180
rect 14028 53954 14084 53956
rect 14028 53902 14030 53954
rect 14030 53902 14082 53954
rect 14082 53902 14084 53954
rect 14028 53900 14084 53902
rect 13804 53228 13860 53284
rect 13804 52556 13860 52612
rect 14364 52834 14420 52836
rect 14364 52782 14366 52834
rect 14366 52782 14418 52834
rect 14418 52782 14420 52834
rect 14364 52780 14420 52782
rect 14588 54908 14644 54964
rect 14588 54236 14644 54292
rect 14700 53676 14756 53732
rect 15372 57538 15428 57540
rect 15372 57486 15374 57538
rect 15374 57486 15426 57538
rect 15426 57486 15428 57538
rect 15372 57484 15428 57486
rect 17612 59500 17668 59556
rect 18060 59500 18116 59556
rect 18508 59500 18564 59556
rect 17948 59442 18004 59444
rect 17948 59390 17950 59442
rect 17950 59390 18002 59442
rect 18002 59390 18004 59442
rect 17948 59388 18004 59390
rect 18396 59276 18452 59332
rect 16604 58940 16660 58996
rect 15484 56924 15540 56980
rect 16492 58828 16548 58884
rect 16044 56866 16100 56868
rect 16044 56814 16046 56866
rect 16046 56814 16098 56866
rect 16098 56814 16100 56866
rect 16044 56812 16100 56814
rect 15932 56252 15988 56308
rect 15148 55410 15204 55412
rect 15148 55358 15150 55410
rect 15150 55358 15202 55410
rect 15202 55358 15204 55410
rect 15148 55356 15204 55358
rect 15820 55132 15876 55188
rect 15708 55074 15764 55076
rect 15708 55022 15710 55074
rect 15710 55022 15762 55074
rect 15762 55022 15764 55074
rect 15708 55020 15764 55022
rect 15596 54012 15652 54068
rect 15036 53900 15092 53956
rect 15820 53954 15876 53956
rect 15820 53902 15822 53954
rect 15822 53902 15874 53954
rect 15874 53902 15876 53954
rect 15820 53900 15876 53902
rect 16940 58716 16996 58772
rect 16604 58546 16660 58548
rect 16604 58494 16606 58546
rect 16606 58494 16658 58546
rect 16658 58494 16660 58546
rect 16604 58492 16660 58494
rect 16268 58434 16324 58436
rect 16268 58382 16270 58434
rect 16270 58382 16322 58434
rect 16322 58382 16324 58434
rect 16268 58380 16324 58382
rect 16492 57036 16548 57092
rect 16492 56700 16548 56756
rect 16828 56700 16884 56756
rect 14588 53116 14644 53172
rect 14924 53452 14980 53508
rect 13804 52274 13860 52276
rect 13804 52222 13806 52274
rect 13806 52222 13858 52274
rect 13858 52222 13860 52274
rect 13804 52220 13860 52222
rect 14252 52332 14308 52388
rect 13692 51436 13748 51492
rect 14028 51996 14084 52052
rect 14812 52946 14868 52948
rect 14812 52894 14814 52946
rect 14814 52894 14866 52946
rect 14866 52894 14868 52946
rect 14812 52892 14868 52894
rect 15372 53506 15428 53508
rect 15372 53454 15374 53506
rect 15374 53454 15426 53506
rect 15426 53454 15428 53506
rect 15372 53452 15428 53454
rect 14924 52668 14980 52724
rect 14476 51884 14532 51940
rect 14812 52050 14868 52052
rect 14812 51998 14814 52050
rect 14814 51998 14866 52050
rect 14866 51998 14868 52050
rect 14812 51996 14868 51998
rect 14028 50594 14084 50596
rect 14028 50542 14030 50594
rect 14030 50542 14082 50594
rect 14082 50542 14084 50594
rect 14028 50540 14084 50542
rect 13804 50482 13860 50484
rect 13804 50430 13806 50482
rect 13806 50430 13858 50482
rect 13858 50430 13860 50482
rect 14140 51436 14196 51492
rect 14252 51378 14308 51380
rect 14252 51326 14254 51378
rect 14254 51326 14306 51378
rect 14306 51326 14308 51378
rect 14252 51324 14308 51326
rect 15260 52780 15316 52836
rect 15148 52162 15204 52164
rect 15148 52110 15150 52162
rect 15150 52110 15202 52162
rect 15202 52110 15204 52162
rect 15148 52108 15204 52110
rect 14140 50764 14196 50820
rect 14700 50652 14756 50708
rect 13804 50428 13860 50430
rect 13804 49810 13860 49812
rect 13804 49758 13806 49810
rect 13806 49758 13858 49810
rect 13858 49758 13860 49810
rect 13804 49756 13860 49758
rect 13468 45724 13524 45780
rect 13244 45612 13300 45668
rect 13132 44156 13188 44212
rect 13020 43820 13076 43876
rect 14700 50204 14756 50260
rect 14476 49868 14532 49924
rect 14364 49138 14420 49140
rect 14364 49086 14366 49138
rect 14366 49086 14418 49138
rect 14418 49086 14420 49138
rect 14364 49084 14420 49086
rect 14588 48972 14644 49028
rect 14140 48636 14196 48692
rect 14588 48748 14644 48804
rect 14140 48242 14196 48244
rect 14140 48190 14142 48242
rect 14142 48190 14194 48242
rect 14194 48190 14196 48242
rect 14140 48188 14196 48190
rect 14364 48242 14420 48244
rect 14364 48190 14366 48242
rect 14366 48190 14418 48242
rect 14418 48190 14420 48242
rect 14364 48188 14420 48190
rect 14812 50092 14868 50148
rect 14812 49698 14868 49700
rect 14812 49646 14814 49698
rect 14814 49646 14866 49698
rect 14866 49646 14868 49698
rect 14812 49644 14868 49646
rect 14924 49196 14980 49252
rect 14924 48860 14980 48916
rect 15372 52444 15428 52500
rect 16380 54124 16436 54180
rect 16156 53228 16212 53284
rect 16716 55186 16772 55188
rect 16716 55134 16718 55186
rect 16718 55134 16770 55186
rect 16770 55134 16772 55186
rect 16716 55132 16772 55134
rect 18172 58604 18228 58660
rect 17500 58434 17556 58436
rect 17500 58382 17502 58434
rect 17502 58382 17554 58434
rect 17554 58382 17556 58434
rect 17500 58380 17556 58382
rect 18060 58434 18116 58436
rect 18060 58382 18062 58434
rect 18062 58382 18114 58434
rect 18114 58382 18116 58434
rect 18060 58380 18116 58382
rect 17052 57484 17108 57540
rect 17612 57538 17668 57540
rect 17612 57486 17614 57538
rect 17614 57486 17666 57538
rect 17666 57486 17668 57538
rect 17612 57484 17668 57486
rect 17500 56866 17556 56868
rect 17500 56814 17502 56866
rect 17502 56814 17554 56866
rect 17554 56814 17556 56866
rect 17500 56812 17556 56814
rect 17276 56754 17332 56756
rect 17276 56702 17278 56754
rect 17278 56702 17330 56754
rect 17330 56702 17332 56754
rect 17276 56700 17332 56702
rect 16940 54124 16996 54180
rect 16604 53954 16660 53956
rect 16604 53902 16606 53954
rect 16606 53902 16658 53954
rect 16658 53902 16660 53954
rect 16604 53900 16660 53902
rect 18172 57538 18228 57540
rect 18172 57486 18174 57538
rect 18174 57486 18226 57538
rect 18226 57486 18228 57538
rect 18172 57484 18228 57486
rect 17724 57090 17780 57092
rect 17724 57038 17726 57090
rect 17726 57038 17778 57090
rect 17778 57038 17780 57090
rect 17724 57036 17780 57038
rect 18396 56812 18452 56868
rect 18060 56700 18116 56756
rect 17836 56252 17892 56308
rect 18620 59106 18676 59108
rect 18620 59054 18622 59106
rect 18622 59054 18674 59106
rect 18674 59054 18676 59106
rect 18620 59052 18676 59054
rect 18956 58268 19012 58324
rect 18620 57036 18676 57092
rect 19180 58268 19236 58324
rect 19292 57596 19348 57652
rect 19516 59330 19572 59332
rect 19516 59278 19518 59330
rect 19518 59278 19570 59330
rect 19570 59278 19572 59330
rect 19516 59276 19572 59278
rect 19404 57260 19460 57316
rect 19836 59610 19892 59612
rect 19836 59558 19838 59610
rect 19838 59558 19890 59610
rect 19890 59558 19892 59610
rect 19836 59556 19892 59558
rect 19940 59610 19996 59612
rect 19940 59558 19942 59610
rect 19942 59558 19994 59610
rect 19994 59558 19996 59610
rect 19940 59556 19996 59558
rect 20044 59610 20100 59612
rect 20044 59558 20046 59610
rect 20046 59558 20098 59610
rect 20098 59558 20100 59610
rect 20044 59556 20100 59558
rect 20076 59330 20132 59332
rect 20076 59278 20078 59330
rect 20078 59278 20130 59330
rect 20130 59278 20132 59330
rect 20076 59276 20132 59278
rect 20076 59052 20132 59108
rect 19852 58322 19908 58324
rect 19852 58270 19854 58322
rect 19854 58270 19906 58322
rect 19906 58270 19908 58322
rect 19852 58268 19908 58270
rect 20300 58492 20356 58548
rect 20188 58380 20244 58436
rect 19836 58042 19892 58044
rect 19836 57990 19838 58042
rect 19838 57990 19890 58042
rect 19890 57990 19892 58042
rect 19836 57988 19892 57990
rect 19940 58042 19996 58044
rect 19940 57990 19942 58042
rect 19942 57990 19994 58042
rect 19994 57990 19996 58042
rect 19940 57988 19996 57990
rect 20044 58042 20100 58044
rect 20044 57990 20046 58042
rect 20046 57990 20098 58042
rect 20098 57990 20100 58042
rect 20044 57988 20100 57990
rect 19852 57650 19908 57652
rect 19852 57598 19854 57650
rect 19854 57598 19906 57650
rect 19906 57598 19908 57650
rect 19852 57596 19908 57598
rect 19628 57260 19684 57316
rect 19404 57036 19460 57092
rect 19180 56924 19236 56980
rect 17388 53788 17444 53844
rect 17276 53676 17332 53732
rect 16044 52834 16100 52836
rect 16044 52782 16046 52834
rect 16046 52782 16098 52834
rect 16098 52782 16100 52834
rect 16044 52780 16100 52782
rect 15932 52444 15988 52500
rect 16044 52332 16100 52388
rect 15260 49644 15316 49700
rect 15372 51996 15428 52052
rect 15260 49308 15316 49364
rect 15260 49026 15316 49028
rect 15260 48974 15262 49026
rect 15262 48974 15314 49026
rect 15314 48974 15316 49026
rect 15260 48972 15316 48974
rect 15148 48748 15204 48804
rect 14924 48636 14980 48692
rect 14364 47516 14420 47572
rect 13692 47234 13748 47236
rect 13692 47182 13694 47234
rect 13694 47182 13746 47234
rect 13746 47182 13748 47234
rect 13692 47180 13748 47182
rect 14476 47404 14532 47460
rect 14924 47964 14980 48020
rect 15148 47570 15204 47572
rect 15148 47518 15150 47570
rect 15150 47518 15202 47570
rect 15202 47518 15204 47570
rect 15148 47516 15204 47518
rect 14812 47180 14868 47236
rect 14476 47068 14532 47124
rect 14364 46956 14420 47012
rect 14140 46898 14196 46900
rect 14140 46846 14142 46898
rect 14142 46846 14194 46898
rect 14194 46846 14196 46898
rect 14140 46844 14196 46846
rect 13916 46674 13972 46676
rect 13916 46622 13918 46674
rect 13918 46622 13970 46674
rect 13970 46622 13972 46674
rect 13916 46620 13972 46622
rect 14252 46620 14308 46676
rect 15260 46674 15316 46676
rect 15260 46622 15262 46674
rect 15262 46622 15314 46674
rect 15314 46622 15316 46674
rect 15260 46620 15316 46622
rect 14140 46284 14196 46340
rect 14588 46284 14644 46340
rect 14252 46172 14308 46228
rect 14028 45836 14084 45892
rect 13916 45778 13972 45780
rect 13916 45726 13918 45778
rect 13918 45726 13970 45778
rect 13970 45726 13972 45778
rect 13916 45724 13972 45726
rect 14028 45388 14084 45444
rect 13804 44492 13860 44548
rect 11900 43148 11956 43204
rect 11564 42364 11620 42420
rect 11788 42588 11844 42644
rect 11228 42028 11284 42084
rect 11452 41916 11508 41972
rect 11116 41132 11172 41188
rect 11228 40514 11284 40516
rect 11228 40462 11230 40514
rect 11230 40462 11282 40514
rect 11282 40462 11284 40514
rect 11228 40460 11284 40462
rect 11116 40290 11172 40292
rect 11116 40238 11118 40290
rect 11118 40238 11170 40290
rect 11170 40238 11172 40290
rect 11116 40236 11172 40238
rect 12124 42978 12180 42980
rect 12124 42926 12126 42978
rect 12126 42926 12178 42978
rect 12178 42926 12180 42978
rect 12124 42924 12180 42926
rect 12348 42812 12404 42868
rect 12348 42588 12404 42644
rect 12124 41916 12180 41972
rect 13580 43708 13636 43764
rect 13804 44044 13860 44100
rect 12908 43538 12964 43540
rect 12908 43486 12910 43538
rect 12910 43486 12962 43538
rect 12962 43486 12964 43538
rect 12908 43484 12964 43486
rect 13356 43484 13412 43540
rect 13020 43426 13076 43428
rect 13020 43374 13022 43426
rect 13022 43374 13074 43426
rect 13074 43374 13076 43426
rect 13020 43372 13076 43374
rect 13356 42588 13412 42644
rect 12460 41580 12516 41636
rect 11564 40796 11620 40852
rect 11676 40626 11732 40628
rect 11676 40574 11678 40626
rect 11678 40574 11730 40626
rect 11730 40574 11732 40626
rect 11676 40572 11732 40574
rect 11340 40236 11396 40292
rect 11564 40348 11620 40404
rect 10220 39228 10276 39284
rect 9996 38892 10052 38948
rect 10444 39004 10500 39060
rect 10108 38668 10164 38724
rect 9772 37938 9828 37940
rect 9772 37886 9774 37938
rect 9774 37886 9826 37938
rect 9826 37886 9828 37938
rect 9772 37884 9828 37886
rect 9548 36988 9604 37044
rect 9660 37100 9716 37156
rect 9436 36540 9492 36596
rect 9324 36482 9380 36484
rect 9324 36430 9326 36482
rect 9326 36430 9378 36482
rect 9378 36430 9380 36482
rect 9324 36428 9380 36430
rect 8988 36092 9044 36148
rect 9324 36092 9380 36148
rect 9324 35420 9380 35476
rect 9548 35644 9604 35700
rect 9100 34188 9156 34244
rect 9212 35308 9268 35364
rect 9212 34300 9268 34356
rect 8988 33740 9044 33796
rect 8876 33404 8932 33460
rect 9212 33122 9268 33124
rect 9212 33070 9214 33122
rect 9214 33070 9266 33122
rect 9266 33070 9268 33122
rect 9212 33068 9268 33070
rect 10332 38220 10388 38276
rect 10220 37996 10276 38052
rect 9996 37378 10052 37380
rect 9996 37326 9998 37378
rect 9998 37326 10050 37378
rect 10050 37326 10052 37378
rect 9996 37324 10052 37326
rect 10444 37996 10500 38052
rect 10668 38892 10724 38948
rect 10668 37826 10724 37828
rect 10668 37774 10670 37826
rect 10670 37774 10722 37826
rect 10722 37774 10724 37826
rect 10668 37772 10724 37774
rect 10220 37212 10276 37268
rect 10220 37042 10276 37044
rect 10220 36990 10222 37042
rect 10222 36990 10274 37042
rect 10274 36990 10276 37042
rect 10220 36988 10276 36990
rect 9996 36876 10052 36932
rect 10556 37490 10612 37492
rect 10556 37438 10558 37490
rect 10558 37438 10610 37490
rect 10610 37438 10612 37490
rect 10556 37436 10612 37438
rect 10668 37324 10724 37380
rect 10556 36988 10612 37044
rect 10668 36876 10724 36932
rect 10108 36482 10164 36484
rect 10108 36430 10110 36482
rect 10110 36430 10162 36482
rect 10162 36430 10164 36482
rect 10108 36428 10164 36430
rect 9884 35980 9940 36036
rect 10108 35756 10164 35812
rect 10108 35420 10164 35476
rect 9772 35196 9828 35252
rect 9884 34972 9940 35028
rect 9996 34188 10052 34244
rect 9548 32732 9604 32788
rect 9660 33292 9716 33348
rect 9100 32562 9156 32564
rect 9100 32510 9102 32562
rect 9102 32510 9154 32562
rect 9154 32510 9156 32562
rect 9100 32508 9156 32510
rect 9212 31948 9268 32004
rect 8428 30380 8484 30436
rect 8316 29036 8372 29092
rect 8540 29148 8596 29204
rect 8428 27858 8484 27860
rect 8428 27806 8430 27858
rect 8430 27806 8482 27858
rect 8482 27806 8484 27858
rect 8428 27804 8484 27806
rect 8316 27468 8372 27524
rect 7868 25788 7924 25844
rect 7868 25452 7924 25508
rect 7420 24780 7476 24836
rect 6524 24108 6580 24164
rect 7308 24108 7364 24164
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 5068 21420 5124 21476
rect 4956 20972 5012 21028
rect 4508 20300 4564 20356
rect 4956 20300 5012 20356
rect 4284 19964 4340 20020
rect 3388 18450 3444 18452
rect 3388 18398 3390 18450
rect 3390 18398 3442 18450
rect 3442 18398 3444 18450
rect 3388 18396 3444 18398
rect 4060 18284 4116 18340
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 5516 20972 5572 21028
rect 5180 19628 5236 19684
rect 5068 19346 5124 19348
rect 5068 19294 5070 19346
rect 5070 19294 5122 19346
rect 5122 19294 5124 19346
rect 5068 19292 5124 19294
rect 4956 19180 5012 19236
rect 4172 18674 4228 18676
rect 4172 18622 4174 18674
rect 4174 18622 4226 18674
rect 4226 18622 4228 18674
rect 4172 18620 4228 18622
rect 4508 18620 4564 18676
rect 2268 17724 2324 17780
rect 4620 18338 4676 18340
rect 4620 18286 4622 18338
rect 4622 18286 4674 18338
rect 4674 18286 4676 18338
rect 4620 18284 4676 18286
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4508 17778 4564 17780
rect 4508 17726 4510 17778
rect 4510 17726 4562 17778
rect 4562 17726 4564 17778
rect 4508 17724 4564 17726
rect 4844 17724 4900 17780
rect 4620 17106 4676 17108
rect 4620 17054 4622 17106
rect 4622 17054 4674 17106
rect 4674 17054 4676 17106
rect 4620 17052 4676 17054
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 5628 20914 5684 20916
rect 5628 20862 5630 20914
rect 5630 20862 5682 20914
rect 5682 20862 5684 20914
rect 5628 20860 5684 20862
rect 6412 22258 6468 22260
rect 6412 22206 6414 22258
rect 6414 22206 6466 22258
rect 6466 22206 6468 22258
rect 6412 22204 6468 22206
rect 6412 21756 6468 21812
rect 6188 21698 6244 21700
rect 6188 21646 6190 21698
rect 6190 21646 6242 21698
rect 6242 21646 6244 21698
rect 6188 21644 6244 21646
rect 5964 21532 6020 21588
rect 6412 20860 6468 20916
rect 5852 19346 5908 19348
rect 5852 19294 5854 19346
rect 5854 19294 5906 19346
rect 5906 19294 5908 19346
rect 5852 19292 5908 19294
rect 5292 16828 5348 16884
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4284 13020 4340 13076
rect 3500 12850 3556 12852
rect 3500 12798 3502 12850
rect 3502 12798 3554 12850
rect 3554 12798 3556 12850
rect 3500 12796 3556 12798
rect 4284 12850 4340 12852
rect 4284 12798 4286 12850
rect 4286 12798 4338 12850
rect 4338 12798 4340 12850
rect 4284 12796 4340 12798
rect 3612 12124 3668 12180
rect 4172 12178 4228 12180
rect 4172 12126 4174 12178
rect 4174 12126 4226 12178
rect 4226 12126 4228 12178
rect 4172 12124 4228 12126
rect 4508 12124 4564 12180
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4844 11340 4900 11396
rect 5068 11116 5124 11172
rect 5628 14642 5684 14644
rect 5628 14590 5630 14642
rect 5630 14590 5682 14642
rect 5682 14590 5684 14642
rect 5628 14588 5684 14590
rect 6076 20188 6132 20244
rect 6188 20636 6244 20692
rect 7084 23938 7140 23940
rect 7084 23886 7086 23938
rect 7086 23886 7138 23938
rect 7138 23886 7140 23938
rect 7084 23884 7140 23886
rect 6636 23154 6692 23156
rect 6636 23102 6638 23154
rect 6638 23102 6690 23154
rect 6690 23102 6692 23154
rect 6636 23100 6692 23102
rect 6972 23548 7028 23604
rect 6636 21868 6692 21924
rect 6748 22428 6804 22484
rect 6636 21586 6692 21588
rect 6636 21534 6638 21586
rect 6638 21534 6690 21586
rect 6690 21534 6692 21586
rect 6636 21532 6692 21534
rect 6636 20300 6692 20356
rect 6524 19292 6580 19348
rect 6636 19628 6692 19684
rect 6860 21756 6916 21812
rect 6860 20748 6916 20804
rect 7644 24108 7700 24164
rect 7868 23548 7924 23604
rect 7868 23324 7924 23380
rect 8092 24668 8148 24724
rect 8988 30994 9044 30996
rect 8988 30942 8990 30994
rect 8990 30942 9042 30994
rect 9042 30942 9044 30994
rect 8988 30940 9044 30942
rect 10108 34130 10164 34132
rect 10108 34078 10110 34130
rect 10110 34078 10162 34130
rect 10162 34078 10164 34130
rect 10108 34076 10164 34078
rect 10444 36316 10500 36372
rect 10332 35308 10388 35364
rect 10108 33906 10164 33908
rect 10108 33854 10110 33906
rect 10110 33854 10162 33906
rect 10162 33854 10164 33906
rect 10108 33852 10164 33854
rect 9660 31612 9716 31668
rect 9324 30940 9380 30996
rect 8876 30380 8932 30436
rect 8876 30156 8932 30212
rect 9660 31276 9716 31332
rect 9772 30492 9828 30548
rect 9884 31948 9940 32004
rect 9212 30098 9268 30100
rect 9212 30046 9214 30098
rect 9214 30046 9266 30098
rect 9266 30046 9268 30098
rect 9212 30044 9268 30046
rect 10220 31948 10276 32004
rect 10108 31836 10164 31892
rect 10892 37996 10948 38052
rect 10892 36988 10948 37044
rect 12460 41020 12516 41076
rect 12012 40460 12068 40516
rect 12124 40402 12180 40404
rect 12124 40350 12126 40402
rect 12126 40350 12178 40402
rect 12178 40350 12180 40402
rect 12124 40348 12180 40350
rect 11676 40012 11732 40068
rect 11452 39506 11508 39508
rect 11452 39454 11454 39506
rect 11454 39454 11506 39506
rect 11506 39454 11508 39506
rect 11452 39452 11508 39454
rect 11676 39452 11732 39508
rect 11564 39340 11620 39396
rect 11116 37826 11172 37828
rect 11116 37774 11118 37826
rect 11118 37774 11170 37826
rect 11170 37774 11172 37826
rect 11116 37772 11172 37774
rect 11116 37548 11172 37604
rect 11900 39452 11956 39508
rect 11676 38108 11732 38164
rect 11228 37100 11284 37156
rect 10892 36594 10948 36596
rect 10892 36542 10894 36594
rect 10894 36542 10946 36594
rect 10946 36542 10948 36594
rect 10892 36540 10948 36542
rect 10780 36428 10836 36484
rect 10892 36204 10948 36260
rect 10780 35698 10836 35700
rect 10780 35646 10782 35698
rect 10782 35646 10834 35698
rect 10834 35646 10836 35698
rect 10780 35644 10836 35646
rect 10444 31388 10500 31444
rect 10556 31500 10612 31556
rect 10444 31164 10500 31220
rect 9996 31052 10052 31108
rect 10108 30994 10164 30996
rect 10108 30942 10110 30994
rect 10110 30942 10162 30994
rect 10162 30942 10164 30994
rect 10108 30940 10164 30942
rect 10332 30994 10388 30996
rect 10332 30942 10334 30994
rect 10334 30942 10386 30994
rect 10386 30942 10388 30994
rect 10332 30940 10388 30942
rect 9324 28924 9380 28980
rect 8988 27970 9044 27972
rect 8988 27918 8990 27970
rect 8990 27918 9042 27970
rect 9042 27918 9044 27970
rect 8988 27916 9044 27918
rect 9100 28364 9156 28420
rect 8652 27244 8708 27300
rect 8876 27804 8932 27860
rect 8764 27132 8820 27188
rect 8540 26796 8596 26852
rect 8316 23212 8372 23268
rect 8540 26178 8596 26180
rect 8540 26126 8542 26178
rect 8542 26126 8594 26178
rect 8594 26126 8596 26178
rect 8540 26124 8596 26126
rect 9436 26796 9492 26852
rect 9660 28530 9716 28532
rect 9660 28478 9662 28530
rect 9662 28478 9714 28530
rect 9714 28478 9716 28530
rect 9660 28476 9716 28478
rect 9884 29372 9940 29428
rect 9996 29148 10052 29204
rect 10556 30940 10612 30996
rect 10444 29986 10500 29988
rect 10444 29934 10446 29986
rect 10446 29934 10498 29986
rect 10498 29934 10500 29986
rect 10444 29932 10500 29934
rect 10108 28140 10164 28196
rect 9772 27916 9828 27972
rect 10108 27916 10164 27972
rect 9996 27858 10052 27860
rect 9996 27806 9998 27858
rect 9998 27806 10050 27858
rect 10050 27806 10052 27858
rect 9996 27804 10052 27806
rect 9996 27020 10052 27076
rect 9100 25676 9156 25732
rect 9212 26124 9268 26180
rect 8876 24834 8932 24836
rect 8876 24782 8878 24834
rect 8878 24782 8930 24834
rect 8930 24782 8932 24834
rect 8876 24780 8932 24782
rect 9324 25340 9380 25396
rect 8652 23938 8708 23940
rect 8652 23886 8654 23938
rect 8654 23886 8706 23938
rect 8706 23886 8708 23938
rect 8652 23884 8708 23886
rect 8764 23548 8820 23604
rect 8988 23660 9044 23716
rect 8988 23324 9044 23380
rect 7420 21644 7476 21700
rect 7308 20972 7364 21028
rect 7308 20802 7364 20804
rect 7308 20750 7310 20802
rect 7310 20750 7362 20802
rect 7362 20750 7364 20802
rect 7308 20748 7364 20750
rect 6860 20076 6916 20132
rect 7196 20188 7252 20244
rect 8092 21644 8148 21700
rect 8204 21308 8260 21364
rect 8540 21308 8596 21364
rect 7980 21084 8036 21140
rect 7980 20748 8036 20804
rect 8428 21196 8484 21252
rect 8428 20578 8484 20580
rect 8428 20526 8430 20578
rect 8430 20526 8482 20578
rect 8482 20526 8484 20578
rect 8428 20524 8484 20526
rect 7084 20018 7140 20020
rect 7084 19966 7086 20018
rect 7086 19966 7138 20018
rect 7138 19966 7140 20018
rect 7084 19964 7140 19966
rect 6636 18956 6692 19012
rect 6076 18620 6132 18676
rect 6748 18284 6804 18340
rect 6524 17778 6580 17780
rect 6524 17726 6526 17778
rect 6526 17726 6578 17778
rect 6578 17726 6580 17778
rect 6524 17724 6580 17726
rect 6412 16210 6468 16212
rect 6412 16158 6414 16210
rect 6414 16158 6466 16210
rect 6466 16158 6468 16210
rect 6412 16156 6468 16158
rect 7084 18508 7140 18564
rect 6972 16156 7028 16212
rect 7532 19404 7588 19460
rect 7532 19180 7588 19236
rect 5740 13020 5796 13076
rect 5404 12178 5460 12180
rect 5404 12126 5406 12178
rect 5406 12126 5458 12178
rect 5458 12126 5460 12178
rect 5404 12124 5460 12126
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4956 9714 5012 9716
rect 4956 9662 4958 9714
rect 4958 9662 5010 9714
rect 5010 9662 5012 9714
rect 4956 9660 5012 9662
rect 4844 9266 4900 9268
rect 4844 9214 4846 9266
rect 4846 9214 4898 9266
rect 4898 9214 4900 9266
rect 4844 9212 4900 9214
rect 4284 9042 4340 9044
rect 4284 8990 4286 9042
rect 4286 8990 4338 9042
rect 4338 8990 4340 9042
rect 4284 8988 4340 8990
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 5740 9714 5796 9716
rect 5740 9662 5742 9714
rect 5742 9662 5794 9714
rect 5794 9662 5796 9714
rect 5740 9660 5796 9662
rect 5292 8316 5348 8372
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4844 6578 4900 6580
rect 4844 6526 4846 6578
rect 4846 6526 4898 6578
rect 4898 6526 4900 6578
rect 4844 6524 4900 6526
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 6748 15148 6804 15204
rect 7532 17724 7588 17780
rect 7980 19346 8036 19348
rect 7980 19294 7982 19346
rect 7982 19294 8034 19346
rect 8034 19294 8036 19346
rect 7980 19292 8036 19294
rect 8204 19068 8260 19124
rect 8428 19010 8484 19012
rect 8428 18958 8430 19010
rect 8430 18958 8482 19010
rect 8482 18958 8484 19010
rect 8428 18956 8484 18958
rect 7980 18396 8036 18452
rect 7868 17778 7924 17780
rect 7868 17726 7870 17778
rect 7870 17726 7922 17778
rect 7922 17726 7924 17778
rect 7868 17724 7924 17726
rect 8428 17778 8484 17780
rect 8428 17726 8430 17778
rect 8430 17726 8482 17778
rect 8482 17726 8484 17778
rect 8428 17724 8484 17726
rect 8540 18396 8596 18452
rect 7644 17052 7700 17108
rect 8988 21810 9044 21812
rect 8988 21758 8990 21810
rect 8990 21758 9042 21810
rect 9042 21758 9044 21810
rect 8988 21756 9044 21758
rect 8988 21420 9044 21476
rect 9100 21644 9156 21700
rect 8876 20748 8932 20804
rect 8988 20690 9044 20692
rect 8988 20638 8990 20690
rect 8990 20638 9042 20690
rect 9042 20638 9044 20690
rect 8988 20636 9044 20638
rect 9660 26348 9716 26404
rect 9660 25618 9716 25620
rect 9660 25566 9662 25618
rect 9662 25566 9714 25618
rect 9714 25566 9716 25618
rect 9660 25564 9716 25566
rect 9772 26236 9828 26292
rect 10444 29596 10500 29652
rect 10444 28252 10500 28308
rect 10332 27580 10388 27636
rect 10332 27186 10388 27188
rect 10332 27134 10334 27186
rect 10334 27134 10386 27186
rect 10386 27134 10388 27186
rect 10332 27132 10388 27134
rect 10332 26514 10388 26516
rect 10332 26462 10334 26514
rect 10334 26462 10386 26514
rect 10386 26462 10388 26514
rect 10332 26460 10388 26462
rect 10220 26012 10276 26068
rect 11004 35196 11060 35252
rect 11004 34914 11060 34916
rect 11004 34862 11006 34914
rect 11006 34862 11058 34914
rect 11058 34862 11060 34914
rect 11004 34860 11060 34862
rect 10668 34636 10724 34692
rect 11564 36764 11620 36820
rect 11452 36428 11508 36484
rect 11340 34300 11396 34356
rect 10780 34130 10836 34132
rect 10780 34078 10782 34130
rect 10782 34078 10834 34130
rect 10834 34078 10836 34130
rect 10780 34076 10836 34078
rect 10668 33964 10724 34020
rect 10780 33628 10836 33684
rect 11452 32620 11508 32676
rect 11228 32396 11284 32452
rect 10780 31724 10836 31780
rect 11004 30604 11060 30660
rect 11228 31164 11284 31220
rect 11228 30828 11284 30884
rect 11116 30492 11172 30548
rect 11116 30268 11172 30324
rect 10668 30156 10724 30212
rect 11004 30210 11060 30212
rect 11004 30158 11006 30210
rect 11006 30158 11058 30210
rect 11058 30158 11060 30210
rect 11004 30156 11060 30158
rect 11228 29932 11284 29988
rect 11340 30156 11396 30212
rect 11116 29596 11172 29652
rect 11452 29596 11508 29652
rect 10780 29538 10836 29540
rect 10780 29486 10782 29538
rect 10782 29486 10834 29538
rect 10834 29486 10836 29538
rect 10780 29484 10836 29486
rect 11004 29314 11060 29316
rect 11004 29262 11006 29314
rect 11006 29262 11058 29314
rect 11058 29262 11060 29314
rect 11004 29260 11060 29262
rect 11228 29202 11284 29204
rect 11228 29150 11230 29202
rect 11230 29150 11282 29202
rect 11282 29150 11284 29202
rect 11228 29148 11284 29150
rect 10668 28476 10724 28532
rect 10780 28418 10836 28420
rect 10780 28366 10782 28418
rect 10782 28366 10834 28418
rect 10834 28366 10836 28418
rect 10780 28364 10836 28366
rect 11004 27916 11060 27972
rect 10556 26908 10612 26964
rect 10892 26962 10948 26964
rect 10892 26910 10894 26962
rect 10894 26910 10946 26962
rect 10946 26910 10948 26962
rect 10892 26908 10948 26910
rect 10444 25900 10500 25956
rect 9996 25340 10052 25396
rect 11004 26290 11060 26292
rect 11004 26238 11006 26290
rect 11006 26238 11058 26290
rect 11058 26238 11060 26290
rect 11004 26236 11060 26238
rect 10668 26012 10724 26068
rect 10444 25282 10500 25284
rect 10444 25230 10446 25282
rect 10446 25230 10498 25282
rect 10498 25230 10500 25282
rect 10444 25228 10500 25230
rect 10220 25116 10276 25172
rect 10444 24834 10500 24836
rect 10444 24782 10446 24834
rect 10446 24782 10498 24834
rect 10498 24782 10500 24834
rect 10444 24780 10500 24782
rect 9996 24668 10052 24724
rect 9772 23996 9828 24052
rect 9884 24108 9940 24164
rect 9548 23100 9604 23156
rect 9660 21756 9716 21812
rect 9436 21644 9492 21700
rect 9884 22092 9940 22148
rect 9436 20802 9492 20804
rect 9436 20750 9438 20802
rect 9438 20750 9490 20802
rect 9490 20750 9492 20802
rect 9436 20748 9492 20750
rect 7756 16828 7812 16884
rect 7308 15260 7364 15316
rect 6412 14642 6468 14644
rect 6412 14590 6414 14642
rect 6414 14590 6466 14642
rect 6466 14590 6468 14642
rect 6412 14588 6468 14590
rect 6860 14642 6916 14644
rect 6860 14590 6862 14642
rect 6862 14590 6914 14642
rect 6914 14590 6916 14642
rect 6860 14588 6916 14590
rect 8540 16828 8596 16884
rect 9772 20914 9828 20916
rect 9772 20862 9774 20914
rect 9774 20862 9826 20914
rect 9826 20862 9828 20914
rect 9772 20860 9828 20862
rect 10220 24332 10276 24388
rect 10556 24108 10612 24164
rect 10556 23826 10612 23828
rect 10556 23774 10558 23826
rect 10558 23774 10610 23826
rect 10610 23774 10612 23826
rect 10556 23772 10612 23774
rect 10892 25900 10948 25956
rect 10780 25116 10836 25172
rect 10780 23660 10836 23716
rect 11228 26796 11284 26852
rect 12012 39228 12068 39284
rect 12460 39506 12516 39508
rect 12460 39454 12462 39506
rect 12462 39454 12514 39506
rect 12514 39454 12516 39506
rect 12460 39452 12516 39454
rect 12236 39340 12292 39396
rect 12684 39900 12740 39956
rect 13020 41916 13076 41972
rect 13244 42140 13300 42196
rect 13580 43372 13636 43428
rect 13468 42194 13524 42196
rect 13468 42142 13470 42194
rect 13470 42142 13522 42194
rect 13522 42142 13524 42194
rect 13468 42140 13524 42142
rect 13692 42028 13748 42084
rect 12908 41244 12964 41300
rect 13020 41468 13076 41524
rect 13356 41244 13412 41300
rect 13020 40796 13076 40852
rect 13020 40514 13076 40516
rect 13020 40462 13022 40514
rect 13022 40462 13074 40514
rect 13074 40462 13076 40514
rect 13020 40460 13076 40462
rect 12908 39730 12964 39732
rect 12908 39678 12910 39730
rect 12910 39678 12962 39730
rect 12962 39678 12964 39730
rect 12908 39676 12964 39678
rect 12572 39228 12628 39284
rect 12124 37996 12180 38052
rect 11900 37772 11956 37828
rect 12124 37548 12180 37604
rect 12012 37324 12068 37380
rect 12124 37212 12180 37268
rect 11676 34524 11732 34580
rect 11788 35644 11844 35700
rect 11900 35196 11956 35252
rect 12124 36988 12180 37044
rect 12012 35084 12068 35140
rect 12124 35026 12180 35028
rect 12124 34974 12126 35026
rect 12126 34974 12178 35026
rect 12178 34974 12180 35026
rect 12124 34972 12180 34974
rect 12460 39058 12516 39060
rect 12460 39006 12462 39058
rect 12462 39006 12514 39058
rect 12514 39006 12516 39058
rect 12460 39004 12516 39006
rect 12348 38834 12404 38836
rect 12348 38782 12350 38834
rect 12350 38782 12402 38834
rect 12402 38782 12404 38834
rect 12348 38780 12404 38782
rect 12684 38668 12740 38724
rect 13244 39228 13300 39284
rect 12908 38220 12964 38276
rect 12572 38108 12628 38164
rect 12572 37660 12628 37716
rect 12796 37548 12852 37604
rect 12684 37266 12740 37268
rect 12684 37214 12686 37266
rect 12686 37214 12738 37266
rect 12738 37214 12740 37266
rect 12684 37212 12740 37214
rect 12572 37100 12628 37156
rect 12796 36652 12852 36708
rect 12908 36428 12964 36484
rect 12684 36092 12740 36148
rect 12348 35698 12404 35700
rect 12348 35646 12350 35698
rect 12350 35646 12402 35698
rect 12402 35646 12404 35698
rect 12348 35644 12404 35646
rect 11900 34524 11956 34580
rect 11900 34354 11956 34356
rect 11900 34302 11902 34354
rect 11902 34302 11954 34354
rect 11954 34302 11956 34354
rect 11900 34300 11956 34302
rect 12236 34354 12292 34356
rect 12236 34302 12238 34354
rect 12238 34302 12290 34354
rect 12290 34302 12292 34354
rect 12236 34300 12292 34302
rect 11788 34188 11844 34244
rect 12348 33628 12404 33684
rect 12572 34690 12628 34692
rect 12572 34638 12574 34690
rect 12574 34638 12626 34690
rect 12626 34638 12628 34690
rect 12572 34636 12628 34638
rect 12908 36092 12964 36148
rect 13692 41020 13748 41076
rect 13692 40348 13748 40404
rect 13692 39564 13748 39620
rect 13580 39394 13636 39396
rect 13580 39342 13582 39394
rect 13582 39342 13634 39394
rect 13634 39342 13636 39394
rect 13580 39340 13636 39342
rect 13580 37548 13636 37604
rect 14476 45724 14532 45780
rect 14364 44604 14420 44660
rect 14364 44044 14420 44100
rect 14252 43484 14308 43540
rect 13916 43426 13972 43428
rect 13916 43374 13918 43426
rect 13918 43374 13970 43426
rect 13970 43374 13972 43426
rect 13916 43372 13972 43374
rect 13916 42812 13972 42868
rect 14252 42866 14308 42868
rect 14252 42814 14254 42866
rect 14254 42814 14306 42866
rect 14306 42814 14308 42866
rect 14252 42812 14308 42814
rect 14364 42754 14420 42756
rect 14364 42702 14366 42754
rect 14366 42702 14418 42754
rect 14418 42702 14420 42754
rect 14364 42700 14420 42702
rect 14140 42642 14196 42644
rect 14140 42590 14142 42642
rect 14142 42590 14194 42642
rect 14194 42590 14196 42642
rect 14140 42588 14196 42590
rect 14140 42140 14196 42196
rect 14364 41858 14420 41860
rect 14364 41806 14366 41858
rect 14366 41806 14418 41858
rect 14418 41806 14420 41858
rect 14364 41804 14420 41806
rect 14812 45052 14868 45108
rect 15932 52108 15988 52164
rect 15820 51602 15876 51604
rect 15820 51550 15822 51602
rect 15822 51550 15874 51602
rect 15874 51550 15876 51602
rect 15820 51548 15876 51550
rect 16044 51324 16100 51380
rect 15820 50764 15876 50820
rect 15596 50482 15652 50484
rect 15596 50430 15598 50482
rect 15598 50430 15650 50482
rect 15650 50430 15652 50482
rect 15596 50428 15652 50430
rect 15596 50204 15652 50260
rect 15708 50034 15764 50036
rect 15708 49982 15710 50034
rect 15710 49982 15762 50034
rect 15762 49982 15764 50034
rect 15708 49980 15764 49982
rect 16492 52668 16548 52724
rect 16492 50988 16548 51044
rect 16156 50204 16212 50260
rect 17052 53004 17108 53060
rect 16940 52220 16996 52276
rect 16716 50818 16772 50820
rect 16716 50766 16718 50818
rect 16718 50766 16770 50818
rect 16770 50766 16772 50818
rect 16716 50764 16772 50766
rect 16380 49980 16436 50036
rect 17164 53228 17220 53284
rect 17276 52892 17332 52948
rect 17276 52108 17332 52164
rect 17052 50540 17108 50596
rect 17164 51996 17220 52052
rect 17164 51548 17220 51604
rect 16940 49868 16996 49924
rect 16044 49644 16100 49700
rect 15484 49308 15540 49364
rect 15596 49026 15652 49028
rect 15596 48974 15598 49026
rect 15598 48974 15650 49026
rect 15650 48974 15652 49026
rect 15596 48972 15652 48974
rect 16940 49698 16996 49700
rect 16940 49646 16942 49698
rect 16942 49646 16994 49698
rect 16994 49646 16996 49698
rect 16940 49644 16996 49646
rect 16492 49196 16548 49252
rect 16044 48802 16100 48804
rect 16044 48750 16046 48802
rect 16046 48750 16098 48802
rect 16098 48750 16100 48802
rect 16044 48748 16100 48750
rect 16380 49084 16436 49140
rect 15596 48524 15652 48580
rect 15484 48412 15540 48468
rect 14924 44210 14980 44212
rect 14924 44158 14926 44210
rect 14926 44158 14978 44210
rect 14978 44158 14980 44210
rect 14924 44156 14980 44158
rect 15484 47964 15540 48020
rect 14700 43762 14756 43764
rect 14700 43710 14702 43762
rect 14702 43710 14754 43762
rect 14754 43710 14756 43762
rect 14700 43708 14756 43710
rect 14588 41970 14644 41972
rect 14588 41918 14590 41970
rect 14590 41918 14642 41970
rect 14642 41918 14644 41970
rect 14588 41916 14644 41918
rect 14140 41186 14196 41188
rect 14140 41134 14142 41186
rect 14142 41134 14194 41186
rect 14194 41134 14196 41186
rect 14140 41132 14196 41134
rect 14252 41074 14308 41076
rect 14252 41022 14254 41074
rect 14254 41022 14306 41074
rect 14306 41022 14308 41074
rect 14252 41020 14308 41022
rect 13916 40626 13972 40628
rect 13916 40574 13918 40626
rect 13918 40574 13970 40626
rect 13970 40574 13972 40626
rect 13916 40572 13972 40574
rect 14028 39116 14084 39172
rect 14364 40572 14420 40628
rect 14476 40684 14532 40740
rect 14364 39788 14420 39844
rect 15708 48636 15764 48692
rect 16156 48524 16212 48580
rect 15932 48242 15988 48244
rect 15932 48190 15934 48242
rect 15934 48190 15986 48242
rect 15986 48190 15988 48242
rect 15932 48188 15988 48190
rect 15596 47516 15652 47572
rect 15708 47458 15764 47460
rect 15708 47406 15710 47458
rect 15710 47406 15762 47458
rect 15762 47406 15764 47458
rect 15708 47404 15764 47406
rect 15708 47068 15764 47124
rect 15596 45330 15652 45332
rect 15596 45278 15598 45330
rect 15598 45278 15650 45330
rect 15650 45278 15652 45330
rect 15596 45276 15652 45278
rect 15932 47068 15988 47124
rect 15820 46732 15876 46788
rect 16940 49138 16996 49140
rect 16940 49086 16942 49138
rect 16942 49086 16994 49138
rect 16994 49086 16996 49138
rect 16940 49084 16996 49086
rect 16044 45778 16100 45780
rect 16044 45726 16046 45778
rect 16046 45726 16098 45778
rect 16098 45726 16100 45778
rect 16044 45724 16100 45726
rect 15148 43036 15204 43092
rect 14924 42194 14980 42196
rect 14924 42142 14926 42194
rect 14926 42142 14978 42194
rect 14978 42142 14980 42194
rect 14924 42140 14980 42142
rect 15036 41692 15092 41748
rect 15260 41580 15316 41636
rect 15260 41356 15316 41412
rect 15484 43260 15540 43316
rect 16156 44716 16212 44772
rect 16492 48802 16548 48804
rect 16492 48750 16494 48802
rect 16494 48750 16546 48802
rect 16546 48750 16548 48802
rect 16492 48748 16548 48750
rect 16940 48466 16996 48468
rect 16940 48414 16942 48466
rect 16942 48414 16994 48466
rect 16994 48414 16996 48466
rect 16940 48412 16996 48414
rect 17612 55970 17668 55972
rect 17612 55918 17614 55970
rect 17614 55918 17666 55970
rect 17666 55918 17668 55970
rect 17612 55916 17668 55918
rect 18508 55580 18564 55636
rect 18172 55468 18228 55524
rect 18732 55298 18788 55300
rect 18732 55246 18734 55298
rect 18734 55246 18786 55298
rect 18786 55246 18788 55298
rect 18732 55244 18788 55246
rect 19180 55244 19236 55300
rect 19068 55186 19124 55188
rect 19068 55134 19070 55186
rect 19070 55134 19122 55186
rect 19122 55134 19124 55186
rect 19068 55132 19124 55134
rect 17836 54908 17892 54964
rect 17724 54236 17780 54292
rect 19292 54572 19348 54628
rect 19516 55858 19572 55860
rect 19516 55806 19518 55858
rect 19518 55806 19570 55858
rect 19570 55806 19572 55858
rect 19516 55804 19572 55806
rect 20972 58210 21028 58212
rect 20972 58158 20974 58210
rect 20974 58158 21026 58210
rect 21026 58158 21028 58210
rect 20972 58156 21028 58158
rect 20524 57148 20580 57204
rect 20188 57036 20244 57092
rect 19852 56642 19908 56644
rect 19852 56590 19854 56642
rect 19854 56590 19906 56642
rect 19906 56590 19908 56642
rect 19852 56588 19908 56590
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 20076 55858 20132 55860
rect 20076 55806 20078 55858
rect 20078 55806 20130 55858
rect 20130 55806 20132 55858
rect 20076 55804 20132 55806
rect 20188 55692 20244 55748
rect 19964 55298 20020 55300
rect 19964 55246 19966 55298
rect 19966 55246 20018 55298
rect 20018 55246 20020 55298
rect 19964 55244 20020 55246
rect 19740 55132 19796 55188
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 19628 54684 19684 54740
rect 18508 53842 18564 53844
rect 18508 53790 18510 53842
rect 18510 53790 18562 53842
rect 18562 53790 18564 53842
rect 18508 53788 18564 53790
rect 18060 52892 18116 52948
rect 17836 52108 17892 52164
rect 17724 51436 17780 51492
rect 17612 51212 17668 51268
rect 17612 50764 17668 50820
rect 18172 51996 18228 52052
rect 18284 52780 18340 52836
rect 18284 52332 18340 52388
rect 18284 51884 18340 51940
rect 18732 53676 18788 53732
rect 19516 54572 19572 54628
rect 19404 54124 19460 54180
rect 19516 53900 19572 53956
rect 19628 53788 19684 53844
rect 20188 54684 20244 54740
rect 19964 54572 20020 54628
rect 19068 53564 19124 53620
rect 19516 53340 19572 53396
rect 19836 53338 19892 53340
rect 19068 53228 19124 53284
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 19852 53058 19908 53060
rect 19852 53006 19854 53058
rect 19854 53006 19906 53058
rect 19906 53006 19908 53058
rect 19852 53004 19908 53006
rect 18956 52834 19012 52836
rect 18956 52782 18958 52834
rect 18958 52782 19010 52834
rect 19010 52782 19012 52834
rect 18956 52780 19012 52782
rect 17276 49868 17332 49924
rect 17836 50204 17892 50260
rect 17724 50092 17780 50148
rect 18172 50764 18228 50820
rect 18396 50540 18452 50596
rect 18172 50204 18228 50260
rect 17612 49756 17668 49812
rect 17388 49644 17444 49700
rect 18060 49308 18116 49364
rect 17500 49196 17556 49252
rect 16604 46674 16660 46676
rect 16604 46622 16606 46674
rect 16606 46622 16658 46674
rect 16658 46622 16660 46674
rect 16604 46620 16660 46622
rect 16492 45836 16548 45892
rect 16604 45388 16660 45444
rect 16492 44994 16548 44996
rect 16492 44942 16494 44994
rect 16494 44942 16546 44994
rect 16546 44942 16548 44994
rect 16492 44940 16548 44942
rect 16156 44492 16212 44548
rect 15820 44322 15876 44324
rect 15820 44270 15822 44322
rect 15822 44270 15874 44322
rect 15874 44270 15876 44322
rect 15820 44268 15876 44270
rect 15708 44044 15764 44100
rect 15820 43932 15876 43988
rect 15596 42252 15652 42308
rect 15596 41970 15652 41972
rect 15596 41918 15598 41970
rect 15598 41918 15650 41970
rect 15650 41918 15652 41970
rect 15596 41916 15652 41918
rect 14700 40572 14756 40628
rect 15036 41020 15092 41076
rect 15372 41020 15428 41076
rect 14812 39900 14868 39956
rect 14140 39004 14196 39060
rect 14028 38892 14084 38948
rect 13804 37548 13860 37604
rect 13132 34972 13188 35028
rect 13580 37266 13636 37268
rect 13580 37214 13582 37266
rect 13582 37214 13634 37266
rect 13634 37214 13636 37266
rect 13580 37212 13636 37214
rect 13020 34636 13076 34692
rect 13356 36764 13412 36820
rect 13692 37154 13748 37156
rect 13692 37102 13694 37154
rect 13694 37102 13746 37154
rect 13746 37102 13748 37154
rect 13692 37100 13748 37102
rect 13580 36652 13636 36708
rect 13916 36988 13972 37044
rect 13804 36652 13860 36708
rect 13804 36370 13860 36372
rect 13804 36318 13806 36370
rect 13806 36318 13858 36370
rect 13858 36318 13860 36370
rect 13804 36316 13860 36318
rect 13468 35922 13524 35924
rect 13468 35870 13470 35922
rect 13470 35870 13522 35922
rect 13522 35870 13524 35922
rect 13468 35868 13524 35870
rect 13356 35644 13412 35700
rect 12796 34242 12852 34244
rect 12796 34190 12798 34242
rect 12798 34190 12850 34242
rect 12850 34190 12852 34242
rect 12796 34188 12852 34190
rect 13020 33852 13076 33908
rect 12908 33516 12964 33572
rect 12460 33292 12516 33348
rect 11676 32396 11732 32452
rect 11676 31724 11732 31780
rect 12124 32844 12180 32900
rect 12348 32450 12404 32452
rect 12348 32398 12350 32450
rect 12350 32398 12402 32450
rect 12402 32398 12404 32450
rect 12348 32396 12404 32398
rect 12572 32956 12628 33012
rect 12572 32060 12628 32116
rect 12684 32508 12740 32564
rect 12012 31836 12068 31892
rect 12012 31554 12068 31556
rect 12012 31502 12014 31554
rect 12014 31502 12066 31554
rect 12066 31502 12068 31554
rect 12012 31500 12068 31502
rect 12236 31388 12292 31444
rect 11900 30940 11956 30996
rect 12124 31276 12180 31332
rect 11676 30268 11732 30324
rect 11788 30492 11844 30548
rect 11676 29708 11732 29764
rect 11676 29538 11732 29540
rect 11676 29486 11678 29538
rect 11678 29486 11730 29538
rect 11730 29486 11732 29538
rect 11676 29484 11732 29486
rect 11900 30268 11956 30324
rect 11788 28754 11844 28756
rect 11788 28702 11790 28754
rect 11790 28702 11842 28754
rect 11842 28702 11844 28754
rect 11788 28700 11844 28702
rect 12460 31276 12516 31332
rect 12572 31500 12628 31556
rect 13244 33740 13300 33796
rect 12908 31724 12964 31780
rect 13132 31612 13188 31668
rect 13132 30268 13188 30324
rect 12348 30044 12404 30100
rect 12908 30044 12964 30100
rect 12236 29708 12292 29764
rect 12796 29820 12852 29876
rect 12684 29650 12740 29652
rect 12684 29598 12686 29650
rect 12686 29598 12738 29650
rect 12738 29598 12740 29650
rect 12684 29596 12740 29598
rect 12796 28700 12852 28756
rect 12572 28588 12628 28644
rect 12348 28530 12404 28532
rect 12348 28478 12350 28530
rect 12350 28478 12402 28530
rect 12402 28478 12404 28530
rect 12348 28476 12404 28478
rect 12908 29484 12964 29540
rect 13468 35196 13524 35252
rect 13468 33740 13524 33796
rect 13692 35810 13748 35812
rect 13692 35758 13694 35810
rect 13694 35758 13746 35810
rect 13746 35758 13748 35810
rect 13692 35756 13748 35758
rect 13692 34300 13748 34356
rect 13804 35532 13860 35588
rect 13692 33740 13748 33796
rect 13916 35308 13972 35364
rect 13804 33180 13860 33236
rect 14476 38946 14532 38948
rect 14476 38894 14478 38946
rect 14478 38894 14530 38946
rect 14530 38894 14532 38946
rect 14476 38892 14532 38894
rect 14252 38220 14308 38276
rect 14364 37548 14420 37604
rect 14252 36652 14308 36708
rect 15260 40514 15316 40516
rect 15260 40462 15262 40514
rect 15262 40462 15314 40514
rect 15314 40462 15316 40514
rect 15260 40460 15316 40462
rect 15372 40124 15428 40180
rect 15372 39788 15428 39844
rect 15148 39394 15204 39396
rect 15148 39342 15150 39394
rect 15150 39342 15202 39394
rect 15202 39342 15204 39394
rect 15148 39340 15204 39342
rect 15036 39116 15092 39172
rect 14812 38780 14868 38836
rect 14924 39004 14980 39060
rect 15484 39058 15540 39060
rect 15484 39006 15486 39058
rect 15486 39006 15538 39058
rect 15538 39006 15540 39058
rect 15484 39004 15540 39006
rect 15372 38946 15428 38948
rect 15372 38894 15374 38946
rect 15374 38894 15426 38946
rect 15426 38894 15428 38946
rect 15372 38892 15428 38894
rect 16380 44098 16436 44100
rect 16380 44046 16382 44098
rect 16382 44046 16434 44098
rect 16434 44046 16436 44098
rect 16380 44044 16436 44046
rect 16156 43260 16212 43316
rect 16268 43650 16324 43652
rect 16268 43598 16270 43650
rect 16270 43598 16322 43650
rect 16322 43598 16324 43650
rect 16268 43596 16324 43598
rect 16156 43036 16212 43092
rect 16044 42642 16100 42644
rect 16044 42590 16046 42642
rect 16046 42590 16098 42642
rect 16098 42590 16100 42642
rect 16044 42588 16100 42590
rect 15932 42530 15988 42532
rect 15932 42478 15934 42530
rect 15934 42478 15986 42530
rect 15986 42478 15988 42530
rect 15932 42476 15988 42478
rect 16044 41580 16100 41636
rect 15708 39340 15764 39396
rect 15596 38892 15652 38948
rect 14476 36540 14532 36596
rect 14588 36652 14644 36708
rect 14476 36370 14532 36372
rect 14476 36318 14478 36370
rect 14478 36318 14530 36370
rect 14530 36318 14532 36370
rect 14476 36316 14532 36318
rect 14364 36204 14420 36260
rect 14252 35644 14308 35700
rect 14588 35644 14644 35700
rect 14252 35084 14308 35140
rect 14252 34860 14308 34916
rect 14028 33964 14084 34020
rect 14476 34802 14532 34804
rect 14476 34750 14478 34802
rect 14478 34750 14530 34802
rect 14530 34750 14532 34802
rect 14476 34748 14532 34750
rect 13916 32844 13972 32900
rect 13804 32786 13860 32788
rect 13804 32734 13806 32786
rect 13806 32734 13858 32786
rect 13858 32734 13860 32786
rect 13804 32732 13860 32734
rect 13468 32674 13524 32676
rect 13468 32622 13470 32674
rect 13470 32622 13522 32674
rect 13522 32622 13524 32674
rect 13468 32620 13524 32622
rect 13580 32508 13636 32564
rect 13692 31836 13748 31892
rect 13244 29538 13300 29540
rect 13244 29486 13246 29538
rect 13246 29486 13298 29538
rect 13298 29486 13300 29538
rect 13244 29484 13300 29486
rect 13020 28700 13076 28756
rect 13132 28812 13188 28868
rect 12124 27186 12180 27188
rect 12124 27134 12126 27186
rect 12126 27134 12178 27186
rect 12178 27134 12180 27186
rect 12124 27132 12180 27134
rect 12012 27074 12068 27076
rect 12012 27022 12014 27074
rect 12014 27022 12066 27074
rect 12066 27022 12068 27074
rect 12012 27020 12068 27022
rect 11564 26684 11620 26740
rect 11676 26796 11732 26852
rect 11452 26348 11508 26404
rect 11452 26178 11508 26180
rect 11452 26126 11454 26178
rect 11454 26126 11506 26178
rect 11506 26126 11508 26178
rect 11452 26124 11508 26126
rect 11676 25618 11732 25620
rect 11676 25566 11678 25618
rect 11678 25566 11730 25618
rect 11730 25566 11732 25618
rect 11676 25564 11732 25566
rect 11788 25506 11844 25508
rect 11788 25454 11790 25506
rect 11790 25454 11842 25506
rect 11842 25454 11844 25506
rect 11788 25452 11844 25454
rect 11340 25228 11396 25284
rect 11004 23772 11060 23828
rect 11228 23938 11284 23940
rect 11228 23886 11230 23938
rect 11230 23886 11282 23938
rect 11282 23886 11284 23938
rect 11228 23884 11284 23886
rect 10892 23266 10948 23268
rect 10892 23214 10894 23266
rect 10894 23214 10946 23266
rect 10946 23214 10948 23266
rect 10892 23212 10948 23214
rect 10780 23100 10836 23156
rect 9660 18396 9716 18452
rect 8316 15314 8372 15316
rect 8316 15262 8318 15314
rect 8318 15262 8370 15314
rect 8370 15262 8372 15314
rect 8316 15260 8372 15262
rect 8652 15148 8708 15204
rect 8092 14588 8148 14644
rect 8092 12908 8148 12964
rect 6188 12402 6244 12404
rect 6188 12350 6190 12402
rect 6190 12350 6242 12402
rect 6242 12350 6244 12402
rect 6188 12348 6244 12350
rect 8092 12348 8148 12404
rect 6972 12124 7028 12180
rect 6636 11394 6692 11396
rect 6636 11342 6638 11394
rect 6638 11342 6690 11394
rect 6690 11342 6692 11394
rect 6636 11340 6692 11342
rect 7644 9100 7700 9156
rect 5516 6412 5572 6468
rect 5628 6524 5684 6580
rect 6748 8370 6804 8372
rect 6748 8318 6750 8370
rect 6750 8318 6802 8370
rect 6802 8318 6804 8370
rect 6748 8316 6804 8318
rect 7196 8034 7252 8036
rect 7196 7982 7198 8034
rect 7198 7982 7250 8034
rect 7250 7982 7252 8034
rect 7196 7980 7252 7982
rect 5068 5180 5124 5236
rect 4284 4060 4340 4116
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 5964 5234 6020 5236
rect 5964 5182 5966 5234
rect 5966 5182 6018 5234
rect 6018 5182 6020 5234
rect 5964 5180 6020 5182
rect 6636 6076 6692 6132
rect 7196 6524 7252 6580
rect 8428 12178 8484 12180
rect 8428 12126 8430 12178
rect 8430 12126 8482 12178
rect 8482 12126 8484 12178
rect 8428 12124 8484 12126
rect 8540 11116 8596 11172
rect 8764 14700 8820 14756
rect 10220 22482 10276 22484
rect 10220 22430 10222 22482
rect 10222 22430 10274 22482
rect 10274 22430 10276 22482
rect 10220 22428 10276 22430
rect 10332 20860 10388 20916
rect 10332 20524 10388 20580
rect 10108 19292 10164 19348
rect 10220 19068 10276 19124
rect 10220 18620 10276 18676
rect 10220 17106 10276 17108
rect 10220 17054 10222 17106
rect 10222 17054 10274 17106
rect 10274 17054 10276 17106
rect 10220 17052 10276 17054
rect 10668 21586 10724 21588
rect 10668 21534 10670 21586
rect 10670 21534 10722 21586
rect 10722 21534 10724 21586
rect 10668 21532 10724 21534
rect 10892 20748 10948 20804
rect 11228 23324 11284 23380
rect 11228 23154 11284 23156
rect 11228 23102 11230 23154
rect 11230 23102 11282 23154
rect 11282 23102 11284 23154
rect 11228 23100 11284 23102
rect 11116 22258 11172 22260
rect 11116 22206 11118 22258
rect 11118 22206 11170 22258
rect 11170 22206 11172 22258
rect 11116 22204 11172 22206
rect 10668 20018 10724 20020
rect 10668 19966 10670 20018
rect 10670 19966 10722 20018
rect 10722 19966 10724 20018
rect 10668 19964 10724 19966
rect 11116 20188 11172 20244
rect 11004 19346 11060 19348
rect 11004 19294 11006 19346
rect 11006 19294 11058 19346
rect 11058 19294 11060 19346
rect 11004 19292 11060 19294
rect 10556 18674 10612 18676
rect 10556 18622 10558 18674
rect 10558 18622 10610 18674
rect 10610 18622 10612 18674
rect 10556 18620 10612 18622
rect 11564 25282 11620 25284
rect 11564 25230 11566 25282
rect 11566 25230 11618 25282
rect 11618 25230 11620 25282
rect 11564 25228 11620 25230
rect 11452 24332 11508 24388
rect 11676 23826 11732 23828
rect 11676 23774 11678 23826
rect 11678 23774 11730 23826
rect 11730 23774 11732 23826
rect 11676 23772 11732 23774
rect 11900 23660 11956 23716
rect 11788 23378 11844 23380
rect 11788 23326 11790 23378
rect 11790 23326 11842 23378
rect 11842 23326 11844 23378
rect 11788 23324 11844 23326
rect 11452 22204 11508 22260
rect 11676 21420 11732 21476
rect 11788 20802 11844 20804
rect 11788 20750 11790 20802
rect 11790 20750 11842 20802
rect 11842 20750 11844 20802
rect 11788 20748 11844 20750
rect 11564 19964 11620 20020
rect 11564 19068 11620 19124
rect 11340 18956 11396 19012
rect 12124 26348 12180 26404
rect 12236 25788 12292 25844
rect 12460 27244 12516 27300
rect 12460 26796 12516 26852
rect 12348 25452 12404 25508
rect 12460 26124 12516 26180
rect 12236 24892 12292 24948
rect 12572 25788 12628 25844
rect 12572 25506 12628 25508
rect 12572 25454 12574 25506
rect 12574 25454 12626 25506
rect 12626 25454 12628 25506
rect 12572 25452 12628 25454
rect 12460 23772 12516 23828
rect 12012 22204 12068 22260
rect 12236 22146 12292 22148
rect 12236 22094 12238 22146
rect 12238 22094 12290 22146
rect 12290 22094 12292 22146
rect 12236 22092 12292 22094
rect 12348 21980 12404 22036
rect 12124 21308 12180 21364
rect 12236 21586 12292 21588
rect 12236 21534 12238 21586
rect 12238 21534 12290 21586
rect 12290 21534 12292 21586
rect 12236 21532 12292 21534
rect 12124 21084 12180 21140
rect 12348 21084 12404 21140
rect 12236 20748 12292 20804
rect 12348 20860 12404 20916
rect 12012 20018 12068 20020
rect 12012 19966 12014 20018
rect 12014 19966 12066 20018
rect 12066 19966 12068 20018
rect 12012 19964 12068 19966
rect 11900 19292 11956 19348
rect 11788 19068 11844 19124
rect 10220 15932 10276 15988
rect 9660 15202 9716 15204
rect 9660 15150 9662 15202
rect 9662 15150 9714 15202
rect 9714 15150 9716 15202
rect 9660 15148 9716 15150
rect 9996 15148 10052 15204
rect 9548 14588 9604 14644
rect 8764 12908 8820 12964
rect 8764 12738 8820 12740
rect 8764 12686 8766 12738
rect 8766 12686 8818 12738
rect 8818 12686 8820 12738
rect 8764 12684 8820 12686
rect 10108 13692 10164 13748
rect 10108 13356 10164 13412
rect 9884 12850 9940 12852
rect 9884 12798 9886 12850
rect 9886 12798 9938 12850
rect 9938 12798 9940 12850
rect 9884 12796 9940 12798
rect 11228 16882 11284 16884
rect 11228 16830 11230 16882
rect 11230 16830 11282 16882
rect 11282 16830 11284 16882
rect 11228 16828 11284 16830
rect 10556 13746 10612 13748
rect 10556 13694 10558 13746
rect 10558 13694 10610 13746
rect 10610 13694 10612 13746
rect 10556 13692 10612 13694
rect 10892 13692 10948 13748
rect 10444 12962 10500 12964
rect 10444 12910 10446 12962
rect 10446 12910 10498 12962
rect 10498 12910 10500 12962
rect 10444 12908 10500 12910
rect 10108 12684 10164 12740
rect 12796 26796 12852 26852
rect 13020 26796 13076 26852
rect 12908 26178 12964 26180
rect 12908 26126 12910 26178
rect 12910 26126 12962 26178
rect 12962 26126 12964 26178
rect 12908 26124 12964 26126
rect 13244 28140 13300 28196
rect 13356 27580 13412 27636
rect 13132 25452 13188 25508
rect 13244 26348 13300 26404
rect 14252 33180 14308 33236
rect 14812 38444 14868 38500
rect 14924 38332 14980 38388
rect 15148 38220 15204 38276
rect 15036 38162 15092 38164
rect 15036 38110 15038 38162
rect 15038 38110 15090 38162
rect 15090 38110 15092 38162
rect 15036 38108 15092 38110
rect 15036 37938 15092 37940
rect 15036 37886 15038 37938
rect 15038 37886 15090 37938
rect 15090 37886 15092 37938
rect 15036 37884 15092 37886
rect 14924 36204 14980 36260
rect 15036 35922 15092 35924
rect 15036 35870 15038 35922
rect 15038 35870 15090 35922
rect 15090 35870 15092 35922
rect 15036 35868 15092 35870
rect 15372 37548 15428 37604
rect 15260 37212 15316 37268
rect 15260 36988 15316 37044
rect 15260 36428 15316 36484
rect 14812 34130 14868 34132
rect 14812 34078 14814 34130
rect 14814 34078 14866 34130
rect 14866 34078 14868 34130
rect 14812 34076 14868 34078
rect 15148 34690 15204 34692
rect 15148 34638 15150 34690
rect 15150 34638 15202 34690
rect 15202 34638 15204 34690
rect 15148 34636 15204 34638
rect 15596 37212 15652 37268
rect 16044 40348 16100 40404
rect 17388 46060 17444 46116
rect 17388 45890 17444 45892
rect 17388 45838 17390 45890
rect 17390 45838 17442 45890
rect 17442 45838 17444 45890
rect 17388 45836 17444 45838
rect 16940 45612 16996 45668
rect 16828 43820 16884 43876
rect 16380 43538 16436 43540
rect 16380 43486 16382 43538
rect 16382 43486 16434 43538
rect 16434 43486 16436 43538
rect 16380 43484 16436 43486
rect 16380 43260 16436 43316
rect 16492 42588 16548 42644
rect 16380 42476 16436 42532
rect 16604 42476 16660 42532
rect 16380 40962 16436 40964
rect 16380 40910 16382 40962
rect 16382 40910 16434 40962
rect 16434 40910 16436 40962
rect 16380 40908 16436 40910
rect 16604 40796 16660 40852
rect 16268 40460 16324 40516
rect 16380 40684 16436 40740
rect 16492 40514 16548 40516
rect 16492 40462 16494 40514
rect 16494 40462 16546 40514
rect 16546 40462 16548 40514
rect 16492 40460 16548 40462
rect 17276 44098 17332 44100
rect 17276 44046 17278 44098
rect 17278 44046 17330 44098
rect 17330 44046 17332 44098
rect 17276 44044 17332 44046
rect 18172 49420 18228 49476
rect 18172 48914 18228 48916
rect 18172 48862 18174 48914
rect 18174 48862 18226 48914
rect 18226 48862 18228 48914
rect 18172 48860 18228 48862
rect 17948 48300 18004 48356
rect 19292 52556 19348 52612
rect 18844 51772 18900 51828
rect 19404 52444 19460 52500
rect 18956 51266 19012 51268
rect 18956 51214 18958 51266
rect 18958 51214 19010 51266
rect 19010 51214 19012 51266
rect 18956 51212 19012 51214
rect 18732 50370 18788 50372
rect 18732 50318 18734 50370
rect 18734 50318 18786 50370
rect 18786 50318 18788 50370
rect 18732 50316 18788 50318
rect 18620 50204 18676 50260
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 20300 54572 20356 54628
rect 20636 55410 20692 55412
rect 20636 55358 20638 55410
rect 20638 55358 20690 55410
rect 20690 55358 20692 55410
rect 20636 55356 20692 55358
rect 20748 54684 20804 54740
rect 20524 53900 20580 53956
rect 20412 53842 20468 53844
rect 20412 53790 20414 53842
rect 20414 53790 20466 53842
rect 20466 53790 20468 53842
rect 20412 53788 20468 53790
rect 20636 52892 20692 52948
rect 20636 52444 20692 52500
rect 20524 52332 20580 52388
rect 20636 52108 20692 52164
rect 20300 51884 20356 51940
rect 19740 51266 19796 51268
rect 19740 51214 19742 51266
rect 19742 51214 19794 51266
rect 19794 51214 19796 51266
rect 19740 51212 19796 51214
rect 20076 50876 20132 50932
rect 19068 50092 19124 50148
rect 19292 50092 19348 50148
rect 18508 49810 18564 49812
rect 18508 49758 18510 49810
rect 18510 49758 18562 49810
rect 18562 49758 18564 49810
rect 18508 49756 18564 49758
rect 18396 49420 18452 49476
rect 18396 49138 18452 49140
rect 18396 49086 18398 49138
rect 18398 49086 18450 49138
rect 18450 49086 18452 49138
rect 18396 49084 18452 49086
rect 18396 48524 18452 48580
rect 18284 48300 18340 48356
rect 17836 48130 17892 48132
rect 17836 48078 17838 48130
rect 17838 48078 17890 48130
rect 17890 48078 17892 48130
rect 17836 48076 17892 48078
rect 17612 47570 17668 47572
rect 17612 47518 17614 47570
rect 17614 47518 17666 47570
rect 17666 47518 17668 47570
rect 17612 47516 17668 47518
rect 18508 48188 18564 48244
rect 19404 49980 19460 50036
rect 19180 48412 19236 48468
rect 18172 47964 18228 48020
rect 17948 47292 18004 47348
rect 17724 47180 17780 47236
rect 17836 46508 17892 46564
rect 18060 46956 18116 47012
rect 17948 46284 18004 46340
rect 17836 46060 17892 46116
rect 18956 47516 19012 47572
rect 18620 46396 18676 46452
rect 18508 46172 18564 46228
rect 17948 44380 18004 44436
rect 17500 44044 17556 44100
rect 17052 43820 17108 43876
rect 17276 43260 17332 43316
rect 16940 41580 16996 41636
rect 16940 41074 16996 41076
rect 16940 41022 16942 41074
rect 16942 41022 16994 41074
rect 16994 41022 16996 41074
rect 16940 41020 16996 41022
rect 16940 40684 16996 40740
rect 16828 39788 16884 39844
rect 16156 39340 16212 39396
rect 16268 39676 16324 39732
rect 16268 39004 16324 39060
rect 16044 38444 16100 38500
rect 16156 38780 16212 38836
rect 15932 38220 15988 38276
rect 15484 36876 15540 36932
rect 15484 35084 15540 35140
rect 14924 32956 14980 33012
rect 14364 32674 14420 32676
rect 14364 32622 14366 32674
rect 14366 32622 14418 32674
rect 14418 32622 14420 32674
rect 14364 32620 14420 32622
rect 13692 30716 13748 30772
rect 13580 29932 13636 29988
rect 13468 26236 13524 26292
rect 13580 29372 13636 29428
rect 13020 24050 13076 24052
rect 13020 23998 13022 24050
rect 13022 23998 13074 24050
rect 13074 23998 13076 24050
rect 13020 23996 13076 23998
rect 13468 23436 13524 23492
rect 13804 29426 13860 29428
rect 13804 29374 13806 29426
rect 13806 29374 13858 29426
rect 13858 29374 13860 29426
rect 13804 29372 13860 29374
rect 13692 29260 13748 29316
rect 13692 28476 13748 28532
rect 13804 28364 13860 28420
rect 13692 28140 13748 28196
rect 14700 32172 14756 32228
rect 14924 32060 14980 32116
rect 14700 31724 14756 31780
rect 14588 31666 14644 31668
rect 14588 31614 14590 31666
rect 14590 31614 14642 31666
rect 14642 31614 14644 31666
rect 14588 31612 14644 31614
rect 14140 30268 14196 30324
rect 14028 29932 14084 29988
rect 14140 29596 14196 29652
rect 14252 29708 14308 29764
rect 14364 29426 14420 29428
rect 14364 29374 14366 29426
rect 14366 29374 14418 29426
rect 14418 29374 14420 29426
rect 14364 29372 14420 29374
rect 14364 29202 14420 29204
rect 14364 29150 14366 29202
rect 14366 29150 14418 29202
rect 14418 29150 14420 29202
rect 14364 29148 14420 29150
rect 14140 28642 14196 28644
rect 14140 28590 14142 28642
rect 14142 28590 14194 28642
rect 14194 28590 14196 28642
rect 14140 28588 14196 28590
rect 14252 28252 14308 28308
rect 14588 28700 14644 28756
rect 14812 30828 14868 30884
rect 15148 33964 15204 34020
rect 15148 31948 15204 32004
rect 15260 33292 15316 33348
rect 15260 31724 15316 31780
rect 15148 31500 15204 31556
rect 15148 30994 15204 30996
rect 15148 30942 15150 30994
rect 15150 30942 15202 30994
rect 15202 30942 15204 30994
rect 15148 30940 15204 30942
rect 15484 31948 15540 32004
rect 16380 39228 16436 39284
rect 16716 39618 16772 39620
rect 16716 39566 16718 39618
rect 16718 39566 16770 39618
rect 16770 39566 16772 39618
rect 16716 39564 16772 39566
rect 18060 43820 18116 43876
rect 18284 45330 18340 45332
rect 18284 45278 18286 45330
rect 18286 45278 18338 45330
rect 18338 45278 18340 45330
rect 18284 45276 18340 45278
rect 18620 44828 18676 44884
rect 17948 43484 18004 43540
rect 17612 42924 17668 42980
rect 17388 42642 17444 42644
rect 17388 42590 17390 42642
rect 17390 42590 17442 42642
rect 17442 42590 17444 42642
rect 17388 42588 17444 42590
rect 17276 41804 17332 41860
rect 17948 42476 18004 42532
rect 18284 44322 18340 44324
rect 18284 44270 18286 44322
rect 18286 44270 18338 44322
rect 18338 44270 18340 44322
rect 18284 44268 18340 44270
rect 18172 42364 18228 42420
rect 17836 42028 17892 42084
rect 17612 41804 17668 41860
rect 17836 41858 17892 41860
rect 17836 41806 17838 41858
rect 17838 41806 17890 41858
rect 17890 41806 17892 41858
rect 17836 41804 17892 41806
rect 17724 41356 17780 41412
rect 17388 40684 17444 40740
rect 17836 40908 17892 40964
rect 17164 39676 17220 39732
rect 16716 39058 16772 39060
rect 16716 39006 16718 39058
rect 16718 39006 16770 39058
rect 16770 39006 16772 39058
rect 16716 39004 16772 39006
rect 17164 39506 17220 39508
rect 17164 39454 17166 39506
rect 17166 39454 17218 39506
rect 17218 39454 17220 39506
rect 17164 39452 17220 39454
rect 17612 39788 17668 39844
rect 18060 41132 18116 41188
rect 18172 40572 18228 40628
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 19852 49922 19908 49924
rect 19852 49870 19854 49922
rect 19854 49870 19906 49922
rect 19906 49870 19908 49922
rect 19852 49868 19908 49870
rect 19292 47346 19348 47348
rect 19292 47294 19294 47346
rect 19294 47294 19346 47346
rect 19346 47294 19348 47346
rect 19292 47292 19348 47294
rect 19292 44716 19348 44772
rect 19292 44380 19348 44436
rect 20076 49026 20132 49028
rect 20076 48974 20078 49026
rect 20078 48974 20130 49026
rect 20130 48974 20132 49026
rect 20076 48972 20132 48974
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 19628 48076 19684 48132
rect 19852 47516 19908 47572
rect 20076 47570 20132 47572
rect 20076 47518 20078 47570
rect 20078 47518 20130 47570
rect 20130 47518 20132 47570
rect 20076 47516 20132 47518
rect 20524 49084 20580 49140
rect 20412 47740 20468 47796
rect 20972 56588 21028 56644
rect 20972 55020 21028 55076
rect 20860 52892 20916 52948
rect 20860 52162 20916 52164
rect 20860 52110 20862 52162
rect 20862 52110 20914 52162
rect 20914 52110 20916 52162
rect 20860 52108 20916 52110
rect 21868 58828 21924 58884
rect 21756 58716 21812 58772
rect 21868 58156 21924 58212
rect 21420 56082 21476 56084
rect 21420 56030 21422 56082
rect 21422 56030 21474 56082
rect 21474 56030 21476 56082
rect 21420 56028 21476 56030
rect 21308 55692 21364 55748
rect 21196 54124 21252 54180
rect 21644 55020 21700 55076
rect 21084 51996 21140 52052
rect 21196 53004 21252 53060
rect 20860 50092 20916 50148
rect 20972 50316 21028 50372
rect 20748 49810 20804 49812
rect 20748 49758 20750 49810
rect 20750 49758 20802 49810
rect 20802 49758 20804 49810
rect 20748 49756 20804 49758
rect 20860 49138 20916 49140
rect 20860 49086 20862 49138
rect 20862 49086 20914 49138
rect 20914 49086 20916 49138
rect 20860 49084 20916 49086
rect 20860 48354 20916 48356
rect 20860 48302 20862 48354
rect 20862 48302 20914 48354
rect 20914 48302 20916 48354
rect 20860 48300 20916 48302
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 20188 47068 20244 47124
rect 19628 45948 19684 46004
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 20412 46956 20468 47012
rect 20412 46562 20468 46564
rect 20412 46510 20414 46562
rect 20414 46510 20466 46562
rect 20466 46510 20468 46562
rect 20412 46508 20468 46510
rect 20300 45836 20356 45892
rect 20636 47068 20692 47124
rect 20860 47516 20916 47572
rect 20412 45388 20468 45444
rect 20188 45106 20244 45108
rect 20188 45054 20190 45106
rect 20190 45054 20242 45106
rect 20242 45054 20244 45106
rect 20188 45052 20244 45054
rect 19068 44322 19124 44324
rect 19068 44270 19070 44322
rect 19070 44270 19122 44322
rect 19122 44270 19124 44322
rect 19068 44268 19124 44270
rect 19180 44210 19236 44212
rect 19180 44158 19182 44210
rect 19182 44158 19234 44210
rect 19234 44158 19236 44210
rect 19180 44156 19236 44158
rect 18844 43596 18900 43652
rect 18956 43538 19012 43540
rect 18956 43486 18958 43538
rect 18958 43486 19010 43538
rect 19010 43486 19012 43538
rect 18956 43484 19012 43486
rect 18732 43372 18788 43428
rect 18396 42866 18452 42868
rect 18396 42814 18398 42866
rect 18398 42814 18450 42866
rect 18450 42814 18452 42866
rect 18396 42812 18452 42814
rect 18732 42700 18788 42756
rect 19404 43596 19460 43652
rect 19516 44044 19572 44100
rect 19180 43260 19236 43316
rect 19068 42924 19124 42980
rect 19740 44380 19796 44436
rect 20300 44380 20356 44436
rect 20524 45276 20580 45332
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 19628 43484 19684 43540
rect 20412 43708 20468 43764
rect 20300 43484 20356 43540
rect 19628 42924 19684 42980
rect 19516 42812 19572 42868
rect 18620 42530 18676 42532
rect 18620 42478 18622 42530
rect 18622 42478 18674 42530
rect 18674 42478 18676 42530
rect 18620 42476 18676 42478
rect 18284 40348 18340 40404
rect 18396 42364 18452 42420
rect 17948 40124 18004 40180
rect 19180 42364 19236 42420
rect 18620 41298 18676 41300
rect 18620 41246 18622 41298
rect 18622 41246 18674 41298
rect 18674 41246 18676 41298
rect 18620 41244 18676 41246
rect 18732 41020 18788 41076
rect 18732 40796 18788 40852
rect 18508 40402 18564 40404
rect 18508 40350 18510 40402
rect 18510 40350 18562 40402
rect 18562 40350 18564 40402
rect 18508 40348 18564 40350
rect 19964 42642 20020 42644
rect 19964 42590 19966 42642
rect 19966 42590 20018 42642
rect 20018 42590 20020 42642
rect 19964 42588 20020 42590
rect 19516 42364 19572 42420
rect 19628 42476 19684 42532
rect 20524 43260 20580 43316
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20412 42364 20468 42420
rect 20044 42308 20100 42310
rect 20860 45388 20916 45444
rect 21308 49980 21364 50036
rect 21420 53116 21476 53172
rect 21084 48466 21140 48468
rect 21084 48414 21086 48466
rect 21086 48414 21138 48466
rect 21138 48414 21140 48466
rect 21084 48412 21140 48414
rect 21644 53004 21700 53060
rect 22092 58604 22148 58660
rect 22316 58716 22372 58772
rect 22092 56924 22148 56980
rect 21980 56140 22036 56196
rect 22316 56754 22372 56756
rect 22316 56702 22318 56754
rect 22318 56702 22370 56754
rect 22370 56702 22372 56754
rect 22316 56700 22372 56702
rect 23324 59612 23380 59668
rect 23548 59500 23604 59556
rect 24108 59612 24164 59668
rect 22988 59164 23044 59220
rect 23884 59218 23940 59220
rect 23884 59166 23886 59218
rect 23886 59166 23938 59218
rect 23938 59166 23940 59218
rect 23884 59164 23940 59166
rect 23548 58716 23604 58772
rect 22764 58604 22820 58660
rect 22540 57708 22596 57764
rect 22092 56028 22148 56084
rect 22540 56364 22596 56420
rect 22428 56082 22484 56084
rect 22428 56030 22430 56082
rect 22430 56030 22482 56082
rect 22482 56030 22484 56082
rect 22428 56028 22484 56030
rect 21980 55916 22036 55972
rect 21868 55244 21924 55300
rect 22204 54908 22260 54964
rect 22092 54348 22148 54404
rect 21756 52556 21812 52612
rect 21980 53058 22036 53060
rect 21980 53006 21982 53058
rect 21982 53006 22034 53058
rect 22034 53006 22036 53058
rect 21980 53004 22036 53006
rect 22316 53788 22372 53844
rect 22764 57090 22820 57092
rect 22764 57038 22766 57090
rect 22766 57038 22818 57090
rect 22818 57038 22820 57090
rect 22764 57036 22820 57038
rect 23436 57484 23492 57540
rect 23772 57484 23828 57540
rect 24556 59500 24612 59556
rect 24668 59724 24724 59780
rect 24556 58546 24612 58548
rect 24556 58494 24558 58546
rect 24558 58494 24610 58546
rect 24610 58494 24612 58546
rect 24556 58492 24612 58494
rect 24444 58322 24500 58324
rect 24444 58270 24446 58322
rect 24446 58270 24498 58322
rect 24498 58270 24500 58322
rect 24444 58268 24500 58270
rect 24108 57538 24164 57540
rect 24108 57486 24110 57538
rect 24110 57486 24162 57538
rect 24162 57486 24164 57538
rect 24108 57484 24164 57486
rect 23660 57036 23716 57092
rect 23996 57090 24052 57092
rect 23996 57038 23998 57090
rect 23998 57038 24050 57090
rect 24050 57038 24052 57090
rect 23996 57036 24052 57038
rect 25228 59612 25284 59668
rect 24892 59500 24948 59556
rect 24780 58434 24836 58436
rect 24780 58382 24782 58434
rect 24782 58382 24834 58434
rect 24834 58382 24836 58434
rect 24780 58380 24836 58382
rect 24108 56924 24164 56980
rect 24780 57484 24836 57540
rect 23772 56866 23828 56868
rect 23772 56814 23774 56866
rect 23774 56814 23826 56866
rect 23826 56814 23828 56866
rect 23772 56812 23828 56814
rect 23324 56364 23380 56420
rect 24108 56364 24164 56420
rect 23212 56252 23268 56308
rect 23660 56306 23716 56308
rect 23660 56254 23662 56306
rect 23662 56254 23714 56306
rect 23714 56254 23716 56306
rect 23660 56252 23716 56254
rect 23324 55580 23380 55636
rect 23884 55580 23940 55636
rect 23996 55804 24052 55860
rect 23772 55468 23828 55524
rect 22428 53730 22484 53732
rect 22428 53678 22430 53730
rect 22430 53678 22482 53730
rect 22482 53678 22484 53730
rect 22428 53676 22484 53678
rect 22540 55244 22596 55300
rect 22540 53116 22596 53172
rect 22652 54908 22708 54964
rect 22764 54738 22820 54740
rect 22764 54686 22766 54738
rect 22766 54686 22818 54738
rect 22818 54686 22820 54738
rect 22764 54684 22820 54686
rect 23324 53900 23380 53956
rect 23212 53676 23268 53732
rect 22988 53618 23044 53620
rect 22988 53566 22990 53618
rect 22990 53566 23042 53618
rect 23042 53566 23044 53618
rect 22988 53564 23044 53566
rect 23436 53564 23492 53620
rect 22652 53506 22708 53508
rect 22652 53454 22654 53506
rect 22654 53454 22706 53506
rect 22706 53454 22708 53506
rect 22652 53452 22708 53454
rect 22540 52946 22596 52948
rect 22540 52894 22542 52946
rect 22542 52894 22594 52946
rect 22594 52894 22596 52946
rect 22540 52892 22596 52894
rect 22428 52834 22484 52836
rect 22428 52782 22430 52834
rect 22430 52782 22482 52834
rect 22482 52782 22484 52834
rect 22428 52780 22484 52782
rect 22204 52556 22260 52612
rect 22876 53506 22932 53508
rect 22876 53454 22878 53506
rect 22878 53454 22930 53506
rect 22930 53454 22932 53506
rect 22876 53452 22932 53454
rect 22764 53228 22820 53284
rect 22876 53116 22932 53172
rect 21868 52108 21924 52164
rect 21756 51996 21812 52052
rect 21532 51660 21588 51716
rect 21644 51884 21700 51940
rect 21532 51436 21588 51492
rect 21644 49868 21700 49924
rect 21644 48914 21700 48916
rect 21644 48862 21646 48914
rect 21646 48862 21698 48914
rect 21698 48862 21700 48914
rect 21644 48860 21700 48862
rect 22540 52162 22596 52164
rect 22540 52110 22542 52162
rect 22542 52110 22594 52162
rect 22594 52110 22596 52162
rect 22540 52108 22596 52110
rect 22316 50706 22372 50708
rect 22316 50654 22318 50706
rect 22318 50654 22370 50706
rect 22370 50654 22372 50706
rect 22316 50652 22372 50654
rect 22204 50204 22260 50260
rect 22092 49868 22148 49924
rect 21980 49026 22036 49028
rect 21980 48974 21982 49026
rect 21982 48974 22034 49026
rect 22034 48974 22036 49026
rect 21980 48972 22036 48974
rect 21420 48412 21476 48468
rect 21308 48300 21364 48356
rect 21532 47068 21588 47124
rect 21308 45724 21364 45780
rect 21644 46396 21700 46452
rect 21532 45666 21588 45668
rect 21532 45614 21534 45666
rect 21534 45614 21586 45666
rect 21586 45614 21588 45666
rect 21532 45612 21588 45614
rect 21644 45218 21700 45220
rect 21644 45166 21646 45218
rect 21646 45166 21698 45218
rect 21698 45166 21700 45218
rect 21644 45164 21700 45166
rect 21308 44716 21364 44772
rect 20748 44268 20804 44324
rect 19740 41804 19796 41860
rect 19292 41692 19348 41748
rect 19180 41244 19236 41300
rect 19292 41468 19348 41524
rect 19068 41132 19124 41188
rect 19404 41356 19460 41412
rect 21196 43596 21252 43652
rect 21084 43426 21140 43428
rect 21084 43374 21086 43426
rect 21086 43374 21138 43426
rect 21138 43374 21140 43426
rect 21084 43372 21140 43374
rect 21308 43484 21364 43540
rect 21420 43260 21476 43316
rect 20860 42252 20916 42308
rect 21084 41970 21140 41972
rect 21084 41918 21086 41970
rect 21086 41918 21138 41970
rect 21138 41918 21140 41970
rect 21084 41916 21140 41918
rect 20524 41746 20580 41748
rect 20524 41694 20526 41746
rect 20526 41694 20578 41746
rect 20578 41694 20580 41746
rect 20524 41692 20580 41694
rect 19628 40796 19684 40852
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 18844 40348 18900 40404
rect 18620 40290 18676 40292
rect 18620 40238 18622 40290
rect 18622 40238 18674 40290
rect 18674 40238 18676 40290
rect 18620 40236 18676 40238
rect 16940 39228 16996 39284
rect 16044 35810 16100 35812
rect 16044 35758 16046 35810
rect 16046 35758 16098 35810
rect 16098 35758 16100 35810
rect 16044 35756 16100 35758
rect 16044 35026 16100 35028
rect 16044 34974 16046 35026
rect 16046 34974 16098 35026
rect 16098 34974 16100 35026
rect 16044 34972 16100 34974
rect 15932 34860 15988 34916
rect 15820 34130 15876 34132
rect 15820 34078 15822 34130
rect 15822 34078 15874 34130
rect 15874 34078 15876 34130
rect 15820 34076 15876 34078
rect 16044 33964 16100 34020
rect 16604 38722 16660 38724
rect 16604 38670 16606 38722
rect 16606 38670 16658 38722
rect 16658 38670 16660 38722
rect 16604 38668 16660 38670
rect 16940 38556 16996 38612
rect 17276 39228 17332 39284
rect 16604 37324 16660 37380
rect 16492 37266 16548 37268
rect 16492 37214 16494 37266
rect 16494 37214 16546 37266
rect 16546 37214 16548 37266
rect 16492 37212 16548 37214
rect 16380 36764 16436 36820
rect 17164 37212 17220 37268
rect 16828 37042 16884 37044
rect 16828 36990 16830 37042
rect 16830 36990 16882 37042
rect 16882 36990 16884 37042
rect 16828 36988 16884 36990
rect 16716 36876 16772 36932
rect 16716 36706 16772 36708
rect 16716 36654 16718 36706
rect 16718 36654 16770 36706
rect 16770 36654 16772 36706
rect 16716 36652 16772 36654
rect 16268 35810 16324 35812
rect 16268 35758 16270 35810
rect 16270 35758 16322 35810
rect 16322 35758 16324 35810
rect 16268 35756 16324 35758
rect 16156 33516 16212 33572
rect 15820 32786 15876 32788
rect 15820 32734 15822 32786
rect 15822 32734 15874 32786
rect 15874 32734 15876 32786
rect 15820 32732 15876 32734
rect 16044 33180 16100 33236
rect 15820 32396 15876 32452
rect 15484 31388 15540 31444
rect 15596 31500 15652 31556
rect 15036 29820 15092 29876
rect 15708 30268 15764 30324
rect 16268 33404 16324 33460
rect 16716 36428 16772 36484
rect 16828 36370 16884 36372
rect 16828 36318 16830 36370
rect 16830 36318 16882 36370
rect 16882 36318 16884 36370
rect 16828 36316 16884 36318
rect 17052 36316 17108 36372
rect 16940 35922 16996 35924
rect 16940 35870 16942 35922
rect 16942 35870 16994 35922
rect 16994 35870 16996 35922
rect 16940 35868 16996 35870
rect 16492 35756 16548 35812
rect 16604 35698 16660 35700
rect 16604 35646 16606 35698
rect 16606 35646 16658 35698
rect 16658 35646 16660 35698
rect 16604 35644 16660 35646
rect 16828 35698 16884 35700
rect 16828 35646 16830 35698
rect 16830 35646 16882 35698
rect 16882 35646 16884 35698
rect 16828 35644 16884 35646
rect 16940 35420 16996 35476
rect 16604 35084 16660 35140
rect 16380 33292 16436 33348
rect 16268 32508 16324 32564
rect 16156 32396 16212 32452
rect 16492 32450 16548 32452
rect 16492 32398 16494 32450
rect 16494 32398 16546 32450
rect 16546 32398 16548 32450
rect 16492 32396 16548 32398
rect 16492 31106 16548 31108
rect 16492 31054 16494 31106
rect 16494 31054 16546 31106
rect 16546 31054 16548 31106
rect 16492 31052 16548 31054
rect 16156 30940 16212 30996
rect 16044 30828 16100 30884
rect 16828 34188 16884 34244
rect 17052 34748 17108 34804
rect 17164 35868 17220 35924
rect 16940 33740 16996 33796
rect 16716 33068 16772 33124
rect 17052 33068 17108 33124
rect 16828 32284 16884 32340
rect 16828 31948 16884 32004
rect 17052 31724 17108 31780
rect 16716 31052 16772 31108
rect 16380 30210 16436 30212
rect 16380 30158 16382 30210
rect 16382 30158 16434 30210
rect 16434 30158 16436 30210
rect 16380 30156 16436 30158
rect 14924 29372 14980 29428
rect 14812 29148 14868 29204
rect 15260 29372 15316 29428
rect 14924 28754 14980 28756
rect 14924 28702 14926 28754
rect 14926 28702 14978 28754
rect 14978 28702 14980 28754
rect 14924 28700 14980 28702
rect 15036 28588 15092 28644
rect 14924 28530 14980 28532
rect 14924 28478 14926 28530
rect 14926 28478 14978 28530
rect 14978 28478 14980 28530
rect 14924 28476 14980 28478
rect 14028 26572 14084 26628
rect 14140 26348 14196 26404
rect 13916 26124 13972 26180
rect 14476 26460 14532 26516
rect 14588 27580 14644 27636
rect 14252 26012 14308 26068
rect 14028 25452 14084 25508
rect 14700 27132 14756 27188
rect 14140 24892 14196 24948
rect 14700 26572 14756 26628
rect 13580 23324 13636 23380
rect 13916 23548 13972 23604
rect 12796 23266 12852 23268
rect 12796 23214 12798 23266
rect 12798 23214 12850 23266
rect 12850 23214 12852 23266
rect 12796 23212 12852 23214
rect 13804 23212 13860 23268
rect 12684 22092 12740 22148
rect 13020 23100 13076 23156
rect 12572 21308 12628 21364
rect 12572 20018 12628 20020
rect 12572 19966 12574 20018
rect 12574 19966 12626 20018
rect 12626 19966 12628 20018
rect 12572 19964 12628 19966
rect 12572 19346 12628 19348
rect 12572 19294 12574 19346
rect 12574 19294 12626 19346
rect 12626 19294 12628 19346
rect 12572 19292 12628 19294
rect 12124 19068 12180 19124
rect 12124 18508 12180 18564
rect 12572 18450 12628 18452
rect 12572 18398 12574 18450
rect 12574 18398 12626 18450
rect 12626 18398 12628 18450
rect 12572 18396 12628 18398
rect 12012 17052 12068 17108
rect 12236 16828 12292 16884
rect 14028 24444 14084 24500
rect 13132 22092 13188 22148
rect 13132 21196 13188 21252
rect 13468 20972 13524 21028
rect 13692 21308 13748 21364
rect 13916 20972 13972 21028
rect 13356 20524 13412 20580
rect 12908 19010 12964 19012
rect 12908 18958 12910 19010
rect 12910 18958 12962 19010
rect 12962 18958 12964 19010
rect 12908 18956 12964 18958
rect 13020 16210 13076 16212
rect 13020 16158 13022 16210
rect 13022 16158 13074 16210
rect 13074 16158 13076 16210
rect 13020 16156 13076 16158
rect 11788 15314 11844 15316
rect 11788 15262 11790 15314
rect 11790 15262 11842 15314
rect 11842 15262 11844 15314
rect 11788 15260 11844 15262
rect 11564 15148 11620 15204
rect 13356 18396 13412 18452
rect 13468 18508 13524 18564
rect 13468 15820 13524 15876
rect 11228 13746 11284 13748
rect 11228 13694 11230 13746
rect 11230 13694 11282 13746
rect 11282 13694 11284 13746
rect 11228 13692 11284 13694
rect 11116 13356 11172 13412
rect 11900 13356 11956 13412
rect 11340 13132 11396 13188
rect 11116 12908 11172 12964
rect 11340 12908 11396 12964
rect 11900 12962 11956 12964
rect 11900 12910 11902 12962
rect 11902 12910 11954 12962
rect 11954 12910 11956 12962
rect 11900 12908 11956 12910
rect 12460 12908 12516 12964
rect 12908 12962 12964 12964
rect 12908 12910 12910 12962
rect 12910 12910 12962 12962
rect 12962 12910 12964 12962
rect 12908 12908 12964 12910
rect 13804 20578 13860 20580
rect 13804 20526 13806 20578
rect 13806 20526 13858 20578
rect 13858 20526 13860 20578
rect 13804 20524 13860 20526
rect 14140 20860 14196 20916
rect 13916 18956 13972 19012
rect 14028 19852 14084 19908
rect 14924 24892 14980 24948
rect 14476 23378 14532 23380
rect 14476 23326 14478 23378
rect 14478 23326 14530 23378
rect 14530 23326 14532 23378
rect 14476 23324 14532 23326
rect 15148 27916 15204 27972
rect 15372 27692 15428 27748
rect 15372 27074 15428 27076
rect 15372 27022 15374 27074
rect 15374 27022 15426 27074
rect 15426 27022 15428 27074
rect 15372 27020 15428 27022
rect 15148 23436 15204 23492
rect 15148 22146 15204 22148
rect 15148 22094 15150 22146
rect 15150 22094 15202 22146
rect 15202 22094 15204 22146
rect 15148 22092 15204 22094
rect 14364 19346 14420 19348
rect 14364 19294 14366 19346
rect 14366 19294 14418 19346
rect 14418 19294 14420 19346
rect 14364 19292 14420 19294
rect 13692 16156 13748 16212
rect 13916 16828 13972 16884
rect 14028 16716 14084 16772
rect 14028 15874 14084 15876
rect 14028 15822 14030 15874
rect 14030 15822 14082 15874
rect 14082 15822 14084 15874
rect 14028 15820 14084 15822
rect 14700 19010 14756 19012
rect 14700 18958 14702 19010
rect 14702 18958 14754 19010
rect 14754 18958 14756 19010
rect 14700 18956 14756 18958
rect 15372 25506 15428 25508
rect 15372 25454 15374 25506
rect 15374 25454 15426 25506
rect 15426 25454 15428 25506
rect 15372 25452 15428 25454
rect 16604 30322 16660 30324
rect 16604 30270 16606 30322
rect 16606 30270 16658 30322
rect 16658 30270 16660 30322
rect 16604 30268 16660 30270
rect 15820 29484 15876 29540
rect 15708 28082 15764 28084
rect 15708 28030 15710 28082
rect 15710 28030 15762 28082
rect 15762 28030 15764 28082
rect 15708 28028 15764 28030
rect 16604 29596 16660 29652
rect 16156 29426 16212 29428
rect 16156 29374 16158 29426
rect 16158 29374 16210 29426
rect 16210 29374 16212 29426
rect 16156 29372 16212 29374
rect 16156 28252 16212 28308
rect 15596 27580 15652 27636
rect 15932 28028 15988 28084
rect 15820 26962 15876 26964
rect 15820 26910 15822 26962
rect 15822 26910 15874 26962
rect 15874 26910 15876 26962
rect 15820 26908 15876 26910
rect 15708 26796 15764 26852
rect 15708 24946 15764 24948
rect 15708 24894 15710 24946
rect 15710 24894 15762 24946
rect 15762 24894 15764 24946
rect 15708 24892 15764 24894
rect 15484 23324 15540 23380
rect 15596 23436 15652 23492
rect 15484 23154 15540 23156
rect 15484 23102 15486 23154
rect 15486 23102 15538 23154
rect 15538 23102 15540 23154
rect 15484 23100 15540 23102
rect 15820 21756 15876 21812
rect 15596 21586 15652 21588
rect 15596 21534 15598 21586
rect 15598 21534 15650 21586
rect 15650 21534 15652 21586
rect 15596 21532 15652 21534
rect 15820 21420 15876 21476
rect 15260 20860 15316 20916
rect 16380 28028 16436 28084
rect 16156 27916 16212 27972
rect 16604 28364 16660 28420
rect 16492 27916 16548 27972
rect 16268 27692 16324 27748
rect 16828 30940 16884 30996
rect 16940 30380 16996 30436
rect 17388 38780 17444 38836
rect 17388 36988 17444 37044
rect 17724 39228 17780 39284
rect 18844 40012 18900 40068
rect 17948 39452 18004 39508
rect 18060 39788 18116 39844
rect 17836 38780 17892 38836
rect 17612 38556 17668 38612
rect 17836 37660 17892 37716
rect 17724 37100 17780 37156
rect 18620 39730 18676 39732
rect 18620 39678 18622 39730
rect 18622 39678 18674 39730
rect 18674 39678 18676 39730
rect 18620 39676 18676 39678
rect 18284 39618 18340 39620
rect 18284 39566 18286 39618
rect 18286 39566 18338 39618
rect 18338 39566 18340 39618
rect 18284 39564 18340 39566
rect 18732 39564 18788 39620
rect 18620 39452 18676 39508
rect 18284 39228 18340 39284
rect 18396 39340 18452 39396
rect 18284 38946 18340 38948
rect 18284 38894 18286 38946
rect 18286 38894 18338 38946
rect 18338 38894 18340 38946
rect 18284 38892 18340 38894
rect 18172 38722 18228 38724
rect 18172 38670 18174 38722
rect 18174 38670 18226 38722
rect 18226 38670 18228 38722
rect 18172 38668 18228 38670
rect 18172 38162 18228 38164
rect 18172 38110 18174 38162
rect 18174 38110 18226 38162
rect 18226 38110 18228 38162
rect 18172 38108 18228 38110
rect 18172 37548 18228 37604
rect 18844 39394 18900 39396
rect 18844 39342 18846 39394
rect 18846 39342 18898 39394
rect 18898 39342 18900 39394
rect 18844 39340 18900 39342
rect 19068 39340 19124 39396
rect 18508 39004 18564 39060
rect 18060 36876 18116 36932
rect 18508 37212 18564 37268
rect 17836 36594 17892 36596
rect 17836 36542 17838 36594
rect 17838 36542 17890 36594
rect 17890 36542 17892 36594
rect 17836 36540 17892 36542
rect 17836 35980 17892 36036
rect 17612 35644 17668 35700
rect 17500 35196 17556 35252
rect 17500 34860 17556 34916
rect 17276 34636 17332 34692
rect 18284 36540 18340 36596
rect 18172 36482 18228 36484
rect 18172 36430 18174 36482
rect 18174 36430 18226 36482
rect 18226 36430 18228 36482
rect 18172 36428 18228 36430
rect 18060 36092 18116 36148
rect 17948 34972 18004 35028
rect 17948 34690 18004 34692
rect 17948 34638 17950 34690
rect 17950 34638 18002 34690
rect 18002 34638 18004 34690
rect 17948 34636 18004 34638
rect 17276 31724 17332 31780
rect 17388 33964 17444 34020
rect 17612 33516 17668 33572
rect 17836 33964 17892 34020
rect 17836 33346 17892 33348
rect 17836 33294 17838 33346
rect 17838 33294 17890 33346
rect 17890 33294 17892 33346
rect 17836 33292 17892 33294
rect 18284 35868 18340 35924
rect 18284 35698 18340 35700
rect 18284 35646 18286 35698
rect 18286 35646 18338 35698
rect 18338 35646 18340 35698
rect 18284 35644 18340 35646
rect 18620 36764 18676 36820
rect 18508 35084 18564 35140
rect 18396 35026 18452 35028
rect 18396 34974 18398 35026
rect 18398 34974 18450 35026
rect 18450 34974 18452 35026
rect 18396 34972 18452 34974
rect 18620 34412 18676 34468
rect 18956 39004 19012 39060
rect 19180 38892 19236 38948
rect 19628 40626 19684 40628
rect 19628 40574 19630 40626
rect 19630 40574 19682 40626
rect 19682 40574 19684 40626
rect 19628 40572 19684 40574
rect 20748 41244 20804 41300
rect 20412 41020 20468 41076
rect 19404 39676 19460 39732
rect 20188 40124 20244 40180
rect 19964 39730 20020 39732
rect 19964 39678 19966 39730
rect 19966 39678 20018 39730
rect 20018 39678 20020 39730
rect 19964 39676 20020 39678
rect 19852 39506 19908 39508
rect 19852 39454 19854 39506
rect 19854 39454 19906 39506
rect 19906 39454 19908 39506
rect 19852 39452 19908 39454
rect 20076 39394 20132 39396
rect 20076 39342 20078 39394
rect 20078 39342 20130 39394
rect 20130 39342 20132 39394
rect 20076 39340 20132 39342
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 20188 38892 20244 38948
rect 19404 38834 19460 38836
rect 19404 38782 19406 38834
rect 19406 38782 19458 38834
rect 19458 38782 19460 38834
rect 19404 38780 19460 38782
rect 19292 38556 19348 38612
rect 19628 38556 19684 38612
rect 19404 38444 19460 38500
rect 18844 37212 18900 37268
rect 19068 37826 19124 37828
rect 19068 37774 19070 37826
rect 19070 37774 19122 37826
rect 19122 37774 19124 37826
rect 19068 37772 19124 37774
rect 19292 37212 19348 37268
rect 18956 36764 19012 36820
rect 19180 36876 19236 36932
rect 19516 36988 19572 37044
rect 18956 35980 19012 36036
rect 19068 35644 19124 35700
rect 19404 35922 19460 35924
rect 19404 35870 19406 35922
rect 19406 35870 19458 35922
rect 19458 35870 19460 35922
rect 19404 35868 19460 35870
rect 19180 35420 19236 35476
rect 18396 33740 18452 33796
rect 18844 35196 18900 35252
rect 18732 34018 18788 34020
rect 18732 33966 18734 34018
rect 18734 33966 18786 34018
rect 18786 33966 18788 34018
rect 18732 33964 18788 33966
rect 17724 33122 17780 33124
rect 17724 33070 17726 33122
rect 17726 33070 17778 33122
rect 17778 33070 17780 33122
rect 17724 33068 17780 33070
rect 17388 32732 17444 32788
rect 17948 32450 18004 32452
rect 17948 32398 17950 32450
rect 17950 32398 18002 32450
rect 18002 32398 18004 32450
rect 17948 32396 18004 32398
rect 17724 32338 17780 32340
rect 17724 32286 17726 32338
rect 17726 32286 17778 32338
rect 17778 32286 17780 32338
rect 17724 32284 17780 32286
rect 18396 33346 18452 33348
rect 18396 33294 18398 33346
rect 18398 33294 18450 33346
rect 18450 33294 18452 33346
rect 18396 33292 18452 33294
rect 18620 33234 18676 33236
rect 18620 33182 18622 33234
rect 18622 33182 18674 33234
rect 18674 33182 18676 33234
rect 18620 33180 18676 33182
rect 18284 33068 18340 33124
rect 18060 32284 18116 32340
rect 17724 31890 17780 31892
rect 17724 31838 17726 31890
rect 17726 31838 17778 31890
rect 17778 31838 17780 31890
rect 17724 31836 17780 31838
rect 17388 31500 17444 31556
rect 18396 32786 18452 32788
rect 18396 32734 18398 32786
rect 18398 32734 18450 32786
rect 18450 32734 18452 32786
rect 18396 32732 18452 32734
rect 18620 32284 18676 32340
rect 19292 35084 19348 35140
rect 18956 34914 19012 34916
rect 18956 34862 18958 34914
rect 18958 34862 19010 34914
rect 19010 34862 19012 34914
rect 18956 34860 19012 34862
rect 19180 34802 19236 34804
rect 19180 34750 19182 34802
rect 19182 34750 19234 34802
rect 19234 34750 19236 34802
rect 19180 34748 19236 34750
rect 19404 34690 19460 34692
rect 19404 34638 19406 34690
rect 19406 34638 19458 34690
rect 19458 34638 19460 34690
rect 19404 34636 19460 34638
rect 19964 37996 20020 38052
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 19964 37490 20020 37492
rect 19964 37438 19966 37490
rect 19966 37438 20018 37490
rect 20018 37438 20020 37490
rect 19964 37436 20020 37438
rect 20636 40908 20692 40964
rect 20524 40460 20580 40516
rect 21980 47570 22036 47572
rect 21980 47518 21982 47570
rect 21982 47518 22034 47570
rect 22034 47518 22036 47570
rect 21980 47516 22036 47518
rect 21756 44492 21812 44548
rect 21868 47180 21924 47236
rect 22092 46620 22148 46676
rect 22204 49756 22260 49812
rect 22092 44604 22148 44660
rect 22316 47516 22372 47572
rect 22540 49980 22596 50036
rect 22540 48860 22596 48916
rect 22988 53004 23044 53060
rect 23324 52780 23380 52836
rect 23100 52556 23156 52612
rect 23436 52668 23492 52724
rect 24220 55074 24276 55076
rect 24220 55022 24222 55074
rect 24222 55022 24274 55074
rect 24274 55022 24276 55074
rect 24220 55020 24276 55022
rect 24444 54738 24500 54740
rect 24444 54686 24446 54738
rect 24446 54686 24498 54738
rect 24498 54686 24500 54738
rect 24444 54684 24500 54686
rect 24220 53730 24276 53732
rect 24220 53678 24222 53730
rect 24222 53678 24274 53730
rect 24274 53678 24276 53730
rect 24220 53676 24276 53678
rect 23772 53452 23828 53508
rect 23324 52108 23380 52164
rect 23100 51938 23156 51940
rect 23100 51886 23102 51938
rect 23102 51886 23154 51938
rect 23154 51886 23156 51938
rect 23100 51884 23156 51886
rect 23212 51772 23268 51828
rect 23660 52892 23716 52948
rect 23884 52834 23940 52836
rect 23884 52782 23886 52834
rect 23886 52782 23938 52834
rect 23938 52782 23940 52834
rect 23884 52780 23940 52782
rect 23996 52668 24052 52724
rect 24220 52892 24276 52948
rect 23772 52162 23828 52164
rect 23772 52110 23774 52162
rect 23774 52110 23826 52162
rect 23826 52110 23828 52162
rect 23772 52108 23828 52110
rect 22876 50652 22932 50708
rect 23212 50876 23268 50932
rect 22876 50428 22932 50484
rect 22764 49980 22820 50036
rect 23100 50204 23156 50260
rect 23100 49084 23156 49140
rect 22652 48300 22708 48356
rect 23100 48636 23156 48692
rect 22764 47740 22820 47796
rect 22540 46396 22596 46452
rect 22540 45500 22596 45556
rect 23324 50316 23380 50372
rect 22988 48300 23044 48356
rect 23772 50540 23828 50596
rect 24668 55298 24724 55300
rect 24668 55246 24670 55298
rect 24670 55246 24722 55298
rect 24722 55246 24724 55298
rect 24668 55244 24724 55246
rect 25004 56924 25060 56980
rect 25116 56866 25172 56868
rect 25116 56814 25118 56866
rect 25118 56814 25170 56866
rect 25170 56814 25172 56866
rect 25116 56812 25172 56814
rect 25228 56642 25284 56644
rect 25228 56590 25230 56642
rect 25230 56590 25282 56642
rect 25282 56590 25284 56642
rect 25228 56588 25284 56590
rect 25004 55804 25060 55860
rect 25004 54402 25060 54404
rect 25004 54350 25006 54402
rect 25006 54350 25058 54402
rect 25058 54350 25060 54402
rect 25004 54348 25060 54350
rect 24668 53452 24724 53508
rect 24668 53058 24724 53060
rect 24668 53006 24670 53058
rect 24670 53006 24722 53058
rect 24722 53006 24724 53058
rect 24668 53004 24724 53006
rect 24332 51996 24388 52052
rect 23660 48748 23716 48804
rect 23436 48466 23492 48468
rect 23436 48414 23438 48466
rect 23438 48414 23490 48466
rect 23490 48414 23492 48466
rect 23436 48412 23492 48414
rect 23324 48354 23380 48356
rect 23324 48302 23326 48354
rect 23326 48302 23378 48354
rect 23378 48302 23380 48354
rect 23324 48300 23380 48302
rect 23548 47964 23604 48020
rect 23324 47458 23380 47460
rect 23324 47406 23326 47458
rect 23326 47406 23378 47458
rect 23378 47406 23380 47458
rect 23324 47404 23380 47406
rect 23772 47404 23828 47460
rect 24108 51772 24164 51828
rect 24108 50316 24164 50372
rect 24444 51938 24500 51940
rect 24444 51886 24446 51938
rect 24446 51886 24498 51938
rect 24498 51886 24500 51938
rect 24444 51884 24500 51886
rect 24892 53116 24948 53172
rect 25004 52780 25060 52836
rect 24780 51772 24836 51828
rect 35196 60394 35252 60396
rect 35196 60342 35198 60394
rect 35198 60342 35250 60394
rect 35250 60342 35252 60394
rect 35196 60340 35252 60342
rect 35300 60394 35356 60396
rect 35300 60342 35302 60394
rect 35302 60342 35354 60394
rect 35354 60342 35356 60394
rect 35300 60340 35356 60342
rect 35404 60394 35460 60396
rect 35404 60342 35406 60394
rect 35406 60342 35458 60394
rect 35458 60342 35460 60394
rect 35404 60340 35460 60342
rect 30156 60060 30212 60116
rect 31052 60114 31108 60116
rect 31052 60062 31054 60114
rect 31054 60062 31106 60114
rect 31106 60062 31108 60114
rect 31052 60060 31108 60062
rect 50204 60060 50260 60116
rect 51100 60114 51156 60116
rect 51100 60062 51102 60114
rect 51102 60062 51154 60114
rect 51154 60062 51156 60114
rect 51100 60060 51156 60062
rect 25676 59612 25732 59668
rect 26684 59276 26740 59332
rect 29820 59778 29876 59780
rect 29820 59726 29822 59778
rect 29822 59726 29874 59778
rect 29874 59726 29876 59778
rect 29820 59724 29876 59726
rect 30380 59724 30436 59780
rect 26908 59276 26964 59332
rect 28028 59218 28084 59220
rect 28028 59166 28030 59218
rect 28030 59166 28082 59218
rect 28082 59166 28084 59218
rect 28028 59164 28084 59166
rect 27244 58716 27300 58772
rect 27692 58828 27748 58884
rect 26796 58492 26852 58548
rect 26908 58604 26964 58660
rect 25900 58434 25956 58436
rect 25900 58382 25902 58434
rect 25902 58382 25954 58434
rect 25954 58382 25956 58434
rect 25900 58380 25956 58382
rect 26460 58380 26516 58436
rect 25452 58268 25508 58324
rect 26348 58322 26404 58324
rect 26348 58270 26350 58322
rect 26350 58270 26402 58322
rect 26402 58270 26404 58322
rect 26348 58268 26404 58270
rect 25564 57538 25620 57540
rect 25564 57486 25566 57538
rect 25566 57486 25618 57538
rect 25618 57486 25620 57538
rect 25564 57484 25620 57486
rect 25788 56978 25844 56980
rect 25788 56926 25790 56978
rect 25790 56926 25842 56978
rect 25842 56926 25844 56978
rect 25788 56924 25844 56926
rect 25452 55580 25508 55636
rect 25564 55410 25620 55412
rect 25564 55358 25566 55410
rect 25566 55358 25618 55410
rect 25618 55358 25620 55410
rect 25564 55356 25620 55358
rect 26348 57148 26404 57204
rect 26124 57036 26180 57092
rect 26236 55356 26292 55412
rect 25452 54908 25508 54964
rect 24220 48860 24276 48916
rect 24108 48748 24164 48804
rect 23996 48636 24052 48692
rect 24556 51378 24612 51380
rect 24556 51326 24558 51378
rect 24558 51326 24610 51378
rect 24610 51326 24612 51378
rect 24556 51324 24612 51326
rect 25340 52332 25396 52388
rect 25004 51548 25060 51604
rect 25228 51938 25284 51940
rect 25228 51886 25230 51938
rect 25230 51886 25282 51938
rect 25282 51886 25284 51938
rect 25228 51884 25284 51886
rect 24780 49698 24836 49700
rect 24780 49646 24782 49698
rect 24782 49646 24834 49698
rect 24834 49646 24836 49698
rect 24780 49644 24836 49646
rect 24668 49196 24724 49252
rect 25116 50482 25172 50484
rect 25116 50430 25118 50482
rect 25118 50430 25170 50482
rect 25170 50430 25172 50482
rect 25116 50428 25172 50430
rect 25004 49196 25060 49252
rect 24444 48130 24500 48132
rect 24444 48078 24446 48130
rect 24446 48078 24498 48130
rect 24498 48078 24500 48130
rect 24444 48076 24500 48078
rect 26012 55020 26068 55076
rect 25564 54124 25620 54180
rect 25676 53340 25732 53396
rect 26012 53788 26068 53844
rect 25676 53004 25732 53060
rect 25900 53340 25956 53396
rect 25676 52108 25732 52164
rect 27356 58546 27412 58548
rect 27356 58494 27358 58546
rect 27358 58494 27410 58546
rect 27410 58494 27412 58546
rect 27356 58492 27412 58494
rect 27468 58322 27524 58324
rect 27468 58270 27470 58322
rect 27470 58270 27522 58322
rect 27522 58270 27524 58322
rect 27468 58268 27524 58270
rect 27132 57932 27188 57988
rect 26572 57036 26628 57092
rect 27020 56476 27076 56532
rect 26460 55298 26516 55300
rect 26460 55246 26462 55298
rect 26462 55246 26514 55298
rect 26514 55246 26516 55298
rect 26460 55244 26516 55246
rect 26572 55020 26628 55076
rect 28700 59164 28756 59220
rect 28140 58492 28196 58548
rect 27804 58268 27860 58324
rect 27916 57932 27972 57988
rect 28364 58716 28420 58772
rect 28588 58604 28644 58660
rect 28812 58322 28868 58324
rect 28812 58270 28814 58322
rect 28814 58270 28866 58322
rect 28866 58270 28868 58322
rect 28812 58268 28868 58270
rect 29148 58268 29204 58324
rect 28588 57932 28644 57988
rect 28700 57650 28756 57652
rect 28700 57598 28702 57650
rect 28702 57598 28754 57650
rect 28754 57598 28756 57650
rect 28700 57596 28756 57598
rect 29932 58940 29988 58996
rect 29484 58156 29540 58212
rect 27916 57260 27972 57316
rect 27356 55970 27412 55972
rect 27356 55918 27358 55970
rect 27358 55918 27410 55970
rect 27410 55918 27412 55970
rect 27356 55916 27412 55918
rect 27020 55692 27076 55748
rect 27132 55298 27188 55300
rect 27132 55246 27134 55298
rect 27134 55246 27186 55298
rect 27186 55246 27188 55298
rect 27132 55244 27188 55246
rect 27244 54514 27300 54516
rect 27244 54462 27246 54514
rect 27246 54462 27298 54514
rect 27298 54462 27300 54514
rect 27244 54460 27300 54462
rect 26348 52892 26404 52948
rect 27468 53676 27524 53732
rect 27692 55132 27748 55188
rect 26124 52556 26180 52612
rect 26348 52332 26404 52388
rect 24780 48076 24836 48132
rect 24892 48860 24948 48916
rect 24668 47852 24724 47908
rect 23772 47234 23828 47236
rect 23772 47182 23774 47234
rect 23774 47182 23826 47234
rect 23826 47182 23828 47234
rect 23772 47180 23828 47182
rect 22876 45388 22932 45444
rect 23324 46732 23380 46788
rect 22652 45052 22708 45108
rect 22092 44322 22148 44324
rect 22092 44270 22094 44322
rect 22094 44270 22146 44322
rect 22146 44270 22148 44322
rect 22092 44268 22148 44270
rect 21756 44156 21812 44212
rect 21644 43538 21700 43540
rect 21644 43486 21646 43538
rect 21646 43486 21698 43538
rect 21698 43486 21700 43538
rect 21644 43484 21700 43486
rect 21644 42140 21700 42196
rect 22204 44156 22260 44212
rect 22316 44268 22372 44324
rect 21980 43484 22036 43540
rect 22204 42754 22260 42756
rect 22204 42702 22206 42754
rect 22206 42702 22258 42754
rect 22258 42702 22260 42754
rect 22204 42700 22260 42702
rect 21980 42140 22036 42196
rect 22092 42588 22148 42644
rect 20748 40684 20804 40740
rect 21420 41020 21476 41076
rect 21308 40626 21364 40628
rect 21308 40574 21310 40626
rect 21310 40574 21362 40626
rect 21362 40574 21364 40626
rect 21308 40572 21364 40574
rect 20972 40460 21028 40516
rect 21196 40402 21252 40404
rect 21196 40350 21198 40402
rect 21198 40350 21250 40402
rect 21250 40350 21252 40402
rect 21196 40348 21252 40350
rect 21532 40348 21588 40404
rect 21868 42028 21924 42084
rect 21756 41132 21812 41188
rect 21756 40684 21812 40740
rect 20972 39618 21028 39620
rect 20972 39566 20974 39618
rect 20974 39566 21026 39618
rect 21026 39566 21028 39618
rect 20972 39564 21028 39566
rect 20524 37042 20580 37044
rect 20524 36990 20526 37042
rect 20526 36990 20578 37042
rect 20578 36990 20580 37042
rect 20524 36988 20580 36990
rect 19964 36370 20020 36372
rect 19964 36318 19966 36370
rect 19966 36318 20018 36370
rect 20018 36318 20020 36370
rect 19964 36316 20020 36318
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 20076 35532 20132 35588
rect 20076 35084 20132 35140
rect 19628 34860 19684 34916
rect 19180 33964 19236 34020
rect 19068 33516 19124 33572
rect 18956 33068 19012 33124
rect 18956 32732 19012 32788
rect 20076 34914 20132 34916
rect 20076 34862 20078 34914
rect 20078 34862 20130 34914
rect 20130 34862 20132 34914
rect 20076 34860 20132 34862
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19740 34018 19796 34020
rect 19740 33966 19742 34018
rect 19742 33966 19794 34018
rect 19794 33966 19796 34018
rect 19740 33964 19796 33966
rect 20748 38668 20804 38724
rect 20748 37324 20804 37380
rect 20748 36652 20804 36708
rect 20972 37378 21028 37380
rect 20972 37326 20974 37378
rect 20974 37326 21026 37378
rect 21026 37326 21028 37378
rect 20972 37324 21028 37326
rect 21084 37266 21140 37268
rect 21084 37214 21086 37266
rect 21086 37214 21138 37266
rect 21138 37214 21140 37266
rect 21084 37212 21140 37214
rect 21980 40572 22036 40628
rect 22316 42588 22372 42644
rect 22428 42700 22484 42756
rect 22316 42140 22372 42196
rect 22428 41970 22484 41972
rect 22428 41918 22430 41970
rect 22430 41918 22482 41970
rect 22482 41918 22484 41970
rect 22428 41916 22484 41918
rect 22316 40796 22372 40852
rect 22204 40626 22260 40628
rect 22204 40574 22206 40626
rect 22206 40574 22258 40626
rect 22258 40574 22260 40626
rect 22204 40572 22260 40574
rect 22316 40460 22372 40516
rect 21868 40348 21924 40404
rect 21532 38834 21588 38836
rect 21532 38782 21534 38834
rect 21534 38782 21586 38834
rect 21586 38782 21588 38834
rect 21532 38780 21588 38782
rect 21644 37324 21700 37380
rect 21868 38050 21924 38052
rect 21868 37998 21870 38050
rect 21870 37998 21922 38050
rect 21922 37998 21924 38050
rect 21868 37996 21924 37998
rect 21868 37490 21924 37492
rect 21868 37438 21870 37490
rect 21870 37438 21922 37490
rect 21922 37438 21924 37490
rect 21868 37436 21924 37438
rect 22092 37490 22148 37492
rect 22092 37438 22094 37490
rect 22094 37438 22146 37490
rect 22146 37438 22148 37490
rect 22092 37436 22148 37438
rect 22764 43708 22820 43764
rect 22764 42812 22820 42868
rect 23548 46674 23604 46676
rect 23548 46622 23550 46674
rect 23550 46622 23602 46674
rect 23602 46622 23604 46674
rect 23548 46620 23604 46622
rect 23212 45666 23268 45668
rect 23212 45614 23214 45666
rect 23214 45614 23266 45666
rect 23266 45614 23268 45666
rect 23212 45612 23268 45614
rect 23100 45500 23156 45556
rect 22988 44268 23044 44324
rect 23772 46786 23828 46788
rect 23772 46734 23774 46786
rect 23774 46734 23826 46786
rect 23826 46734 23828 46786
rect 23772 46732 23828 46734
rect 24556 47346 24612 47348
rect 24556 47294 24558 47346
rect 24558 47294 24610 47346
rect 24610 47294 24612 47346
rect 24556 47292 24612 47294
rect 24332 47234 24388 47236
rect 24332 47182 24334 47234
rect 24334 47182 24386 47234
rect 24386 47182 24388 47234
rect 24332 47180 24388 47182
rect 24444 46620 24500 46676
rect 24220 46396 24276 46452
rect 24220 45778 24276 45780
rect 24220 45726 24222 45778
rect 24222 45726 24274 45778
rect 24274 45726 24276 45778
rect 24220 45724 24276 45726
rect 23996 45388 24052 45444
rect 24332 45388 24388 45444
rect 24668 46060 24724 46116
rect 25228 49026 25284 49028
rect 25228 48974 25230 49026
rect 25230 48974 25282 49026
rect 25282 48974 25284 49026
rect 25228 48972 25284 48974
rect 25116 47404 25172 47460
rect 24892 46732 24948 46788
rect 25228 47180 25284 47236
rect 24780 45948 24836 46004
rect 24892 46396 24948 46452
rect 23660 44828 23716 44884
rect 23772 45106 23828 45108
rect 23772 45054 23774 45106
rect 23774 45054 23826 45106
rect 23826 45054 23828 45106
rect 23772 45052 23828 45054
rect 23212 44156 23268 44212
rect 23100 43148 23156 43204
rect 23100 42642 23156 42644
rect 23100 42590 23102 42642
rect 23102 42590 23154 42642
rect 23154 42590 23156 42642
rect 23100 42588 23156 42590
rect 23548 44098 23604 44100
rect 23548 44046 23550 44098
rect 23550 44046 23602 44098
rect 23602 44046 23604 44098
rect 23548 44044 23604 44046
rect 24220 45106 24276 45108
rect 24220 45054 24222 45106
rect 24222 45054 24274 45106
rect 24274 45054 24276 45106
rect 24220 45052 24276 45054
rect 23884 44940 23940 44996
rect 24332 44828 24388 44884
rect 24220 44604 24276 44660
rect 23884 44098 23940 44100
rect 23884 44046 23886 44098
rect 23886 44046 23938 44098
rect 23938 44046 23940 44098
rect 23884 44044 23940 44046
rect 23772 43932 23828 43988
rect 22876 41468 22932 41524
rect 22876 41020 22932 41076
rect 22652 40514 22708 40516
rect 22652 40462 22654 40514
rect 22654 40462 22706 40514
rect 22706 40462 22708 40514
rect 22652 40460 22708 40462
rect 22876 40348 22932 40404
rect 23436 41580 23492 41636
rect 23212 41298 23268 41300
rect 23212 41246 23214 41298
rect 23214 41246 23266 41298
rect 23266 41246 23268 41298
rect 23212 41244 23268 41246
rect 22988 40012 23044 40068
rect 23100 39116 23156 39172
rect 23100 38892 23156 38948
rect 22988 38668 23044 38724
rect 22876 38444 22932 38500
rect 22652 38162 22708 38164
rect 22652 38110 22654 38162
rect 22654 38110 22706 38162
rect 22706 38110 22708 38162
rect 22652 38108 22708 38110
rect 21980 37266 22036 37268
rect 21980 37214 21982 37266
rect 21982 37214 22034 37266
rect 22034 37214 22036 37266
rect 21980 37212 22036 37214
rect 20860 36258 20916 36260
rect 20860 36206 20862 36258
rect 20862 36206 20914 36258
rect 20914 36206 20916 36258
rect 20860 36204 20916 36206
rect 20412 35980 20468 36036
rect 20300 35922 20356 35924
rect 20300 35870 20302 35922
rect 20302 35870 20354 35922
rect 20354 35870 20356 35922
rect 20300 35868 20356 35870
rect 20636 35868 20692 35924
rect 20524 35698 20580 35700
rect 20524 35646 20526 35698
rect 20526 35646 20578 35698
rect 20578 35646 20580 35698
rect 20524 35644 20580 35646
rect 20412 35586 20468 35588
rect 20412 35534 20414 35586
rect 20414 35534 20466 35586
rect 20466 35534 20468 35586
rect 20412 35532 20468 35534
rect 20524 35026 20580 35028
rect 20524 34974 20526 35026
rect 20526 34974 20578 35026
rect 20578 34974 20580 35026
rect 20524 34972 20580 34974
rect 20300 34748 20356 34804
rect 19404 32956 19460 33012
rect 19404 32396 19460 32452
rect 19516 33852 19572 33908
rect 18844 31948 18900 32004
rect 18732 31778 18788 31780
rect 18732 31726 18734 31778
rect 18734 31726 18786 31778
rect 18786 31726 18788 31778
rect 18732 31724 18788 31726
rect 18172 31612 18228 31668
rect 18060 31388 18116 31444
rect 17276 31276 17332 31332
rect 16716 27804 16772 27860
rect 17388 31164 17444 31220
rect 17276 30210 17332 30212
rect 17276 30158 17278 30210
rect 17278 30158 17330 30210
rect 17330 30158 17332 30210
rect 17276 30156 17332 30158
rect 17052 29484 17108 29540
rect 16492 26066 16548 26068
rect 16492 26014 16494 26066
rect 16494 26014 16546 26066
rect 16546 26014 16548 26066
rect 16492 26012 16548 26014
rect 16268 25116 16324 25172
rect 16156 23884 16212 23940
rect 16044 23660 16100 23716
rect 15596 19964 15652 20020
rect 15260 19628 15316 19684
rect 14924 17052 14980 17108
rect 17164 29820 17220 29876
rect 16940 29148 16996 29204
rect 16940 28588 16996 28644
rect 17836 31218 17892 31220
rect 17836 31166 17838 31218
rect 17838 31166 17890 31218
rect 17890 31166 17892 31218
rect 17836 31164 17892 31166
rect 19068 31890 19124 31892
rect 19068 31838 19070 31890
rect 19070 31838 19122 31890
rect 19122 31838 19124 31890
rect 19068 31836 19124 31838
rect 19068 31164 19124 31220
rect 19180 32060 19236 32116
rect 18396 30492 18452 30548
rect 18172 30380 18228 30436
rect 17724 29820 17780 29876
rect 17500 29596 17556 29652
rect 17500 28812 17556 28868
rect 18172 29708 18228 29764
rect 19068 30380 19124 30436
rect 18172 29538 18228 29540
rect 18172 29486 18174 29538
rect 18174 29486 18226 29538
rect 18226 29486 18228 29538
rect 18172 29484 18228 29486
rect 18284 28812 18340 28868
rect 17836 28700 17892 28756
rect 18172 28588 18228 28644
rect 16940 26908 16996 26964
rect 16604 24946 16660 24948
rect 16604 24894 16606 24946
rect 16606 24894 16658 24946
rect 16658 24894 16660 24946
rect 16604 24892 16660 24894
rect 18060 27356 18116 27412
rect 18732 30268 18788 30324
rect 18396 28140 18452 28196
rect 18508 28812 18564 28868
rect 18620 28588 18676 28644
rect 18844 28866 18900 28868
rect 18844 28814 18846 28866
rect 18846 28814 18898 28866
rect 18898 28814 18900 28866
rect 18844 28812 18900 28814
rect 18732 28252 18788 28308
rect 18844 28476 18900 28532
rect 18620 28028 18676 28084
rect 20188 33852 20244 33908
rect 20860 35980 20916 36036
rect 21084 35532 21140 35588
rect 21420 35644 21476 35700
rect 21532 35586 21588 35588
rect 21532 35534 21534 35586
rect 21534 35534 21586 35586
rect 21586 35534 21588 35586
rect 21532 35532 21588 35534
rect 21868 36316 21924 36372
rect 21644 34748 21700 34804
rect 20860 34636 20916 34692
rect 21420 34636 21476 34692
rect 20636 34076 20692 34132
rect 20524 33964 20580 34020
rect 19628 33458 19684 33460
rect 19628 33406 19630 33458
rect 19630 33406 19682 33458
rect 19682 33406 19684 33458
rect 19628 33404 19684 33406
rect 20412 33458 20468 33460
rect 20412 33406 20414 33458
rect 20414 33406 20466 33458
rect 20466 33406 20468 33458
rect 20412 33404 20468 33406
rect 19740 33122 19796 33124
rect 19740 33070 19742 33122
rect 19742 33070 19794 33122
rect 19794 33070 19796 33122
rect 19740 33068 19796 33070
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 20300 32674 20356 32676
rect 20300 32622 20302 32674
rect 20302 32622 20354 32674
rect 20354 32622 20356 32674
rect 20300 32620 20356 32622
rect 19964 32284 20020 32340
rect 20636 32844 20692 32900
rect 20076 31948 20132 32004
rect 20188 32060 20244 32116
rect 19404 31500 19460 31556
rect 19628 31500 19684 31556
rect 19404 30940 19460 30996
rect 19516 31164 19572 31220
rect 19180 30268 19236 30324
rect 19292 30604 19348 30660
rect 19404 30492 19460 30548
rect 19292 29708 19348 29764
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 20524 31948 20580 32004
rect 20412 31666 20468 31668
rect 20412 31614 20414 31666
rect 20414 31614 20466 31666
rect 20466 31614 20468 31666
rect 20412 31612 20468 31614
rect 19628 30604 19684 30660
rect 19628 30434 19684 30436
rect 19628 30382 19630 30434
rect 19630 30382 19682 30434
rect 19682 30382 19684 30434
rect 19628 30380 19684 30382
rect 19740 30044 19796 30100
rect 19852 29932 19908 29988
rect 20300 30716 20356 30772
rect 20412 29986 20468 29988
rect 20412 29934 20414 29986
rect 20414 29934 20466 29986
rect 20466 29934 20468 29986
rect 20412 29932 20468 29934
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19068 28476 19124 28532
rect 18172 26908 18228 26964
rect 19292 27804 19348 27860
rect 18732 26460 18788 26516
rect 18732 26290 18788 26292
rect 18732 26238 18734 26290
rect 18734 26238 18786 26290
rect 18786 26238 18788 26290
rect 18732 26236 18788 26238
rect 18396 25506 18452 25508
rect 18396 25454 18398 25506
rect 18398 25454 18450 25506
rect 18450 25454 18452 25506
rect 18396 25452 18452 25454
rect 17164 24108 17220 24164
rect 17612 23826 17668 23828
rect 17612 23774 17614 23826
rect 17614 23774 17666 23826
rect 17666 23774 17668 23826
rect 17612 23772 17668 23774
rect 16492 23660 16548 23716
rect 16828 23714 16884 23716
rect 16828 23662 16830 23714
rect 16830 23662 16882 23714
rect 16882 23662 16884 23714
rect 16828 23660 16884 23662
rect 18284 24050 18340 24052
rect 18284 23998 18286 24050
rect 18286 23998 18338 24050
rect 18338 23998 18340 24050
rect 18284 23996 18340 23998
rect 18060 23660 18116 23716
rect 17612 23324 17668 23380
rect 16380 22764 16436 22820
rect 16156 20972 16212 21028
rect 16492 20018 16548 20020
rect 16492 19966 16494 20018
rect 16494 19966 16546 20018
rect 16546 19966 16548 20018
rect 16492 19964 16548 19966
rect 16268 19852 16324 19908
rect 15596 18956 15652 19012
rect 16156 18396 16212 18452
rect 15708 18284 15764 18340
rect 14588 16210 14644 16212
rect 14588 16158 14590 16210
rect 14590 16158 14642 16210
rect 14642 16158 14644 16210
rect 14588 16156 14644 16158
rect 15148 16716 15204 16772
rect 16940 23154 16996 23156
rect 16940 23102 16942 23154
rect 16942 23102 16994 23154
rect 16994 23102 16996 23154
rect 16940 23100 16996 23102
rect 17612 22764 17668 22820
rect 16716 20076 16772 20132
rect 16828 21756 16884 21812
rect 16268 17388 16324 17444
rect 16268 16828 16324 16884
rect 16940 21698 16996 21700
rect 16940 21646 16942 21698
rect 16942 21646 16994 21698
rect 16994 21646 16996 21698
rect 16940 21644 16996 21646
rect 17164 21420 17220 21476
rect 17052 19906 17108 19908
rect 17052 19854 17054 19906
rect 17054 19854 17106 19906
rect 17106 19854 17108 19906
rect 17052 19852 17108 19854
rect 18172 23100 18228 23156
rect 17948 22930 18004 22932
rect 17948 22878 17950 22930
rect 17950 22878 18002 22930
rect 18002 22878 18004 22930
rect 17948 22876 18004 22878
rect 17724 21644 17780 21700
rect 17836 21980 17892 22036
rect 18172 21980 18228 22036
rect 18172 21756 18228 21812
rect 17836 21532 17892 21588
rect 17724 20802 17780 20804
rect 17724 20750 17726 20802
rect 17726 20750 17778 20802
rect 17778 20750 17780 20802
rect 17724 20748 17780 20750
rect 18620 25564 18676 25620
rect 18732 24892 18788 24948
rect 19628 29314 19684 29316
rect 19628 29262 19630 29314
rect 19630 29262 19682 29314
rect 19682 29262 19684 29314
rect 19628 29260 19684 29262
rect 20300 29260 20356 29316
rect 20300 28476 20356 28532
rect 18956 26572 19012 26628
rect 19180 26908 19236 26964
rect 19068 26236 19124 26292
rect 18956 25004 19012 25060
rect 18508 23266 18564 23268
rect 18508 23214 18510 23266
rect 18510 23214 18562 23266
rect 18562 23214 18564 23266
rect 18508 23212 18564 23214
rect 19068 23996 19124 24052
rect 18956 23212 19012 23268
rect 18396 22764 18452 22820
rect 18732 22876 18788 22932
rect 18844 21644 18900 21700
rect 18284 21532 18340 21588
rect 18284 21084 18340 21140
rect 18060 20914 18116 20916
rect 18060 20862 18062 20914
rect 18062 20862 18114 20914
rect 18114 20862 18116 20914
rect 18060 20860 18116 20862
rect 18284 20524 18340 20580
rect 18508 19852 18564 19908
rect 18396 19628 18452 19684
rect 17948 18284 18004 18340
rect 16828 17052 16884 17108
rect 18060 17106 18116 17108
rect 18060 17054 18062 17106
rect 18062 17054 18114 17106
rect 18114 17054 18116 17106
rect 18060 17052 18116 17054
rect 17052 16994 17108 16996
rect 17052 16942 17054 16994
rect 17054 16942 17106 16994
rect 17106 16942 17108 16994
rect 17052 16940 17108 16942
rect 17948 16828 18004 16884
rect 15372 15372 15428 15428
rect 15260 15260 15316 15316
rect 14140 14700 14196 14756
rect 14252 13522 14308 13524
rect 14252 13470 14254 13522
rect 14254 13470 14306 13522
rect 14306 13470 14308 13522
rect 14252 13468 14308 13470
rect 13692 13020 13748 13076
rect 13916 13020 13972 13076
rect 10332 11394 10388 11396
rect 10332 11342 10334 11394
rect 10334 11342 10386 11394
rect 10386 11342 10388 11394
rect 10332 11340 10388 11342
rect 11116 11340 11172 11396
rect 9660 10668 9716 10724
rect 8428 9212 8484 9268
rect 8316 9100 8372 9156
rect 9884 9826 9940 9828
rect 9884 9774 9886 9826
rect 9886 9774 9938 9826
rect 9938 9774 9940 9826
rect 9884 9772 9940 9774
rect 9548 8988 9604 9044
rect 8988 8652 9044 8708
rect 7756 8316 7812 8372
rect 7980 8034 8036 8036
rect 7980 7982 7982 8034
rect 7982 7982 8034 8034
rect 8034 7982 8036 8034
rect 7980 7980 8036 7982
rect 8316 7196 8372 7252
rect 8540 7196 8596 7252
rect 7644 6690 7700 6692
rect 7644 6638 7646 6690
rect 7646 6638 7698 6690
rect 7698 6638 7700 6690
rect 7644 6636 7700 6638
rect 8316 6636 8372 6692
rect 7980 6466 8036 6468
rect 7980 6414 7982 6466
rect 7982 6414 8034 6466
rect 8034 6414 8036 6466
rect 7980 6412 8036 6414
rect 7308 6076 7364 6132
rect 5740 3724 5796 3780
rect 9772 8652 9828 8708
rect 10332 10722 10388 10724
rect 10332 10670 10334 10722
rect 10334 10670 10386 10722
rect 10386 10670 10388 10722
rect 10332 10668 10388 10670
rect 11004 9154 11060 9156
rect 11004 9102 11006 9154
rect 11006 9102 11058 9154
rect 11058 9102 11060 9154
rect 11004 9100 11060 9102
rect 10556 9042 10612 9044
rect 10556 8990 10558 9042
rect 10558 8990 10610 9042
rect 10610 8990 10612 9042
rect 10556 8988 10612 8990
rect 8876 6690 8932 6692
rect 8876 6638 8878 6690
rect 8878 6638 8930 6690
rect 8930 6638 8932 6690
rect 8876 6636 8932 6638
rect 9548 6690 9604 6692
rect 9548 6638 9550 6690
rect 9550 6638 9602 6690
rect 9602 6638 9604 6690
rect 9548 6636 9604 6638
rect 8652 6076 8708 6132
rect 9100 6130 9156 6132
rect 9100 6078 9102 6130
rect 9102 6078 9154 6130
rect 9154 6078 9156 6130
rect 9100 6076 9156 6078
rect 8316 5964 8372 6020
rect 8316 5122 8372 5124
rect 8316 5070 8318 5122
rect 8318 5070 8370 5122
rect 8370 5070 8372 5122
rect 8316 5068 8372 5070
rect 9996 6690 10052 6692
rect 9996 6638 9998 6690
rect 9998 6638 10050 6690
rect 10050 6638 10052 6690
rect 9996 6636 10052 6638
rect 10220 6076 10276 6132
rect 9100 4338 9156 4340
rect 9100 4286 9102 4338
rect 9102 4286 9154 4338
rect 9154 4286 9156 4338
rect 9100 4284 9156 4286
rect 7644 4172 7700 4228
rect 6300 3554 6356 3556
rect 6300 3502 6302 3554
rect 6302 3502 6354 3554
rect 6354 3502 6356 3554
rect 6300 3500 6356 3502
rect 10780 5628 10836 5684
rect 9772 4338 9828 4340
rect 9772 4286 9774 4338
rect 9774 4286 9826 4338
rect 9826 4286 9828 4338
rect 9772 4284 9828 4286
rect 10220 4226 10276 4228
rect 10220 4174 10222 4226
rect 10222 4174 10274 4226
rect 10274 4174 10276 4226
rect 10220 4172 10276 4174
rect 13132 11676 13188 11732
rect 12908 11340 12964 11396
rect 12460 9602 12516 9604
rect 12460 9550 12462 9602
rect 12462 9550 12514 9602
rect 12514 9550 12516 9602
rect 12460 9548 12516 9550
rect 13020 10050 13076 10052
rect 13020 9998 13022 10050
rect 13022 9998 13074 10050
rect 13074 9998 13076 10050
rect 13020 9996 13076 9998
rect 13580 10610 13636 10612
rect 13580 10558 13582 10610
rect 13582 10558 13634 10610
rect 13634 10558 13636 10610
rect 13580 10556 13636 10558
rect 13132 9772 13188 9828
rect 13580 8988 13636 9044
rect 13356 8930 13412 8932
rect 13356 8878 13358 8930
rect 13358 8878 13410 8930
rect 13410 8878 13412 8930
rect 13356 8876 13412 8878
rect 13356 7698 13412 7700
rect 13356 7646 13358 7698
rect 13358 7646 13410 7698
rect 13410 7646 13412 7698
rect 13356 7644 13412 7646
rect 13356 7196 13412 7252
rect 14588 13074 14644 13076
rect 14588 13022 14590 13074
rect 14590 13022 14642 13074
rect 14642 13022 14644 13074
rect 14588 13020 14644 13022
rect 14140 12738 14196 12740
rect 14140 12686 14142 12738
rect 14142 12686 14194 12738
rect 14194 12686 14196 12738
rect 14140 12684 14196 12686
rect 14924 12684 14980 12740
rect 16604 15426 16660 15428
rect 16604 15374 16606 15426
rect 16606 15374 16658 15426
rect 16658 15374 16660 15426
rect 16604 15372 16660 15374
rect 17612 15426 17668 15428
rect 17612 15374 17614 15426
rect 17614 15374 17666 15426
rect 17666 15374 17668 15426
rect 17612 15372 17668 15374
rect 16044 14530 16100 14532
rect 16044 14478 16046 14530
rect 16046 14478 16098 14530
rect 16098 14478 16100 14530
rect 16044 14476 16100 14478
rect 18508 18226 18564 18228
rect 18508 18174 18510 18226
rect 18510 18174 18562 18226
rect 18562 18174 18564 18226
rect 18508 18172 18564 18174
rect 18396 16268 18452 16324
rect 18508 17442 18564 17444
rect 18508 17390 18510 17442
rect 18510 17390 18562 17442
rect 18562 17390 18564 17442
rect 18508 17388 18564 17390
rect 18284 16156 18340 16212
rect 18732 20972 18788 21028
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19852 27858 19908 27860
rect 19852 27806 19854 27858
rect 19854 27806 19906 27858
rect 19906 27806 19908 27858
rect 19852 27804 19908 27806
rect 20860 32732 20916 32788
rect 21084 33516 21140 33572
rect 20972 32060 21028 32116
rect 20748 31836 20804 31892
rect 20860 30268 20916 30324
rect 21084 29314 21140 29316
rect 21084 29262 21086 29314
rect 21086 29262 21138 29314
rect 21138 29262 21140 29314
rect 21084 29260 21140 29262
rect 20524 28642 20580 28644
rect 20524 28590 20526 28642
rect 20526 28590 20578 28642
rect 20578 28590 20580 28642
rect 20524 28588 20580 28590
rect 20412 28364 20468 28420
rect 19964 27580 20020 27636
rect 20972 28364 21028 28420
rect 20860 27186 20916 27188
rect 20860 27134 20862 27186
rect 20862 27134 20914 27186
rect 20914 27134 20916 27186
rect 20860 27132 20916 27134
rect 20860 26908 20916 26964
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19964 26460 20020 26516
rect 19404 25004 19460 25060
rect 19628 25676 19684 25732
rect 20076 26178 20132 26180
rect 20076 26126 20078 26178
rect 20078 26126 20130 26178
rect 20130 26126 20132 26178
rect 20076 26124 20132 26126
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20188 25116 20244 25172
rect 20044 25060 20100 25062
rect 19292 24610 19348 24612
rect 19292 24558 19294 24610
rect 19294 24558 19346 24610
rect 19346 24558 19348 24610
rect 19292 24556 19348 24558
rect 20748 25228 20804 25284
rect 20860 26514 20916 26516
rect 20860 26462 20862 26514
rect 20862 26462 20914 26514
rect 20914 26462 20916 26514
rect 20860 26460 20916 26462
rect 20972 26236 21028 26292
rect 20860 24892 20916 24948
rect 20524 24556 20580 24612
rect 19516 24050 19572 24052
rect 19516 23998 19518 24050
rect 19518 23998 19570 24050
rect 19570 23998 19572 24050
rect 19516 23996 19572 23998
rect 19404 23772 19460 23828
rect 20524 23996 20580 24052
rect 19628 23660 19684 23716
rect 20188 23938 20244 23940
rect 20188 23886 20190 23938
rect 20190 23886 20242 23938
rect 20242 23886 20244 23938
rect 20188 23884 20244 23886
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19516 22316 19572 22372
rect 20188 22428 20244 22484
rect 19516 21756 19572 21812
rect 19740 22146 19796 22148
rect 19740 22094 19742 22146
rect 19742 22094 19794 22146
rect 19794 22094 19796 22146
rect 19740 22092 19796 22094
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 20076 21586 20132 21588
rect 20076 21534 20078 21586
rect 20078 21534 20130 21586
rect 20130 21534 20132 21586
rect 20076 21532 20132 21534
rect 20748 23714 20804 23716
rect 20748 23662 20750 23714
rect 20750 23662 20802 23714
rect 20802 23662 20804 23714
rect 20748 23660 20804 23662
rect 20636 23100 20692 23156
rect 20748 22876 20804 22932
rect 20524 21868 20580 21924
rect 20636 22092 20692 22148
rect 20524 21698 20580 21700
rect 20524 21646 20526 21698
rect 20526 21646 20578 21698
rect 20578 21646 20580 21698
rect 20524 21644 20580 21646
rect 20188 20914 20244 20916
rect 20188 20862 20190 20914
rect 20190 20862 20242 20914
rect 20242 20862 20244 20914
rect 20188 20860 20244 20862
rect 18844 16994 18900 16996
rect 18844 16942 18846 16994
rect 18846 16942 18898 16994
rect 18898 16942 18900 16994
rect 18844 16940 18900 16942
rect 18620 16604 18676 16660
rect 19068 19852 19124 19908
rect 19180 20076 19236 20132
rect 19068 19628 19124 19684
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 20188 20188 20244 20244
rect 19292 19628 19348 19684
rect 19404 19852 19460 19908
rect 19180 18338 19236 18340
rect 19180 18286 19182 18338
rect 19182 18286 19234 18338
rect 19234 18286 19236 18338
rect 19180 18284 19236 18286
rect 20860 22370 20916 22372
rect 20860 22318 20862 22370
rect 20862 22318 20914 22370
rect 20914 22318 20916 22370
rect 20860 22316 20916 22318
rect 21308 34018 21364 34020
rect 21308 33966 21310 34018
rect 21310 33966 21362 34018
rect 21362 33966 21364 34018
rect 21308 33964 21364 33966
rect 21308 33068 21364 33124
rect 21308 32620 21364 32676
rect 21308 30940 21364 30996
rect 22092 36428 22148 36484
rect 21980 34690 22036 34692
rect 21980 34638 21982 34690
rect 21982 34638 22034 34690
rect 22034 34638 22036 34690
rect 21980 34636 22036 34638
rect 21644 34130 21700 34132
rect 21644 34078 21646 34130
rect 21646 34078 21698 34130
rect 21698 34078 21700 34130
rect 21644 34076 21700 34078
rect 21644 33852 21700 33908
rect 22428 36316 22484 36372
rect 22204 36092 22260 36148
rect 22204 35922 22260 35924
rect 22204 35870 22206 35922
rect 22206 35870 22258 35922
rect 22258 35870 22260 35922
rect 22204 35868 22260 35870
rect 22764 37436 22820 37492
rect 22988 37436 23044 37492
rect 22876 36258 22932 36260
rect 22876 36206 22878 36258
rect 22878 36206 22930 36258
rect 22930 36206 22932 36258
rect 22876 36204 22932 36206
rect 22652 35586 22708 35588
rect 22652 35534 22654 35586
rect 22654 35534 22706 35586
rect 22706 35534 22708 35586
rect 22652 35532 22708 35534
rect 22092 33404 22148 33460
rect 21756 32620 21812 32676
rect 21868 32396 21924 32452
rect 22092 32732 22148 32788
rect 22092 32396 22148 32452
rect 21756 31836 21812 31892
rect 21980 31778 22036 31780
rect 21980 31726 21982 31778
rect 21982 31726 22034 31778
rect 22034 31726 22036 31778
rect 21980 31724 22036 31726
rect 21644 31218 21700 31220
rect 21644 31166 21646 31218
rect 21646 31166 21698 31218
rect 21698 31166 21700 31218
rect 21644 31164 21700 31166
rect 21868 31106 21924 31108
rect 21868 31054 21870 31106
rect 21870 31054 21922 31106
rect 21922 31054 21924 31106
rect 21868 31052 21924 31054
rect 22204 31836 22260 31892
rect 22652 33852 22708 33908
rect 22764 33964 22820 34020
rect 22204 31554 22260 31556
rect 22204 31502 22206 31554
rect 22206 31502 22258 31554
rect 22258 31502 22260 31554
rect 22204 31500 22260 31502
rect 22092 30940 22148 30996
rect 21644 30492 21700 30548
rect 21756 30828 21812 30884
rect 21532 29986 21588 29988
rect 21532 29934 21534 29986
rect 21534 29934 21586 29986
rect 21586 29934 21588 29986
rect 21532 29932 21588 29934
rect 21196 28252 21252 28308
rect 21980 30044 22036 30100
rect 22540 33404 22596 33460
rect 22316 30044 22372 30100
rect 22092 29708 22148 29764
rect 22428 29820 22484 29876
rect 21980 29484 22036 29540
rect 22428 28700 22484 28756
rect 22204 28530 22260 28532
rect 22204 28478 22206 28530
rect 22206 28478 22258 28530
rect 22258 28478 22260 28530
rect 22204 28476 22260 28478
rect 22876 33346 22932 33348
rect 22876 33294 22878 33346
rect 22878 33294 22930 33346
rect 22930 33294 22932 33346
rect 22876 33292 22932 33294
rect 22876 32956 22932 33012
rect 23100 34018 23156 34020
rect 23100 33966 23102 34018
rect 23102 33966 23154 34018
rect 23154 33966 23156 34018
rect 23100 33964 23156 33966
rect 23324 39676 23380 39732
rect 23324 35868 23380 35924
rect 23212 33628 23268 33684
rect 23100 33122 23156 33124
rect 23100 33070 23102 33122
rect 23102 33070 23154 33122
rect 23154 33070 23156 33122
rect 23100 33068 23156 33070
rect 23996 43708 24052 43764
rect 23660 42754 23716 42756
rect 23660 42702 23662 42754
rect 23662 42702 23714 42754
rect 23714 42702 23716 42754
rect 23660 42700 23716 42702
rect 23660 42364 23716 42420
rect 23772 41804 23828 41860
rect 23548 39788 23604 39844
rect 23660 40402 23716 40404
rect 23660 40350 23662 40402
rect 23662 40350 23714 40402
rect 23714 40350 23716 40402
rect 23660 40348 23716 40350
rect 23548 39004 23604 39060
rect 23548 38444 23604 38500
rect 23548 37884 23604 37940
rect 24108 43372 24164 43428
rect 24108 42028 24164 42084
rect 24220 41970 24276 41972
rect 24220 41918 24222 41970
rect 24222 41918 24274 41970
rect 24274 41918 24276 41970
rect 24220 41916 24276 41918
rect 24892 45500 24948 45556
rect 24668 44546 24724 44548
rect 24668 44494 24670 44546
rect 24670 44494 24722 44546
rect 24722 44494 24724 44546
rect 24668 44492 24724 44494
rect 25004 45330 25060 45332
rect 25004 45278 25006 45330
rect 25006 45278 25058 45330
rect 25058 45278 25060 45330
rect 25004 45276 25060 45278
rect 25004 44716 25060 44772
rect 25676 50034 25732 50036
rect 25676 49982 25678 50034
rect 25678 49982 25730 50034
rect 25730 49982 25732 50034
rect 25676 49980 25732 49982
rect 25452 48914 25508 48916
rect 25452 48862 25454 48914
rect 25454 48862 25506 48914
rect 25506 48862 25508 48914
rect 25452 48860 25508 48862
rect 26124 51378 26180 51380
rect 26124 51326 26126 51378
rect 26126 51326 26178 51378
rect 26178 51326 26180 51378
rect 26124 51324 26180 51326
rect 27020 52946 27076 52948
rect 27020 52894 27022 52946
rect 27022 52894 27074 52946
rect 27074 52894 27076 52946
rect 27020 52892 27076 52894
rect 26796 52556 26852 52612
rect 27244 52780 27300 52836
rect 26460 50876 26516 50932
rect 26012 50316 26068 50372
rect 26236 50428 26292 50484
rect 25676 48636 25732 48692
rect 26012 48972 26068 49028
rect 25788 48524 25844 48580
rect 25676 47964 25732 48020
rect 25564 47180 25620 47236
rect 25676 47404 25732 47460
rect 26012 47292 26068 47348
rect 25676 46844 25732 46900
rect 25900 46844 25956 46900
rect 25788 46508 25844 46564
rect 25340 46172 25396 46228
rect 25452 45890 25508 45892
rect 25452 45838 25454 45890
rect 25454 45838 25506 45890
rect 25506 45838 25508 45890
rect 25452 45836 25508 45838
rect 25340 45666 25396 45668
rect 25340 45614 25342 45666
rect 25342 45614 25394 45666
rect 25394 45614 25396 45666
rect 25340 45612 25396 45614
rect 25788 45778 25844 45780
rect 25788 45726 25790 45778
rect 25790 45726 25842 45778
rect 25842 45726 25844 45778
rect 25788 45724 25844 45726
rect 25564 45612 25620 45668
rect 25228 45276 25284 45332
rect 25676 45106 25732 45108
rect 25676 45054 25678 45106
rect 25678 45054 25730 45106
rect 25730 45054 25732 45106
rect 25676 45052 25732 45054
rect 25228 44604 25284 44660
rect 24556 43484 24612 43540
rect 24780 43932 24836 43988
rect 24668 42028 24724 42084
rect 24556 41746 24612 41748
rect 24556 41694 24558 41746
rect 24558 41694 24610 41746
rect 24610 41694 24612 41746
rect 24556 41692 24612 41694
rect 24444 41580 24500 41636
rect 25116 43708 25172 43764
rect 24332 40796 24388 40852
rect 24892 42588 24948 42644
rect 23996 40572 24052 40628
rect 24444 40572 24500 40628
rect 23772 38444 23828 38500
rect 23884 39618 23940 39620
rect 23884 39566 23886 39618
rect 23886 39566 23938 39618
rect 23938 39566 23940 39618
rect 23884 39564 23940 39566
rect 23996 38946 24052 38948
rect 23996 38894 23998 38946
rect 23998 38894 24050 38946
rect 24050 38894 24052 38946
rect 23996 38892 24052 38894
rect 23996 37884 24052 37940
rect 24108 37772 24164 37828
rect 23996 36092 24052 36148
rect 23548 34412 23604 34468
rect 23548 32620 23604 32676
rect 23212 32396 23268 32452
rect 22876 31890 22932 31892
rect 22876 31838 22878 31890
rect 22878 31838 22930 31890
rect 22930 31838 22932 31890
rect 22876 31836 22932 31838
rect 22764 31276 22820 31332
rect 23100 31836 23156 31892
rect 22652 30882 22708 30884
rect 22652 30830 22654 30882
rect 22654 30830 22706 30882
rect 22706 30830 22708 30882
rect 22652 30828 22708 30830
rect 22652 30210 22708 30212
rect 22652 30158 22654 30210
rect 22654 30158 22706 30210
rect 22706 30158 22708 30210
rect 22652 30156 22708 30158
rect 22764 28924 22820 28980
rect 21084 21980 21140 22036
rect 20748 21644 20804 21700
rect 21868 25676 21924 25732
rect 21420 25116 21476 25172
rect 22092 26236 22148 26292
rect 21868 24556 21924 24612
rect 21420 23884 21476 23940
rect 21308 23154 21364 23156
rect 21308 23102 21310 23154
rect 21310 23102 21362 23154
rect 21362 23102 21364 23154
rect 21308 23100 21364 23102
rect 21644 22482 21700 22484
rect 21644 22430 21646 22482
rect 21646 22430 21698 22482
rect 21698 22430 21700 22482
rect 21644 22428 21700 22430
rect 21420 22316 21476 22372
rect 21308 21420 21364 21476
rect 21644 21980 21700 22036
rect 21532 21868 21588 21924
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19628 18338 19684 18340
rect 19628 18286 19630 18338
rect 19630 18286 19682 18338
rect 19682 18286 19684 18338
rect 19628 18284 19684 18286
rect 18956 16268 19012 16324
rect 17948 14476 18004 14532
rect 18508 15314 18564 15316
rect 18508 15262 18510 15314
rect 18510 15262 18562 15314
rect 18562 15262 18564 15314
rect 18508 15260 18564 15262
rect 19628 17778 19684 17780
rect 19628 17726 19630 17778
rect 19630 17726 19682 17778
rect 19682 17726 19684 17778
rect 19628 17724 19684 17726
rect 19180 17666 19236 17668
rect 19180 17614 19182 17666
rect 19182 17614 19234 17666
rect 19234 17614 19236 17666
rect 19180 17612 19236 17614
rect 20076 18172 20132 18228
rect 19740 17612 19796 17668
rect 20188 17724 20244 17780
rect 20524 17778 20580 17780
rect 20524 17726 20526 17778
rect 20526 17726 20578 17778
rect 20578 17726 20580 17778
rect 20524 17724 20580 17726
rect 19852 17500 19908 17556
rect 20188 17388 20244 17444
rect 19180 17106 19236 17108
rect 19180 17054 19182 17106
rect 19182 17054 19234 17106
rect 19234 17054 19236 17106
rect 19180 17052 19236 17054
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19628 16156 19684 16212
rect 19852 16210 19908 16212
rect 19852 16158 19854 16210
rect 19854 16158 19906 16210
rect 19906 16158 19908 16210
rect 19852 16156 19908 16158
rect 20972 17778 21028 17780
rect 20972 17726 20974 17778
rect 20974 17726 21026 17778
rect 21026 17726 21028 17778
rect 20972 17724 21028 17726
rect 20860 17164 20916 17220
rect 20972 17500 21028 17556
rect 20524 17106 20580 17108
rect 20524 17054 20526 17106
rect 20526 17054 20578 17106
rect 20578 17054 20580 17106
rect 20524 17052 20580 17054
rect 21308 17276 21364 17332
rect 21420 17164 21476 17220
rect 21084 16940 21140 16996
rect 20412 16268 20468 16324
rect 20860 16268 20916 16324
rect 20188 15932 20244 15988
rect 21420 15932 21476 15988
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 16044 14252 16100 14308
rect 16268 13746 16324 13748
rect 16268 13694 16270 13746
rect 16270 13694 16322 13746
rect 16322 13694 16324 13746
rect 16268 13692 16324 13694
rect 18284 13356 18340 13412
rect 15372 12684 15428 12740
rect 19180 13356 19236 13412
rect 19068 13186 19124 13188
rect 19068 13134 19070 13186
rect 19070 13134 19122 13186
rect 19122 13134 19124 13186
rect 19068 13132 19124 13134
rect 17052 12348 17108 12404
rect 14140 10556 14196 10612
rect 14028 10444 14084 10500
rect 13916 9548 13972 9604
rect 13804 7644 13860 7700
rect 15036 8988 15092 9044
rect 12796 6076 12852 6132
rect 16044 12236 16100 12292
rect 16492 11900 16548 11956
rect 18732 13020 18788 13076
rect 18284 11900 18340 11956
rect 21196 15314 21252 15316
rect 21196 15262 21198 15314
rect 21198 15262 21250 15314
rect 21250 15262 21252 15314
rect 21196 15260 21252 15262
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19628 13074 19684 13076
rect 19628 13022 19630 13074
rect 19630 13022 19682 13074
rect 19682 13022 19684 13074
rect 19628 13020 19684 13022
rect 19180 12066 19236 12068
rect 19180 12014 19182 12066
rect 19182 12014 19234 12066
rect 19234 12014 19236 12066
rect 19180 12012 19236 12014
rect 19292 12908 19348 12964
rect 18508 11564 18564 11620
rect 15932 10668 15988 10724
rect 17612 10610 17668 10612
rect 17612 10558 17614 10610
rect 17614 10558 17666 10610
rect 17666 10558 17668 10610
rect 17612 10556 17668 10558
rect 19068 11506 19124 11508
rect 19068 11454 19070 11506
rect 19070 11454 19122 11506
rect 19122 11454 19124 11506
rect 19068 11452 19124 11454
rect 18508 10498 18564 10500
rect 18508 10446 18510 10498
rect 18510 10446 18562 10498
rect 18562 10446 18564 10498
rect 18508 10444 18564 10446
rect 19740 12908 19796 12964
rect 20188 13020 20244 13076
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 20524 12962 20580 12964
rect 20524 12910 20526 12962
rect 20526 12910 20578 12962
rect 20578 12910 20580 12962
rect 20524 12908 20580 12910
rect 21420 12290 21476 12292
rect 21420 12238 21422 12290
rect 21422 12238 21474 12290
rect 21474 12238 21476 12290
rect 21420 12236 21476 12238
rect 19628 12012 19684 12068
rect 22764 27858 22820 27860
rect 22764 27806 22766 27858
rect 22766 27806 22818 27858
rect 22818 27806 22820 27858
rect 22764 27804 22820 27806
rect 22540 26348 22596 26404
rect 22204 23660 22260 23716
rect 22316 25228 22372 25284
rect 22540 23772 22596 23828
rect 22428 23436 22484 23492
rect 21980 23212 22036 23268
rect 21980 22316 22036 22372
rect 21756 21644 21812 21700
rect 22316 23266 22372 23268
rect 22316 23214 22318 23266
rect 22318 23214 22370 23266
rect 22370 23214 22372 23266
rect 22316 23212 22372 23214
rect 21756 21420 21812 21476
rect 21756 20524 21812 20580
rect 22204 21362 22260 21364
rect 22204 21310 22206 21362
rect 22206 21310 22258 21362
rect 22258 21310 22260 21362
rect 22204 21308 22260 21310
rect 21980 21196 22036 21252
rect 21980 20636 22036 20692
rect 22428 21084 22484 21140
rect 22540 21756 22596 21812
rect 22092 20802 22148 20804
rect 22092 20750 22094 20802
rect 22094 20750 22146 20802
rect 22146 20750 22148 20802
rect 22092 20748 22148 20750
rect 22092 20300 22148 20356
rect 22764 26402 22820 26404
rect 22764 26350 22766 26402
rect 22766 26350 22818 26402
rect 22818 26350 22820 26402
rect 22764 26348 22820 26350
rect 22764 25788 22820 25844
rect 22988 30044 23044 30100
rect 23884 34412 23940 34468
rect 23772 31612 23828 31668
rect 23660 30604 23716 30660
rect 23212 30156 23268 30212
rect 23436 30044 23492 30100
rect 23548 29148 23604 29204
rect 23772 29148 23828 29204
rect 24332 38332 24388 38388
rect 24556 37884 24612 37940
rect 24332 36988 24388 37044
rect 24444 36258 24500 36260
rect 24444 36206 24446 36258
rect 24446 36206 24498 36258
rect 24498 36206 24500 36258
rect 24444 36204 24500 36206
rect 24108 34300 24164 34356
rect 24220 33964 24276 34020
rect 23996 33628 24052 33684
rect 24332 34412 24388 34468
rect 24444 34748 24500 34804
rect 24444 34076 24500 34132
rect 24332 33180 24388 33236
rect 24332 32562 24388 32564
rect 24332 32510 24334 32562
rect 24334 32510 24386 32562
rect 24386 32510 24388 32562
rect 24332 32508 24388 32510
rect 24108 32450 24164 32452
rect 24108 32398 24110 32450
rect 24110 32398 24162 32450
rect 24162 32398 24164 32450
rect 24108 32396 24164 32398
rect 24556 32338 24612 32340
rect 24556 32286 24558 32338
rect 24558 32286 24610 32338
rect 24610 32286 24612 32338
rect 24556 32284 24612 32286
rect 23996 31724 24052 31780
rect 23996 31218 24052 31220
rect 23996 31166 23998 31218
rect 23998 31166 24050 31218
rect 24050 31166 24052 31218
rect 23996 31164 24052 31166
rect 24444 31890 24500 31892
rect 24444 31838 24446 31890
rect 24446 31838 24498 31890
rect 24498 31838 24500 31890
rect 24444 31836 24500 31838
rect 24444 30882 24500 30884
rect 24444 30830 24446 30882
rect 24446 30830 24498 30882
rect 24498 30830 24500 30882
rect 24444 30828 24500 30830
rect 24556 30492 24612 30548
rect 24444 30380 24500 30436
rect 24220 30098 24276 30100
rect 24220 30046 24222 30098
rect 24222 30046 24274 30098
rect 24274 30046 24276 30098
rect 24220 30044 24276 30046
rect 23772 28476 23828 28532
rect 23660 28364 23716 28420
rect 24220 28476 24276 28532
rect 24108 28364 24164 28420
rect 23996 27020 24052 27076
rect 23884 26572 23940 26628
rect 23548 26290 23604 26292
rect 23548 26238 23550 26290
rect 23550 26238 23602 26290
rect 23602 26238 23604 26290
rect 23548 26236 23604 26238
rect 22988 25900 23044 25956
rect 23660 25676 23716 25732
rect 23548 25618 23604 25620
rect 23548 25566 23550 25618
rect 23550 25566 23602 25618
rect 23602 25566 23604 25618
rect 23548 25564 23604 25566
rect 22988 23714 23044 23716
rect 22988 23662 22990 23714
rect 22990 23662 23042 23714
rect 23042 23662 23044 23714
rect 22988 23660 23044 23662
rect 23100 23212 23156 23268
rect 23660 23548 23716 23604
rect 22876 21756 22932 21812
rect 23660 23042 23716 23044
rect 23660 22990 23662 23042
rect 23662 22990 23714 23042
rect 23714 22990 23716 23042
rect 23660 22988 23716 22990
rect 23548 22092 23604 22148
rect 23100 21698 23156 21700
rect 23100 21646 23102 21698
rect 23102 21646 23154 21698
rect 23154 21646 23156 21698
rect 23100 21644 23156 21646
rect 22652 21196 22708 21252
rect 21644 18284 21700 18340
rect 22652 19964 22708 20020
rect 22204 19794 22260 19796
rect 22204 19742 22206 19794
rect 22206 19742 22258 19794
rect 22258 19742 22260 19794
rect 22204 19740 22260 19742
rect 23324 21868 23380 21924
rect 23212 21532 23268 21588
rect 25116 42866 25172 42868
rect 25116 42814 25118 42866
rect 25118 42814 25170 42866
rect 25170 42814 25172 42866
rect 25116 42812 25172 42814
rect 25004 41244 25060 41300
rect 24780 40236 24836 40292
rect 25676 44492 25732 44548
rect 25788 44604 25844 44660
rect 25452 43372 25508 43428
rect 25228 41804 25284 41860
rect 25228 41244 25284 41300
rect 25340 42812 25396 42868
rect 25228 41074 25284 41076
rect 25228 41022 25230 41074
rect 25230 41022 25282 41074
rect 25282 41022 25284 41074
rect 25228 41020 25284 41022
rect 25116 39730 25172 39732
rect 25116 39678 25118 39730
rect 25118 39678 25170 39730
rect 25170 39678 25172 39730
rect 25116 39676 25172 39678
rect 25004 38332 25060 38388
rect 25004 35868 25060 35924
rect 24780 34412 24836 34468
rect 24892 34018 24948 34020
rect 24892 33966 24894 34018
rect 24894 33966 24946 34018
rect 24946 33966 24948 34018
rect 24892 33964 24948 33966
rect 25340 40348 25396 40404
rect 25564 43260 25620 43316
rect 25676 43036 25732 43092
rect 26012 45948 26068 46004
rect 26012 44882 26068 44884
rect 26012 44830 26014 44882
rect 26014 44830 26066 44882
rect 26066 44830 26068 44882
rect 26012 44828 26068 44830
rect 26012 43820 26068 43876
rect 27132 52050 27188 52052
rect 27132 51998 27134 52050
rect 27134 51998 27186 52050
rect 27186 51998 27188 52050
rect 27132 51996 27188 51998
rect 29820 58604 29876 58660
rect 30156 59330 30212 59332
rect 30156 59278 30158 59330
rect 30158 59278 30210 59330
rect 30210 59278 30212 59330
rect 30156 59276 30212 59278
rect 30716 59330 30772 59332
rect 30716 59278 30718 59330
rect 30718 59278 30770 59330
rect 30770 59278 30772 59330
rect 30716 59276 30772 59278
rect 30828 59218 30884 59220
rect 30828 59166 30830 59218
rect 30830 59166 30882 59218
rect 30882 59166 30884 59218
rect 30828 59164 30884 59166
rect 30716 58994 30772 58996
rect 30716 58942 30718 58994
rect 30718 58942 30770 58994
rect 30770 58942 30772 58994
rect 30716 58940 30772 58942
rect 30044 58716 30100 58772
rect 31276 58716 31332 58772
rect 30156 58658 30212 58660
rect 30156 58606 30158 58658
rect 30158 58606 30210 58658
rect 30210 58606 30212 58658
rect 30156 58604 30212 58606
rect 30604 58604 30660 58660
rect 30492 58434 30548 58436
rect 30492 58382 30494 58434
rect 30494 58382 30546 58434
rect 30546 58382 30548 58434
rect 30492 58380 30548 58382
rect 30044 57708 30100 57764
rect 28812 56866 28868 56868
rect 28812 56814 28814 56866
rect 28814 56814 28866 56866
rect 28866 56814 28868 56866
rect 28812 56812 28868 56814
rect 28028 56700 28084 56756
rect 28588 56754 28644 56756
rect 28588 56702 28590 56754
rect 28590 56702 28642 56754
rect 28642 56702 28644 56754
rect 28588 56700 28644 56702
rect 29260 56476 29316 56532
rect 28140 54514 28196 54516
rect 28140 54462 28142 54514
rect 28142 54462 28194 54514
rect 28194 54462 28196 54514
rect 28140 54460 28196 54462
rect 28476 55580 28532 55636
rect 28476 55020 28532 55076
rect 29036 54514 29092 54516
rect 29036 54462 29038 54514
rect 29038 54462 29090 54514
rect 29090 54462 29092 54514
rect 29036 54460 29092 54462
rect 28700 53676 28756 53732
rect 28252 53564 28308 53620
rect 27916 52108 27972 52164
rect 28028 53340 28084 53396
rect 27244 50764 27300 50820
rect 26908 50594 26964 50596
rect 26908 50542 26910 50594
rect 26910 50542 26962 50594
rect 26962 50542 26964 50594
rect 26908 50540 26964 50542
rect 27804 51996 27860 52052
rect 27244 50540 27300 50596
rect 27356 49756 27412 49812
rect 26460 49308 26516 49364
rect 26348 49138 26404 49140
rect 26348 49086 26350 49138
rect 26350 49086 26402 49138
rect 26402 49086 26404 49138
rect 26348 49084 26404 49086
rect 26236 46956 26292 47012
rect 26348 48860 26404 48916
rect 27020 49196 27076 49252
rect 26236 46674 26292 46676
rect 26236 46622 26238 46674
rect 26238 46622 26290 46674
rect 26290 46622 26292 46674
rect 26236 46620 26292 46622
rect 26796 48802 26852 48804
rect 26796 48750 26798 48802
rect 26798 48750 26850 48802
rect 26850 48750 26852 48802
rect 26796 48748 26852 48750
rect 26684 48524 26740 48580
rect 26572 48354 26628 48356
rect 26572 48302 26574 48354
rect 26574 48302 26626 48354
rect 26626 48302 26628 48354
rect 26572 48300 26628 48302
rect 26348 46060 26404 46116
rect 26348 44604 26404 44660
rect 26460 44322 26516 44324
rect 26460 44270 26462 44322
rect 26462 44270 26514 44322
rect 26514 44270 26516 44322
rect 26460 44268 26516 44270
rect 26348 44210 26404 44212
rect 26348 44158 26350 44210
rect 26350 44158 26402 44210
rect 26402 44158 26404 44210
rect 26348 44156 26404 44158
rect 26908 46172 26964 46228
rect 26908 46002 26964 46004
rect 26908 45950 26910 46002
rect 26910 45950 26962 46002
rect 26962 45950 26964 46002
rect 26908 45948 26964 45950
rect 26796 45164 26852 45220
rect 26908 45724 26964 45780
rect 27132 48748 27188 48804
rect 27356 48748 27412 48804
rect 27356 48076 27412 48132
rect 27356 47458 27412 47460
rect 27356 47406 27358 47458
rect 27358 47406 27410 47458
rect 27410 47406 27412 47458
rect 27356 47404 27412 47406
rect 29036 53058 29092 53060
rect 29036 53006 29038 53058
rect 29038 53006 29090 53058
rect 29090 53006 29092 53058
rect 29036 53004 29092 53006
rect 28588 52892 28644 52948
rect 28364 52444 28420 52500
rect 28252 52108 28308 52164
rect 28028 51324 28084 51380
rect 28028 50764 28084 50820
rect 27916 50540 27972 50596
rect 28028 50092 28084 50148
rect 27916 49810 27972 49812
rect 27916 49758 27918 49810
rect 27918 49758 27970 49810
rect 27970 49758 27972 49810
rect 27916 49756 27972 49758
rect 27916 49138 27972 49140
rect 27916 49086 27918 49138
rect 27918 49086 27970 49138
rect 27970 49086 27972 49138
rect 27916 49084 27972 49086
rect 27580 47346 27636 47348
rect 27580 47294 27582 47346
rect 27582 47294 27634 47346
rect 27634 47294 27636 47346
rect 27580 47292 27636 47294
rect 27916 47292 27972 47348
rect 27804 46562 27860 46564
rect 27804 46510 27806 46562
rect 27806 46510 27858 46562
rect 27858 46510 27860 46562
rect 27804 46508 27860 46510
rect 27468 46172 27524 46228
rect 27020 45052 27076 45108
rect 27356 45276 27412 45332
rect 26236 43036 26292 43092
rect 26460 43820 26516 43876
rect 25676 42252 25732 42308
rect 25788 42476 25844 42532
rect 25564 40236 25620 40292
rect 25452 39340 25508 39396
rect 25228 36092 25284 36148
rect 25340 34412 25396 34468
rect 25116 32396 25172 32452
rect 25004 32338 25060 32340
rect 25004 32286 25006 32338
rect 25006 32286 25058 32338
rect 25058 32286 25060 32338
rect 25004 32284 25060 32286
rect 25116 31612 25172 31668
rect 25004 30940 25060 30996
rect 24780 30380 24836 30436
rect 25116 30828 25172 30884
rect 26124 42588 26180 42644
rect 25900 42252 25956 42308
rect 25900 40796 25956 40852
rect 26460 42476 26516 42532
rect 27244 44716 27300 44772
rect 27132 43820 27188 43876
rect 27020 43708 27076 43764
rect 26908 43596 26964 43652
rect 26796 43426 26852 43428
rect 26796 43374 26798 43426
rect 26798 43374 26850 43426
rect 26850 43374 26852 43426
rect 26796 43372 26852 43374
rect 26684 42866 26740 42868
rect 26684 42814 26686 42866
rect 26686 42814 26738 42866
rect 26738 42814 26740 42866
rect 26684 42812 26740 42814
rect 27580 44716 27636 44772
rect 27468 44322 27524 44324
rect 27468 44270 27470 44322
rect 27470 44270 27522 44322
rect 27522 44270 27524 44322
rect 27468 44268 27524 44270
rect 27804 45106 27860 45108
rect 27804 45054 27806 45106
rect 27806 45054 27858 45106
rect 27858 45054 27860 45106
rect 27804 45052 27860 45054
rect 28252 50482 28308 50484
rect 28252 50430 28254 50482
rect 28254 50430 28306 50482
rect 28306 50430 28308 50482
rect 28252 50428 28308 50430
rect 28364 49196 28420 49252
rect 28364 48412 28420 48468
rect 28252 48300 28308 48356
rect 28140 46620 28196 46676
rect 28364 47180 28420 47236
rect 28252 47068 28308 47124
rect 28140 46396 28196 46452
rect 28476 46396 28532 46452
rect 28028 45948 28084 46004
rect 28252 46172 28308 46228
rect 28252 45724 28308 45780
rect 28028 45276 28084 45332
rect 28140 45612 28196 45668
rect 28028 45052 28084 45108
rect 28028 44716 28084 44772
rect 27356 43484 27412 43540
rect 27244 43426 27300 43428
rect 27244 43374 27246 43426
rect 27246 43374 27298 43426
rect 27298 43374 27300 43426
rect 27244 43372 27300 43374
rect 26796 42754 26852 42756
rect 26796 42702 26798 42754
rect 26798 42702 26850 42754
rect 26850 42702 26852 42754
rect 26796 42700 26852 42702
rect 26236 40348 26292 40404
rect 26124 40124 26180 40180
rect 26684 41692 26740 41748
rect 26460 41074 26516 41076
rect 26460 41022 26462 41074
rect 26462 41022 26514 41074
rect 26514 41022 26516 41074
rect 26460 41020 26516 41022
rect 26572 40572 26628 40628
rect 26796 40572 26852 40628
rect 27020 41356 27076 41412
rect 26908 40460 26964 40516
rect 26348 39788 26404 39844
rect 26124 39452 26180 39508
rect 25788 38892 25844 38948
rect 25900 38668 25956 38724
rect 26348 38892 26404 38948
rect 25676 38108 25732 38164
rect 26124 37884 26180 37940
rect 26124 37100 26180 37156
rect 25564 35644 25620 35700
rect 26012 36370 26068 36372
rect 26012 36318 26014 36370
rect 26014 36318 26066 36370
rect 26066 36318 26068 36370
rect 26012 36316 26068 36318
rect 25900 36204 25956 36260
rect 26572 38444 26628 38500
rect 26348 37266 26404 37268
rect 26348 37214 26350 37266
rect 26350 37214 26402 37266
rect 26402 37214 26404 37266
rect 26348 37212 26404 37214
rect 26572 36482 26628 36484
rect 26572 36430 26574 36482
rect 26574 36430 26626 36482
rect 26626 36430 26628 36482
rect 26572 36428 26628 36430
rect 25788 35980 25844 36036
rect 25788 35698 25844 35700
rect 25788 35646 25790 35698
rect 25790 35646 25842 35698
rect 25842 35646 25844 35698
rect 25788 35644 25844 35646
rect 26124 36092 26180 36148
rect 26012 35922 26068 35924
rect 26012 35870 26014 35922
rect 26014 35870 26066 35922
rect 26066 35870 26068 35922
rect 26012 35868 26068 35870
rect 25676 35196 25732 35252
rect 25564 33852 25620 33908
rect 25676 34972 25732 35028
rect 25676 33740 25732 33796
rect 26348 35532 26404 35588
rect 26460 35308 26516 35364
rect 26348 34690 26404 34692
rect 26348 34638 26350 34690
rect 26350 34638 26402 34690
rect 26402 34638 26404 34690
rect 26348 34636 26404 34638
rect 26012 34354 26068 34356
rect 26012 34302 26014 34354
rect 26014 34302 26066 34354
rect 26066 34302 26068 34354
rect 26012 34300 26068 34302
rect 25452 31948 25508 32004
rect 26236 32844 26292 32900
rect 26460 34242 26516 34244
rect 26460 34190 26462 34242
rect 26462 34190 26514 34242
rect 26514 34190 26516 34242
rect 26460 34188 26516 34190
rect 26460 33852 26516 33908
rect 27132 40962 27188 40964
rect 27132 40910 27134 40962
rect 27134 40910 27186 40962
rect 27186 40910 27188 40962
rect 27132 40908 27188 40910
rect 27244 40460 27300 40516
rect 27132 40402 27188 40404
rect 27132 40350 27134 40402
rect 27134 40350 27186 40402
rect 27186 40350 27188 40402
rect 27132 40348 27188 40350
rect 27244 40012 27300 40068
rect 27468 42140 27524 42196
rect 27916 44434 27972 44436
rect 27916 44382 27918 44434
rect 27918 44382 27970 44434
rect 27970 44382 27972 44434
rect 27916 44380 27972 44382
rect 28028 43932 28084 43988
rect 28700 51996 28756 52052
rect 28700 50428 28756 50484
rect 30716 58156 30772 58212
rect 30492 56866 30548 56868
rect 30492 56814 30494 56866
rect 30494 56814 30546 56866
rect 30546 56814 30548 56866
rect 30492 56812 30548 56814
rect 30044 56700 30100 56756
rect 32844 59218 32900 59220
rect 32844 59166 32846 59218
rect 32846 59166 32898 59218
rect 32898 59166 32900 59218
rect 32844 59164 32900 59166
rect 33740 59612 33796 59668
rect 35532 59778 35588 59780
rect 35532 59726 35534 59778
rect 35534 59726 35586 59778
rect 35586 59726 35588 59778
rect 35532 59724 35588 59726
rect 36316 59724 36372 59780
rect 33964 59218 34020 59220
rect 33964 59166 33966 59218
rect 33966 59166 34018 59218
rect 34018 59166 34020 59218
rect 33964 59164 34020 59166
rect 33852 59052 33908 59108
rect 32732 58492 32788 58548
rect 32844 58940 32900 58996
rect 32508 58380 32564 58436
rect 32060 58156 32116 58212
rect 32284 58322 32340 58324
rect 32284 58270 32286 58322
rect 32286 58270 32338 58322
rect 32338 58270 32340 58322
rect 32284 58268 32340 58270
rect 31164 57650 31220 57652
rect 31164 57598 31166 57650
rect 31166 57598 31218 57650
rect 31218 57598 31220 57650
rect 31164 57596 31220 57598
rect 31724 57484 31780 57540
rect 31500 56924 31556 56980
rect 31500 56754 31556 56756
rect 31500 56702 31502 56754
rect 31502 56702 31554 56754
rect 31554 56702 31556 56754
rect 31500 56700 31556 56702
rect 31052 56588 31108 56644
rect 31388 56476 31444 56532
rect 31276 55970 31332 55972
rect 31276 55918 31278 55970
rect 31278 55918 31330 55970
rect 31330 55918 31332 55970
rect 31276 55916 31332 55918
rect 29708 53842 29764 53844
rect 29708 53790 29710 53842
rect 29710 53790 29762 53842
rect 29762 53790 29764 53842
rect 29708 53788 29764 53790
rect 29596 53730 29652 53732
rect 29596 53678 29598 53730
rect 29598 53678 29650 53730
rect 29650 53678 29652 53730
rect 29596 53676 29652 53678
rect 30156 54514 30212 54516
rect 30156 54462 30158 54514
rect 30158 54462 30210 54514
rect 30210 54462 30212 54514
rect 30156 54460 30212 54462
rect 30940 54684 30996 54740
rect 30828 54402 30884 54404
rect 30828 54350 30830 54402
rect 30830 54350 30882 54402
rect 30882 54350 30884 54402
rect 30828 54348 30884 54350
rect 29932 53676 29988 53732
rect 29708 52162 29764 52164
rect 29708 52110 29710 52162
rect 29710 52110 29762 52162
rect 29762 52110 29764 52162
rect 29708 52108 29764 52110
rect 30604 53676 30660 53732
rect 30044 51660 30100 51716
rect 30156 51548 30212 51604
rect 30716 51660 30772 51716
rect 28924 50316 28980 50372
rect 28812 49138 28868 49140
rect 28812 49086 28814 49138
rect 28814 49086 28866 49138
rect 28866 49086 28868 49138
rect 28812 49084 28868 49086
rect 28812 48076 28868 48132
rect 28812 47570 28868 47572
rect 28812 47518 28814 47570
rect 28814 47518 28866 47570
rect 28866 47518 28868 47570
rect 28812 47516 28868 47518
rect 28924 46620 28980 46676
rect 29148 49644 29204 49700
rect 28700 46508 28756 46564
rect 28588 46172 28644 46228
rect 28588 45612 28644 45668
rect 28812 45500 28868 45556
rect 28700 44828 28756 44884
rect 28252 43932 28308 43988
rect 28140 43762 28196 43764
rect 28140 43710 28142 43762
rect 28142 43710 28194 43762
rect 28194 43710 28196 43762
rect 28140 43708 28196 43710
rect 27916 43538 27972 43540
rect 27916 43486 27918 43538
rect 27918 43486 27970 43538
rect 27970 43486 27972 43538
rect 27916 43484 27972 43486
rect 28476 43650 28532 43652
rect 28476 43598 28478 43650
rect 28478 43598 28530 43650
rect 28530 43598 28532 43650
rect 28476 43596 28532 43598
rect 27916 42866 27972 42868
rect 27916 42814 27918 42866
rect 27918 42814 27970 42866
rect 27970 42814 27972 42866
rect 27916 42812 27972 42814
rect 28028 42476 28084 42532
rect 28028 41916 28084 41972
rect 27916 41410 27972 41412
rect 27916 41358 27918 41410
rect 27918 41358 27970 41410
rect 27970 41358 27972 41410
rect 27916 41356 27972 41358
rect 28364 41468 28420 41524
rect 28476 42028 28532 42084
rect 28252 41410 28308 41412
rect 28252 41358 28254 41410
rect 28254 41358 28306 41410
rect 28306 41358 28308 41410
rect 28252 41356 28308 41358
rect 27356 39900 27412 39956
rect 27580 40684 27636 40740
rect 27020 37212 27076 37268
rect 27132 39564 27188 39620
rect 26796 35420 26852 35476
rect 27020 35084 27076 35140
rect 27804 40684 27860 40740
rect 28028 40626 28084 40628
rect 28028 40574 28030 40626
rect 28030 40574 28082 40626
rect 28082 40574 28084 40626
rect 28028 40572 28084 40574
rect 27692 40514 27748 40516
rect 27692 40462 27694 40514
rect 27694 40462 27746 40514
rect 27746 40462 27748 40514
rect 28140 41020 28196 41076
rect 27692 40460 27748 40462
rect 28028 40348 28084 40404
rect 27692 40124 27748 40180
rect 27692 39564 27748 39620
rect 27804 39116 27860 39172
rect 27244 38220 27300 38276
rect 27580 37884 27636 37940
rect 27356 37548 27412 37604
rect 27468 37100 27524 37156
rect 27356 36988 27412 37044
rect 26796 33516 26852 33572
rect 26572 32732 26628 32788
rect 26908 33180 26964 33236
rect 26012 32562 26068 32564
rect 26012 32510 26014 32562
rect 26014 32510 26066 32562
rect 26066 32510 26068 32562
rect 26012 32508 26068 32510
rect 26908 32396 26964 32452
rect 25900 32172 25956 32228
rect 27244 33964 27300 34020
rect 27132 33906 27188 33908
rect 27132 33854 27134 33906
rect 27134 33854 27186 33906
rect 27186 33854 27188 33906
rect 27132 33852 27188 33854
rect 27804 37938 27860 37940
rect 27804 37886 27806 37938
rect 27806 37886 27858 37938
rect 27858 37886 27860 37938
rect 27804 37884 27860 37886
rect 27916 37548 27972 37604
rect 27804 37266 27860 37268
rect 27804 37214 27806 37266
rect 27806 37214 27858 37266
rect 27858 37214 27860 37266
rect 27804 37212 27860 37214
rect 28924 44156 28980 44212
rect 29036 43708 29092 43764
rect 28812 42754 28868 42756
rect 28812 42702 28814 42754
rect 28814 42702 28866 42754
rect 28866 42702 28868 42754
rect 28812 42700 28868 42702
rect 29036 41970 29092 41972
rect 29036 41918 29038 41970
rect 29038 41918 29090 41970
rect 29090 41918 29092 41970
rect 29036 41916 29092 41918
rect 28924 41356 28980 41412
rect 28812 41298 28868 41300
rect 28812 41246 28814 41298
rect 28814 41246 28866 41298
rect 28866 41246 28868 41298
rect 28812 41244 28868 41246
rect 29708 50428 29764 50484
rect 30604 50428 30660 50484
rect 30492 50316 30548 50372
rect 30604 49980 30660 50036
rect 29708 49810 29764 49812
rect 29708 49758 29710 49810
rect 29710 49758 29762 49810
rect 29762 49758 29764 49810
rect 29708 49756 29764 49758
rect 30268 49644 30324 49700
rect 29484 47404 29540 47460
rect 29820 49196 29876 49252
rect 29708 47234 29764 47236
rect 29708 47182 29710 47234
rect 29710 47182 29762 47234
rect 29762 47182 29764 47234
rect 29708 47180 29764 47182
rect 29708 45948 29764 46004
rect 29596 45500 29652 45556
rect 29484 45330 29540 45332
rect 29484 45278 29486 45330
rect 29486 45278 29538 45330
rect 29538 45278 29540 45330
rect 29484 45276 29540 45278
rect 29372 45218 29428 45220
rect 29372 45166 29374 45218
rect 29374 45166 29426 45218
rect 29426 45166 29428 45218
rect 29372 45164 29428 45166
rect 29260 45106 29316 45108
rect 29260 45054 29262 45106
rect 29262 45054 29314 45106
rect 29314 45054 29316 45106
rect 29260 45052 29316 45054
rect 29484 44210 29540 44212
rect 29484 44158 29486 44210
rect 29486 44158 29538 44210
rect 29538 44158 29540 44210
rect 29484 44156 29540 44158
rect 29260 42028 29316 42084
rect 29484 41804 29540 41860
rect 29372 40796 29428 40852
rect 28476 39452 28532 39508
rect 28588 40572 28644 40628
rect 28364 36706 28420 36708
rect 28364 36654 28366 36706
rect 28366 36654 28418 36706
rect 28418 36654 28420 36706
rect 28364 36652 28420 36654
rect 27580 35532 27636 35588
rect 27692 35420 27748 35476
rect 27468 35308 27524 35364
rect 27804 34636 27860 34692
rect 27468 34076 27524 34132
rect 27356 33516 27412 33572
rect 27020 32284 27076 32340
rect 25788 31948 25844 32004
rect 25900 31778 25956 31780
rect 25900 31726 25902 31778
rect 25902 31726 25954 31778
rect 25954 31726 25956 31778
rect 25900 31724 25956 31726
rect 25676 31052 25732 31108
rect 25900 31500 25956 31556
rect 25564 30940 25620 30996
rect 25676 30882 25732 30884
rect 25676 30830 25678 30882
rect 25678 30830 25730 30882
rect 25730 30830 25732 30882
rect 25676 30828 25732 30830
rect 27580 32338 27636 32340
rect 27580 32286 27582 32338
rect 27582 32286 27634 32338
rect 27634 32286 27636 32338
rect 27580 32284 27636 32286
rect 26124 31724 26180 31780
rect 26572 31724 26628 31780
rect 26684 31500 26740 31556
rect 26124 31164 26180 31220
rect 26236 31276 26292 31332
rect 25340 30210 25396 30212
rect 25340 30158 25342 30210
rect 25342 30158 25394 30210
rect 25394 30158 25396 30210
rect 25340 30156 25396 30158
rect 25116 29932 25172 29988
rect 25676 30268 25732 30324
rect 25900 30604 25956 30660
rect 26012 30322 26068 30324
rect 26012 30270 26014 30322
rect 26014 30270 26066 30322
rect 26066 30270 26068 30322
rect 26012 30268 26068 30270
rect 25676 29650 25732 29652
rect 25676 29598 25678 29650
rect 25678 29598 25730 29650
rect 25730 29598 25732 29650
rect 25676 29596 25732 29598
rect 25116 29484 25172 29540
rect 26124 29820 26180 29876
rect 25900 29650 25956 29652
rect 25900 29598 25902 29650
rect 25902 29598 25954 29650
rect 25954 29598 25956 29650
rect 25900 29596 25956 29598
rect 26460 31052 26516 31108
rect 26572 30770 26628 30772
rect 26572 30718 26574 30770
rect 26574 30718 26626 30770
rect 26626 30718 26628 30770
rect 26572 30716 26628 30718
rect 29036 38668 29092 38724
rect 28588 36540 28644 36596
rect 28700 37436 28756 37492
rect 28028 36428 28084 36484
rect 28476 36482 28532 36484
rect 28476 36430 28478 36482
rect 28478 36430 28530 36482
rect 28530 36430 28532 36482
rect 28476 36428 28532 36430
rect 28252 35532 28308 35588
rect 29148 37378 29204 37380
rect 29148 37326 29150 37378
rect 29150 37326 29202 37378
rect 29202 37326 29204 37378
rect 29148 37324 29204 37326
rect 29260 38108 29316 38164
rect 28812 35532 28868 35588
rect 28924 35644 28980 35700
rect 28588 34690 28644 34692
rect 28588 34638 28590 34690
rect 28590 34638 28642 34690
rect 28642 34638 28644 34690
rect 28588 34636 28644 34638
rect 27916 32450 27972 32452
rect 27916 32398 27918 32450
rect 27918 32398 27970 32450
rect 27970 32398 27972 32450
rect 27916 32396 27972 32398
rect 28140 32562 28196 32564
rect 28140 32510 28142 32562
rect 28142 32510 28194 32562
rect 28194 32510 28196 32562
rect 28140 32508 28196 32510
rect 28476 33852 28532 33908
rect 28252 32172 28308 32228
rect 27356 30940 27412 30996
rect 27132 30156 27188 30212
rect 26796 29820 26852 29876
rect 24556 28812 24612 28868
rect 24556 27858 24612 27860
rect 24556 27806 24558 27858
rect 24558 27806 24610 27858
rect 24610 27806 24612 27858
rect 24556 27804 24612 27806
rect 24556 27468 24612 27524
rect 25004 28252 25060 28308
rect 25004 27020 25060 27076
rect 24668 25788 24724 25844
rect 24668 25506 24724 25508
rect 24668 25454 24670 25506
rect 24670 25454 24722 25506
rect 24722 25454 24724 25506
rect 24668 25452 24724 25454
rect 24668 24668 24724 24724
rect 24220 23660 24276 23716
rect 24444 23884 24500 23940
rect 23772 22092 23828 22148
rect 24108 22876 24164 22932
rect 23660 21868 23716 21924
rect 23212 20690 23268 20692
rect 23212 20638 23214 20690
rect 23214 20638 23266 20690
rect 23266 20638 23268 20690
rect 23212 20636 23268 20638
rect 23324 20578 23380 20580
rect 23324 20526 23326 20578
rect 23326 20526 23378 20578
rect 23378 20526 23380 20578
rect 23324 20524 23380 20526
rect 23660 20636 23716 20692
rect 22988 20300 23044 20356
rect 23100 19906 23156 19908
rect 23100 19854 23102 19906
rect 23102 19854 23154 19906
rect 23154 19854 23156 19906
rect 23100 19852 23156 19854
rect 22316 19234 22372 19236
rect 22316 19182 22318 19234
rect 22318 19182 22370 19234
rect 22370 19182 22372 19234
rect 22316 19180 22372 19182
rect 23100 19234 23156 19236
rect 23100 19182 23102 19234
rect 23102 19182 23154 19234
rect 23154 19182 23156 19234
rect 23100 19180 23156 19182
rect 21644 17052 21700 17108
rect 21980 17442 22036 17444
rect 21980 17390 21982 17442
rect 21982 17390 22034 17442
rect 22034 17390 22036 17442
rect 21980 17388 22036 17390
rect 21868 17276 21924 17332
rect 22316 17276 22372 17332
rect 22204 16994 22260 16996
rect 22204 16942 22206 16994
rect 22206 16942 22258 16994
rect 22258 16942 22260 16994
rect 22204 16940 22260 16942
rect 21868 16828 21924 16884
rect 21756 16156 21812 16212
rect 22764 17612 22820 17668
rect 23660 20300 23716 20356
rect 23548 20188 23604 20244
rect 24220 22092 24276 22148
rect 24668 23548 24724 23604
rect 24892 26402 24948 26404
rect 24892 26350 24894 26402
rect 24894 26350 24946 26402
rect 24946 26350 24948 26402
rect 24892 26348 24948 26350
rect 24892 23548 24948 23604
rect 24556 23212 24612 23268
rect 24780 23266 24836 23268
rect 24780 23214 24782 23266
rect 24782 23214 24834 23266
rect 24834 23214 24836 23266
rect 24780 23212 24836 23214
rect 24892 23100 24948 23156
rect 24668 21756 24724 21812
rect 24332 20914 24388 20916
rect 24332 20862 24334 20914
rect 24334 20862 24386 20914
rect 24386 20862 24388 20914
rect 24332 20860 24388 20862
rect 24220 20578 24276 20580
rect 24220 20526 24222 20578
rect 24222 20526 24274 20578
rect 24274 20526 24276 20578
rect 24220 20524 24276 20526
rect 24444 20300 24500 20356
rect 23212 19068 23268 19124
rect 23548 18562 23604 18564
rect 23548 18510 23550 18562
rect 23550 18510 23602 18562
rect 23602 18510 23604 18562
rect 23548 18508 23604 18510
rect 23100 17666 23156 17668
rect 23100 17614 23102 17666
rect 23102 17614 23154 17666
rect 23154 17614 23156 17666
rect 23100 17612 23156 17614
rect 23772 19740 23828 19796
rect 23772 19068 23828 19124
rect 23884 18562 23940 18564
rect 23884 18510 23886 18562
rect 23886 18510 23938 18562
rect 23938 18510 23940 18562
rect 23884 18508 23940 18510
rect 23548 17164 23604 17220
rect 22988 16940 23044 16996
rect 23212 17052 23268 17108
rect 22652 16268 22708 16324
rect 23324 16156 23380 16212
rect 22204 15986 22260 15988
rect 22204 15934 22206 15986
rect 22206 15934 22258 15986
rect 22258 15934 22260 15986
rect 22204 15932 22260 15934
rect 22540 15932 22596 15988
rect 22204 15260 22260 15316
rect 21644 14306 21700 14308
rect 21644 14254 21646 14306
rect 21646 14254 21698 14306
rect 21698 14254 21700 14306
rect 21644 14252 21700 14254
rect 22876 15314 22932 15316
rect 22876 15262 22878 15314
rect 22878 15262 22930 15314
rect 22930 15262 22932 15314
rect 22876 15260 22932 15262
rect 22988 14418 23044 14420
rect 22988 14366 22990 14418
rect 22990 14366 23042 14418
rect 23042 14366 23044 14418
rect 22988 14364 23044 14366
rect 21644 11506 21700 11508
rect 21644 11454 21646 11506
rect 21646 11454 21698 11506
rect 21698 11454 21700 11506
rect 21644 11452 21700 11454
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19628 10722 19684 10724
rect 19628 10670 19630 10722
rect 19630 10670 19682 10722
rect 19682 10670 19684 10722
rect 19628 10668 19684 10670
rect 19964 10610 20020 10612
rect 19964 10558 19966 10610
rect 19966 10558 20018 10610
rect 20018 10558 20020 10610
rect 19964 10556 20020 10558
rect 20524 10610 20580 10612
rect 20524 10558 20526 10610
rect 20526 10558 20578 10610
rect 20578 10558 20580 10610
rect 20524 10556 20580 10558
rect 21196 10610 21252 10612
rect 21196 10558 21198 10610
rect 21198 10558 21250 10610
rect 21250 10558 21252 10610
rect 21196 10556 21252 10558
rect 21420 10498 21476 10500
rect 21420 10446 21422 10498
rect 21422 10446 21474 10498
rect 21474 10446 21476 10498
rect 21420 10444 21476 10446
rect 18956 9714 19012 9716
rect 18956 9662 18958 9714
rect 18958 9662 19010 9714
rect 19010 9662 19012 9714
rect 18956 9660 19012 9662
rect 18396 9602 18452 9604
rect 18396 9550 18398 9602
rect 18398 9550 18450 9602
rect 18450 9550 18452 9602
rect 18396 9548 18452 9550
rect 18732 9548 18788 9604
rect 15484 8988 15540 9044
rect 17052 9042 17108 9044
rect 17052 8990 17054 9042
rect 17054 8990 17106 9042
rect 17106 8990 17108 9042
rect 17052 8988 17108 8990
rect 17612 8988 17668 9044
rect 16492 8652 16548 8708
rect 17612 8428 17668 8484
rect 17948 8540 18004 8596
rect 13244 6130 13300 6132
rect 13244 6078 13246 6130
rect 13246 6078 13298 6130
rect 13298 6078 13300 6130
rect 13244 6076 13300 6078
rect 14476 6636 14532 6692
rect 14028 6076 14084 6132
rect 14364 6130 14420 6132
rect 14364 6078 14366 6130
rect 14366 6078 14418 6130
rect 14418 6078 14420 6130
rect 14364 6076 14420 6078
rect 13804 5516 13860 5572
rect 14252 5628 14308 5684
rect 13132 5404 13188 5460
rect 13580 5234 13636 5236
rect 13580 5182 13582 5234
rect 13582 5182 13634 5234
rect 13634 5182 13636 5234
rect 13580 5180 13636 5182
rect 13020 4956 13076 5012
rect 11228 4060 11284 4116
rect 7644 3500 7700 3556
rect 12908 3442 12964 3444
rect 12908 3390 12910 3442
rect 12910 3390 12962 3442
rect 12962 3390 12964 3442
rect 12908 3388 12964 3390
rect 13692 3442 13748 3444
rect 13692 3390 13694 3442
rect 13694 3390 13746 3442
rect 13746 3390 13748 3442
rect 13692 3388 13748 3390
rect 15372 6524 15428 6580
rect 15708 7980 15764 8036
rect 15708 5906 15764 5908
rect 15708 5854 15710 5906
rect 15710 5854 15762 5906
rect 15762 5854 15764 5906
rect 15708 5852 15764 5854
rect 15484 5180 15540 5236
rect 16044 5292 16100 5348
rect 15372 5122 15428 5124
rect 15372 5070 15374 5122
rect 15374 5070 15426 5122
rect 15426 5070 15428 5122
rect 15372 5068 15428 5070
rect 16716 5906 16772 5908
rect 16716 5854 16718 5906
rect 16718 5854 16770 5906
rect 16770 5854 16772 5906
rect 16716 5852 16772 5854
rect 16604 5628 16660 5684
rect 16380 5180 16436 5236
rect 16604 5180 16660 5236
rect 16828 5068 16884 5124
rect 17612 5068 17668 5124
rect 17948 5852 18004 5908
rect 17724 3554 17780 3556
rect 17724 3502 17726 3554
rect 17726 3502 17778 3554
rect 17778 3502 17780 3554
rect 17724 3500 17780 3502
rect 18620 8652 18676 8708
rect 18732 8540 18788 8596
rect 18620 8258 18676 8260
rect 18620 8206 18622 8258
rect 18622 8206 18674 8258
rect 18674 8206 18676 8258
rect 18620 8204 18676 8206
rect 19292 9548 19348 9604
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 21308 9266 21364 9268
rect 21308 9214 21310 9266
rect 21310 9214 21362 9266
rect 21362 9214 21364 9266
rect 21308 9212 21364 9214
rect 19068 8370 19124 8372
rect 19068 8318 19070 8370
rect 19070 8318 19122 8370
rect 19122 8318 19124 8370
rect 19068 8316 19124 8318
rect 20636 8092 20692 8148
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19628 7420 19684 7476
rect 18732 6914 18788 6916
rect 18732 6862 18734 6914
rect 18734 6862 18786 6914
rect 18786 6862 18788 6914
rect 18732 6860 18788 6862
rect 19628 6860 19684 6916
rect 18060 6076 18116 6132
rect 18060 4844 18116 4900
rect 18172 6412 18228 6468
rect 19404 6466 19460 6468
rect 19404 6414 19406 6466
rect 19406 6414 19458 6466
rect 19458 6414 19460 6466
rect 19404 6412 19460 6414
rect 18284 5906 18340 5908
rect 18284 5854 18286 5906
rect 18286 5854 18338 5906
rect 18338 5854 18340 5906
rect 18284 5852 18340 5854
rect 19068 5122 19124 5124
rect 19068 5070 19070 5122
rect 19070 5070 19122 5122
rect 19122 5070 19124 5122
rect 19068 5068 19124 5070
rect 18284 4898 18340 4900
rect 18284 4846 18286 4898
rect 18286 4846 18338 4898
rect 18338 4846 18340 4898
rect 18284 4844 18340 4846
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 20860 7586 20916 7588
rect 20860 7534 20862 7586
rect 20862 7534 20914 7586
rect 20914 7534 20916 7586
rect 20860 7532 20916 7534
rect 21644 8034 21700 8036
rect 21644 7982 21646 8034
rect 21646 7982 21698 8034
rect 21698 7982 21700 8034
rect 21644 7980 21700 7982
rect 22652 12572 22708 12628
rect 23212 12850 23268 12852
rect 23212 12798 23214 12850
rect 23214 12798 23266 12850
rect 23266 12798 23268 12850
rect 23212 12796 23268 12798
rect 24332 18508 24388 18564
rect 24332 18284 24388 18340
rect 25900 29148 25956 29204
rect 25228 28924 25284 28980
rect 25788 28924 25844 28980
rect 25116 26796 25172 26852
rect 25452 27916 25508 27972
rect 25900 27970 25956 27972
rect 25900 27918 25902 27970
rect 25902 27918 25954 27970
rect 25954 27918 25956 27970
rect 25900 27916 25956 27918
rect 26460 29426 26516 29428
rect 26460 29374 26462 29426
rect 26462 29374 26514 29426
rect 26514 29374 26516 29426
rect 26460 29372 26516 29374
rect 26124 28588 26180 28644
rect 26236 29148 26292 29204
rect 26012 27020 26068 27076
rect 26348 27244 26404 27300
rect 26572 27132 26628 27188
rect 25116 25452 25172 25508
rect 26012 26460 26068 26516
rect 25452 23938 25508 23940
rect 25452 23886 25454 23938
rect 25454 23886 25506 23938
rect 25506 23886 25508 23938
rect 25452 23884 25508 23886
rect 25788 25340 25844 25396
rect 25676 23660 25732 23716
rect 26236 26514 26292 26516
rect 26236 26462 26238 26514
rect 26238 26462 26290 26514
rect 26290 26462 26292 26514
rect 26236 26460 26292 26462
rect 27132 29538 27188 29540
rect 27132 29486 27134 29538
rect 27134 29486 27186 29538
rect 27186 29486 27188 29538
rect 27132 29484 27188 29486
rect 26908 29426 26964 29428
rect 26908 29374 26910 29426
rect 26910 29374 26962 29426
rect 26962 29374 26964 29426
rect 26908 29372 26964 29374
rect 28028 31388 28084 31444
rect 27580 30716 27636 30772
rect 27804 30940 27860 30996
rect 26796 26460 26852 26516
rect 27580 29820 27636 29876
rect 27132 28588 27188 28644
rect 27020 28530 27076 28532
rect 27020 28478 27022 28530
rect 27022 28478 27074 28530
rect 27074 28478 27076 28530
rect 27020 28476 27076 28478
rect 27020 27916 27076 27972
rect 28028 29260 28084 29316
rect 28028 28700 28084 28756
rect 27580 27916 27636 27972
rect 27804 28642 27860 28644
rect 27804 28590 27806 28642
rect 27806 28590 27858 28642
rect 27858 28590 27860 28642
rect 27804 28588 27860 28590
rect 27692 28476 27748 28532
rect 28140 28476 28196 28532
rect 28028 27858 28084 27860
rect 28028 27806 28030 27858
rect 28030 27806 28082 27858
rect 28082 27806 28084 27858
rect 28028 27804 28084 27806
rect 28028 27356 28084 27412
rect 28028 27132 28084 27188
rect 27244 26962 27300 26964
rect 27244 26910 27246 26962
rect 27246 26910 27298 26962
rect 27298 26910 27300 26962
rect 27244 26908 27300 26910
rect 26908 26290 26964 26292
rect 26908 26238 26910 26290
rect 26910 26238 26962 26290
rect 26962 26238 26964 26290
rect 26908 26236 26964 26238
rect 27132 26012 27188 26068
rect 27356 26290 27412 26292
rect 27356 26238 27358 26290
rect 27358 26238 27410 26290
rect 27410 26238 27412 26290
rect 27356 26236 27412 26238
rect 28700 32562 28756 32564
rect 28700 32510 28702 32562
rect 28702 32510 28754 32562
rect 28754 32510 28756 32562
rect 28700 32508 28756 32510
rect 28924 34300 28980 34356
rect 28364 31554 28420 31556
rect 28364 31502 28366 31554
rect 28366 31502 28418 31554
rect 28418 31502 28420 31554
rect 28364 31500 28420 31502
rect 28476 30994 28532 30996
rect 28476 30942 28478 30994
rect 28478 30942 28530 30994
rect 28530 30942 28532 30994
rect 28476 30940 28532 30942
rect 28588 29314 28644 29316
rect 28588 29262 28590 29314
rect 28590 29262 28642 29314
rect 28642 29262 28644 29314
rect 28588 29260 28644 29262
rect 28476 28588 28532 28644
rect 28588 28530 28644 28532
rect 28588 28478 28590 28530
rect 28590 28478 28642 28530
rect 28642 28478 28644 28530
rect 28588 28476 28644 28478
rect 28364 28028 28420 28084
rect 28476 27916 28532 27972
rect 28812 31164 28868 31220
rect 29036 33180 29092 33236
rect 29260 37100 29316 37156
rect 30044 48412 30100 48468
rect 30492 48412 30548 48468
rect 31836 55970 31892 55972
rect 31836 55918 31838 55970
rect 31838 55918 31890 55970
rect 31890 55918 31892 55970
rect 31836 55916 31892 55918
rect 31388 55858 31444 55860
rect 31388 55806 31390 55858
rect 31390 55806 31442 55858
rect 31442 55806 31444 55858
rect 31388 55804 31444 55806
rect 32172 57596 32228 57652
rect 32396 58156 32452 58212
rect 32956 58546 33012 58548
rect 32956 58494 32958 58546
rect 32958 58494 33010 58546
rect 33010 58494 33012 58546
rect 32956 58492 33012 58494
rect 33180 58434 33236 58436
rect 33180 58382 33182 58434
rect 33182 58382 33234 58434
rect 33234 58382 33236 58434
rect 33180 58380 33236 58382
rect 33516 58434 33572 58436
rect 33516 58382 33518 58434
rect 33518 58382 33570 58434
rect 33570 58382 33572 58434
rect 33516 58380 33572 58382
rect 33740 58380 33796 58436
rect 33628 58268 33684 58324
rect 34076 58994 34132 58996
rect 34076 58942 34078 58994
rect 34078 58942 34130 58994
rect 34130 58942 34132 58994
rect 34076 58940 34132 58942
rect 32508 57538 32564 57540
rect 32508 57486 32510 57538
rect 32510 57486 32562 57538
rect 32562 57486 32564 57538
rect 32508 57484 32564 57486
rect 34524 59164 34580 59220
rect 34412 58434 34468 58436
rect 34412 58382 34414 58434
rect 34414 58382 34466 58434
rect 34466 58382 34468 58434
rect 34412 58380 34468 58382
rect 34748 58940 34804 58996
rect 36988 59724 37044 59780
rect 39676 59724 39732 59780
rect 34972 58604 35028 58660
rect 34860 58210 34916 58212
rect 34860 58158 34862 58210
rect 34862 58158 34914 58210
rect 34914 58158 34916 58210
rect 34860 58156 34916 58158
rect 35420 58994 35476 58996
rect 35420 58942 35422 58994
rect 35422 58942 35474 58994
rect 35474 58942 35476 58994
rect 35420 58940 35476 58942
rect 35196 58826 35252 58828
rect 35196 58774 35198 58826
rect 35198 58774 35250 58826
rect 35250 58774 35252 58826
rect 35196 58772 35252 58774
rect 35300 58826 35356 58828
rect 35300 58774 35302 58826
rect 35302 58774 35354 58826
rect 35354 58774 35356 58826
rect 35300 58772 35356 58774
rect 35404 58826 35460 58828
rect 35404 58774 35406 58826
rect 35406 58774 35458 58826
rect 35458 58774 35460 58826
rect 35404 58772 35460 58774
rect 35084 58380 35140 58436
rect 34300 57596 34356 57652
rect 34748 57650 34804 57652
rect 34748 57598 34750 57650
rect 34750 57598 34802 57650
rect 34802 57598 34804 57650
rect 34748 57596 34804 57598
rect 32284 56812 32340 56868
rect 32172 56754 32228 56756
rect 32172 56702 32174 56754
rect 32174 56702 32226 56754
rect 32226 56702 32228 56754
rect 32172 56700 32228 56702
rect 32060 55804 32116 55860
rect 31276 54684 31332 54740
rect 31052 51266 31108 51268
rect 31052 51214 31054 51266
rect 31054 51214 31106 51266
rect 31106 51214 31108 51266
rect 31052 51212 31108 51214
rect 31388 51660 31444 51716
rect 31276 51548 31332 51604
rect 31276 50482 31332 50484
rect 31276 50430 31278 50482
rect 31278 50430 31330 50482
rect 31330 50430 31332 50482
rect 31276 50428 31332 50430
rect 30828 49084 30884 49140
rect 30604 48860 30660 48916
rect 29932 48130 29988 48132
rect 29932 48078 29934 48130
rect 29934 48078 29986 48130
rect 29986 48078 29988 48130
rect 29932 48076 29988 48078
rect 30156 48076 30212 48132
rect 29932 46674 29988 46676
rect 29932 46622 29934 46674
rect 29934 46622 29986 46674
rect 29986 46622 29988 46674
rect 29932 46620 29988 46622
rect 31052 48412 31108 48468
rect 30716 47180 30772 47236
rect 30828 48300 30884 48356
rect 30828 46396 30884 46452
rect 29932 46060 29988 46116
rect 30268 45948 30324 46004
rect 29932 45778 29988 45780
rect 29932 45726 29934 45778
rect 29934 45726 29986 45778
rect 29986 45726 29988 45778
rect 29932 45724 29988 45726
rect 30380 45666 30436 45668
rect 30380 45614 30382 45666
rect 30382 45614 30434 45666
rect 30434 45614 30436 45666
rect 30380 45612 30436 45614
rect 29932 45164 29988 45220
rect 30044 45052 30100 45108
rect 30156 44940 30212 44996
rect 30492 45330 30548 45332
rect 30492 45278 30494 45330
rect 30494 45278 30546 45330
rect 30546 45278 30548 45330
rect 30492 45276 30548 45278
rect 31164 47964 31220 48020
rect 31276 46956 31332 47012
rect 30940 45276 30996 45332
rect 29820 40796 29876 40852
rect 30156 41244 30212 41300
rect 30268 42140 30324 42196
rect 30380 44434 30436 44436
rect 30380 44382 30382 44434
rect 30382 44382 30434 44434
rect 30434 44382 30436 44434
rect 30380 44380 30436 44382
rect 29820 39900 29876 39956
rect 30044 38834 30100 38836
rect 30044 38782 30046 38834
rect 30046 38782 30098 38834
rect 30098 38782 30100 38834
rect 30044 38780 30100 38782
rect 29820 38722 29876 38724
rect 29820 38670 29822 38722
rect 29822 38670 29874 38722
rect 29874 38670 29876 38722
rect 29820 38668 29876 38670
rect 29708 38108 29764 38164
rect 29484 37100 29540 37156
rect 29484 36540 29540 36596
rect 29708 37490 29764 37492
rect 29708 37438 29710 37490
rect 29710 37438 29762 37490
rect 29762 37438 29764 37490
rect 29708 37436 29764 37438
rect 29596 36316 29652 36372
rect 29484 35420 29540 35476
rect 29596 35308 29652 35364
rect 30044 37324 30100 37380
rect 30156 37154 30212 37156
rect 30156 37102 30158 37154
rect 30158 37102 30210 37154
rect 30210 37102 30212 37154
rect 30156 37100 30212 37102
rect 30716 44380 30772 44436
rect 30828 43932 30884 43988
rect 34972 57036 35028 57092
rect 35196 57258 35252 57260
rect 35196 57206 35198 57258
rect 35198 57206 35250 57258
rect 35250 57206 35252 57258
rect 35196 57204 35252 57206
rect 35300 57258 35356 57260
rect 35300 57206 35302 57258
rect 35302 57206 35354 57258
rect 35354 57206 35356 57258
rect 35300 57204 35356 57206
rect 35404 57258 35460 57260
rect 35404 57206 35406 57258
rect 35406 57206 35458 57258
rect 35458 57206 35460 57258
rect 35404 57204 35460 57206
rect 35644 58716 35700 58772
rect 36092 58044 36148 58100
rect 35644 57596 35700 57652
rect 35756 57708 35812 57764
rect 35532 56306 35588 56308
rect 35532 56254 35534 56306
rect 35534 56254 35586 56306
rect 35586 56254 35588 56306
rect 35532 56252 35588 56254
rect 35084 55970 35140 55972
rect 35084 55918 35086 55970
rect 35086 55918 35138 55970
rect 35138 55918 35140 55970
rect 35084 55916 35140 55918
rect 32620 55804 32676 55860
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 36316 57762 36372 57764
rect 36316 57710 36318 57762
rect 36318 57710 36370 57762
rect 36370 57710 36372 57762
rect 36316 57708 36372 57710
rect 38220 59330 38276 59332
rect 38220 59278 38222 59330
rect 38222 59278 38274 59330
rect 38274 59278 38276 59330
rect 38220 59276 38276 59278
rect 39340 59276 39396 59332
rect 36764 59052 36820 59108
rect 38108 59052 38164 59108
rect 37660 58658 37716 58660
rect 37660 58606 37662 58658
rect 37662 58606 37714 58658
rect 37714 58606 37716 58658
rect 37660 58604 37716 58606
rect 36652 58380 36708 58436
rect 37548 58434 37604 58436
rect 37548 58382 37550 58434
rect 37550 58382 37602 58434
rect 37602 58382 37604 58434
rect 37548 58380 37604 58382
rect 39228 58994 39284 58996
rect 39228 58942 39230 58994
rect 39230 58942 39282 58994
rect 39282 58942 39284 58994
rect 39228 58940 39284 58942
rect 38892 58380 38948 58436
rect 39116 58604 39172 58660
rect 37660 58322 37716 58324
rect 37660 58270 37662 58322
rect 37662 58270 37714 58322
rect 37714 58270 37716 58322
rect 37660 58268 37716 58270
rect 38108 58156 38164 58212
rect 38780 58210 38836 58212
rect 38780 58158 38782 58210
rect 38782 58158 38834 58210
rect 38834 58158 38836 58210
rect 38780 58156 38836 58158
rect 39452 58434 39508 58436
rect 39452 58382 39454 58434
rect 39454 58382 39506 58434
rect 39506 58382 39508 58434
rect 39452 58380 39508 58382
rect 36988 57762 37044 57764
rect 36988 57710 36990 57762
rect 36990 57710 37042 57762
rect 37042 57710 37044 57762
rect 36988 57708 37044 57710
rect 36540 57426 36596 57428
rect 36540 57374 36542 57426
rect 36542 57374 36594 57426
rect 36594 57374 36596 57426
rect 36540 57372 36596 57374
rect 36540 57148 36596 57204
rect 35868 57090 35924 57092
rect 35868 57038 35870 57090
rect 35870 57038 35922 57090
rect 35922 57038 35924 57090
rect 35868 57036 35924 57038
rect 36316 57036 36372 57092
rect 35868 56252 35924 56308
rect 32172 55298 32228 55300
rect 32172 55246 32174 55298
rect 32174 55246 32226 55298
rect 32226 55246 32228 55298
rect 32172 55244 32228 55246
rect 32844 55244 32900 55300
rect 32284 54012 32340 54068
rect 32060 50988 32116 51044
rect 31724 49922 31780 49924
rect 31724 49870 31726 49922
rect 31726 49870 31778 49922
rect 31778 49870 31780 49922
rect 31724 49868 31780 49870
rect 31612 48636 31668 48692
rect 31724 47180 31780 47236
rect 31500 45836 31556 45892
rect 31612 46956 31668 47012
rect 31612 46002 31668 46004
rect 31612 45950 31614 46002
rect 31614 45950 31666 46002
rect 31666 45950 31668 46002
rect 31612 45948 31668 45950
rect 31836 45948 31892 46004
rect 31388 45106 31444 45108
rect 31388 45054 31390 45106
rect 31390 45054 31442 45106
rect 31442 45054 31444 45106
rect 31388 45052 31444 45054
rect 31164 43484 31220 43540
rect 31388 44044 31444 44100
rect 30492 43036 30548 43092
rect 31276 43314 31332 43316
rect 31276 43262 31278 43314
rect 31278 43262 31330 43314
rect 31330 43262 31332 43314
rect 31276 43260 31332 43262
rect 30492 42700 30548 42756
rect 30828 42140 30884 42196
rect 31164 42082 31220 42084
rect 31164 42030 31166 42082
rect 31166 42030 31218 42082
rect 31218 42030 31220 42082
rect 31164 42028 31220 42030
rect 30940 41580 30996 41636
rect 30828 40626 30884 40628
rect 30828 40574 30830 40626
rect 30830 40574 30882 40626
rect 30882 40574 30884 40626
rect 30828 40572 30884 40574
rect 30716 38834 30772 38836
rect 30716 38782 30718 38834
rect 30718 38782 30770 38834
rect 30770 38782 30772 38834
rect 30716 38780 30772 38782
rect 30604 38668 30660 38724
rect 30716 37436 30772 37492
rect 31500 42700 31556 42756
rect 32172 50316 32228 50372
rect 32060 46060 32116 46116
rect 32172 46508 32228 46564
rect 32508 54402 32564 54404
rect 32508 54350 32510 54402
rect 32510 54350 32562 54402
rect 32562 54350 32564 54402
rect 32508 54348 32564 54350
rect 32620 54236 32676 54292
rect 33404 55298 33460 55300
rect 33404 55246 33406 55298
rect 33406 55246 33458 55298
rect 33458 55246 33460 55298
rect 33404 55244 33460 55246
rect 33180 55020 33236 55076
rect 32732 53618 32788 53620
rect 32732 53566 32734 53618
rect 32734 53566 32786 53618
rect 32786 53566 32788 53618
rect 32732 53564 32788 53566
rect 33068 52892 33124 52948
rect 32620 51378 32676 51380
rect 32620 51326 32622 51378
rect 32622 51326 32674 51378
rect 32674 51326 32676 51378
rect 32620 51324 32676 51326
rect 32732 51266 32788 51268
rect 32732 51214 32734 51266
rect 32734 51214 32786 51266
rect 32786 51214 32788 51266
rect 32732 51212 32788 51214
rect 32396 50988 32452 51044
rect 33068 50482 33124 50484
rect 33068 50430 33070 50482
rect 33070 50430 33122 50482
rect 33122 50430 33124 50482
rect 33068 50428 33124 50430
rect 34300 55298 34356 55300
rect 34300 55246 34302 55298
rect 34302 55246 34354 55298
rect 34354 55246 34356 55298
rect 34300 55244 34356 55246
rect 35420 55244 35476 55300
rect 35644 55298 35700 55300
rect 35644 55246 35646 55298
rect 35646 55246 35698 55298
rect 35698 55246 35700 55298
rect 35644 55244 35700 55246
rect 33628 54290 33684 54292
rect 33628 54238 33630 54290
rect 33630 54238 33682 54290
rect 33682 54238 33684 54290
rect 33628 54236 33684 54238
rect 33404 53618 33460 53620
rect 33404 53566 33406 53618
rect 33406 53566 33458 53618
rect 33458 53566 33460 53618
rect 33404 53564 33460 53566
rect 34076 54236 34132 54292
rect 33628 52946 33684 52948
rect 33628 52894 33630 52946
rect 33630 52894 33682 52946
rect 33682 52894 33684 52946
rect 33628 52892 33684 52894
rect 33292 52050 33348 52052
rect 33292 51998 33294 52050
rect 33294 51998 33346 52050
rect 33346 51998 33348 52050
rect 33292 51996 33348 51998
rect 33740 51996 33796 52052
rect 33964 51378 34020 51380
rect 33964 51326 33966 51378
rect 33966 51326 34018 51378
rect 34018 51326 34020 51378
rect 33964 51324 34020 51326
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 35084 53618 35140 53620
rect 35084 53566 35086 53618
rect 35086 53566 35138 53618
rect 35138 53566 35140 53618
rect 35084 53564 35140 53566
rect 35196 53506 35252 53508
rect 35196 53454 35198 53506
rect 35198 53454 35250 53506
rect 35250 53454 35252 53506
rect 35196 53452 35252 53454
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 34636 51266 34692 51268
rect 34636 51214 34638 51266
rect 34638 51214 34690 51266
rect 34690 51214 34692 51266
rect 34636 51212 34692 51214
rect 33740 50988 33796 51044
rect 33404 50818 33460 50820
rect 33404 50766 33406 50818
rect 33406 50766 33458 50818
rect 33458 50766 33460 50818
rect 33404 50764 33460 50766
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 34412 50764 34468 50820
rect 34076 50652 34132 50708
rect 32620 50316 32676 50372
rect 32396 49810 32452 49812
rect 32396 49758 32398 49810
rect 32398 49758 32450 49810
rect 32450 49758 32452 49810
rect 32396 49756 32452 49758
rect 32284 46396 32340 46452
rect 32508 49644 32564 49700
rect 32620 49084 32676 49140
rect 32732 48188 32788 48244
rect 32956 48076 33012 48132
rect 32620 46956 32676 47012
rect 32508 46060 32564 46116
rect 33068 45778 33124 45780
rect 33068 45726 33070 45778
rect 33070 45726 33122 45778
rect 33122 45726 33124 45778
rect 33068 45724 33124 45726
rect 32172 45666 32228 45668
rect 32172 45614 32174 45666
rect 32174 45614 32226 45666
rect 32226 45614 32228 45666
rect 32172 45612 32228 45614
rect 32844 45612 32900 45668
rect 32060 45276 32116 45332
rect 32508 44994 32564 44996
rect 32508 44942 32510 44994
rect 32510 44942 32562 44994
rect 32562 44942 32564 44994
rect 32508 44940 32564 44942
rect 32172 43596 32228 43652
rect 31948 43372 32004 43428
rect 31500 38892 31556 38948
rect 31276 38780 31332 38836
rect 30380 36652 30436 36708
rect 30268 36428 30324 36484
rect 30156 36370 30212 36372
rect 30156 36318 30158 36370
rect 30158 36318 30210 36370
rect 30210 36318 30212 36370
rect 30156 36316 30212 36318
rect 30380 35586 30436 35588
rect 30380 35534 30382 35586
rect 30382 35534 30434 35586
rect 30434 35534 30436 35586
rect 30380 35532 30436 35534
rect 30492 35420 30548 35476
rect 30044 34914 30100 34916
rect 30044 34862 30046 34914
rect 30046 34862 30098 34914
rect 30098 34862 30100 34914
rect 30044 34860 30100 34862
rect 29708 34802 29764 34804
rect 29708 34750 29710 34802
rect 29710 34750 29762 34802
rect 29762 34750 29764 34802
rect 29708 34748 29764 34750
rect 28924 29932 28980 29988
rect 28700 27804 28756 27860
rect 28588 27468 28644 27524
rect 28700 27020 28756 27076
rect 28812 26908 28868 26964
rect 27580 26124 27636 26180
rect 26460 25676 26516 25732
rect 27244 25452 27300 25508
rect 26460 25228 26516 25284
rect 26236 24722 26292 24724
rect 26236 24670 26238 24722
rect 26238 24670 26290 24722
rect 26290 24670 26292 24722
rect 26236 24668 26292 24670
rect 25900 24108 25956 24164
rect 26236 24444 26292 24500
rect 26124 23266 26180 23268
rect 26124 23214 26126 23266
rect 26126 23214 26178 23266
rect 26178 23214 26180 23266
rect 26124 23212 26180 23214
rect 25900 22876 25956 22932
rect 26348 23212 26404 23268
rect 25116 21756 25172 21812
rect 25676 21810 25732 21812
rect 25676 21758 25678 21810
rect 25678 21758 25730 21810
rect 25730 21758 25732 21810
rect 25676 21756 25732 21758
rect 24668 20188 24724 20244
rect 26012 22204 26068 22260
rect 26236 22204 26292 22260
rect 26012 20972 26068 21028
rect 25004 20690 25060 20692
rect 25004 20638 25006 20690
rect 25006 20638 25058 20690
rect 25058 20638 25060 20690
rect 25004 20636 25060 20638
rect 25452 20578 25508 20580
rect 25452 20526 25454 20578
rect 25454 20526 25506 20578
rect 25506 20526 25508 20578
rect 25452 20524 25508 20526
rect 26012 20524 26068 20580
rect 25116 20412 25172 20468
rect 24892 19180 24948 19236
rect 24556 19068 24612 19124
rect 24108 16940 24164 16996
rect 24780 18508 24836 18564
rect 25004 18620 25060 18676
rect 25676 19516 25732 19572
rect 25676 19068 25732 19124
rect 25676 18674 25732 18676
rect 25676 18622 25678 18674
rect 25678 18622 25730 18674
rect 25730 18622 25732 18674
rect 25676 18620 25732 18622
rect 25900 18562 25956 18564
rect 25900 18510 25902 18562
rect 25902 18510 25954 18562
rect 25954 18510 25956 18562
rect 25900 18508 25956 18510
rect 25340 17612 25396 17668
rect 25676 17666 25732 17668
rect 25676 17614 25678 17666
rect 25678 17614 25730 17666
rect 25730 17614 25732 17666
rect 25676 17612 25732 17614
rect 25004 17106 25060 17108
rect 25004 17054 25006 17106
rect 25006 17054 25058 17106
rect 25058 17054 25060 17106
rect 25004 17052 25060 17054
rect 24444 16994 24500 16996
rect 24444 16942 24446 16994
rect 24446 16942 24498 16994
rect 24498 16942 24500 16994
rect 24444 16940 24500 16942
rect 23884 16044 23940 16100
rect 23772 15314 23828 15316
rect 23772 15262 23774 15314
rect 23774 15262 23826 15314
rect 23826 15262 23828 15314
rect 23772 15260 23828 15262
rect 24892 16210 24948 16212
rect 24892 16158 24894 16210
rect 24894 16158 24946 16210
rect 24946 16158 24948 16210
rect 24892 16156 24948 16158
rect 24556 15538 24612 15540
rect 24556 15486 24558 15538
rect 24558 15486 24610 15538
rect 24610 15486 24612 15538
rect 24556 15484 24612 15486
rect 24444 15372 24500 15428
rect 24892 15426 24948 15428
rect 24892 15374 24894 15426
rect 24894 15374 24946 15426
rect 24946 15374 24948 15426
rect 24892 15372 24948 15374
rect 24108 15260 24164 15316
rect 23436 13132 23492 13188
rect 23324 12572 23380 12628
rect 22876 12290 22932 12292
rect 22876 12238 22878 12290
rect 22878 12238 22930 12290
rect 22930 12238 22932 12290
rect 22876 12236 22932 12238
rect 23660 12290 23716 12292
rect 23660 12238 23662 12290
rect 23662 12238 23714 12290
rect 23714 12238 23716 12290
rect 23660 12236 23716 12238
rect 22652 11452 22708 11508
rect 23212 11506 23268 11508
rect 23212 11454 23214 11506
rect 23214 11454 23266 11506
rect 23266 11454 23268 11506
rect 23212 11452 23268 11454
rect 22092 10556 22148 10612
rect 22652 10610 22708 10612
rect 22652 10558 22654 10610
rect 22654 10558 22706 10610
rect 22706 10558 22708 10610
rect 22652 10556 22708 10558
rect 21980 10444 22036 10500
rect 22540 10444 22596 10500
rect 21868 9266 21924 9268
rect 21868 9214 21870 9266
rect 21870 9214 21922 9266
rect 21922 9214 21924 9266
rect 21868 9212 21924 9214
rect 23548 10668 23604 10724
rect 22988 10498 23044 10500
rect 22988 10446 22990 10498
rect 22990 10446 23042 10498
rect 23042 10446 23044 10498
rect 22988 10444 23044 10446
rect 23772 10722 23828 10724
rect 23772 10670 23774 10722
rect 23774 10670 23826 10722
rect 23826 10670 23828 10722
rect 23772 10668 23828 10670
rect 23660 10610 23716 10612
rect 23660 10558 23662 10610
rect 23662 10558 23714 10610
rect 23714 10558 23716 10610
rect 23660 10556 23716 10558
rect 23548 9660 23604 9716
rect 23100 9212 23156 9268
rect 21980 8764 22036 8820
rect 22204 7420 22260 7476
rect 22652 8764 22708 8820
rect 23548 9266 23604 9268
rect 23548 9214 23550 9266
rect 23550 9214 23602 9266
rect 23602 9214 23604 9266
rect 23548 9212 23604 9214
rect 23436 8764 23492 8820
rect 22988 7586 23044 7588
rect 22988 7534 22990 7586
rect 22990 7534 23042 7586
rect 23042 7534 23044 7586
rect 22988 7532 23044 7534
rect 22540 7420 22596 7476
rect 23324 8258 23380 8260
rect 23324 8206 23326 8258
rect 23326 8206 23378 8258
rect 23378 8206 23380 8258
rect 23324 8204 23380 8206
rect 23324 7644 23380 7700
rect 23884 8204 23940 8260
rect 23996 8146 24052 8148
rect 23996 8094 23998 8146
rect 23998 8094 24050 8146
rect 24050 8094 24052 8146
rect 23996 8092 24052 8094
rect 21756 6636 21812 6692
rect 22540 6690 22596 6692
rect 22540 6638 22542 6690
rect 22542 6638 22594 6690
rect 22594 6638 22596 6690
rect 22540 6636 22596 6638
rect 20300 6578 20356 6580
rect 20300 6526 20302 6578
rect 20302 6526 20354 6578
rect 20354 6526 20356 6578
rect 20300 6524 20356 6526
rect 21980 6578 22036 6580
rect 21980 6526 21982 6578
rect 21982 6526 22034 6578
rect 22034 6526 22036 6578
rect 21980 6524 22036 6526
rect 20188 5740 20244 5796
rect 19852 5628 19908 5684
rect 20188 5404 20244 5460
rect 20300 5628 20356 5684
rect 20300 5122 20356 5124
rect 20300 5070 20302 5122
rect 20302 5070 20354 5122
rect 20354 5070 20356 5122
rect 20300 5068 20356 5070
rect 23100 6636 23156 6692
rect 22988 6466 23044 6468
rect 22988 6414 22990 6466
rect 22990 6414 23042 6466
rect 23042 6414 23044 6466
rect 22988 6412 23044 6414
rect 22540 6300 22596 6356
rect 21980 5852 22036 5908
rect 23100 5852 23156 5908
rect 23212 6300 23268 6356
rect 21644 5292 21700 5348
rect 21868 5010 21924 5012
rect 21868 4958 21870 5010
rect 21870 4958 21922 5010
rect 21922 4958 21924 5010
rect 21868 4956 21924 4958
rect 22876 5068 22932 5124
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 19628 4508 19684 4564
rect 18172 3666 18228 3668
rect 18172 3614 18174 3666
rect 18174 3614 18226 3666
rect 18226 3614 18228 3666
rect 18172 3612 18228 3614
rect 19628 3666 19684 3668
rect 19628 3614 19630 3666
rect 19630 3614 19682 3666
rect 19682 3614 19684 3666
rect 19628 3612 19684 3614
rect 21756 4508 21812 4564
rect 21308 4338 21364 4340
rect 21308 4286 21310 4338
rect 21310 4286 21362 4338
rect 21362 4286 21364 4338
rect 21308 4284 21364 4286
rect 21532 4284 21588 4340
rect 20748 3612 20804 3668
rect 17948 3500 18004 3556
rect 18620 3554 18676 3556
rect 18620 3502 18622 3554
rect 18622 3502 18674 3554
rect 18674 3502 18676 3554
rect 18620 3500 18676 3502
rect 21308 3554 21364 3556
rect 21308 3502 21310 3554
rect 21310 3502 21362 3554
rect 21362 3502 21364 3554
rect 21308 3500 21364 3502
rect 22204 4338 22260 4340
rect 22204 4286 22206 4338
rect 22206 4286 22258 4338
rect 22258 4286 22260 4338
rect 22204 4284 22260 4286
rect 21644 4172 21700 4228
rect 22652 4226 22708 4228
rect 22652 4174 22654 4226
rect 22654 4174 22706 4226
rect 22706 4174 22708 4226
rect 22652 4172 22708 4174
rect 22092 3666 22148 3668
rect 22092 3614 22094 3666
rect 22094 3614 22146 3666
rect 22146 3614 22148 3666
rect 22092 3612 22148 3614
rect 23436 6466 23492 6468
rect 23436 6414 23438 6466
rect 23438 6414 23490 6466
rect 23490 6414 23492 6466
rect 23436 6412 23492 6414
rect 23212 5068 23268 5124
rect 23548 6300 23604 6356
rect 23996 6300 24052 6356
rect 23548 5852 23604 5908
rect 25676 16770 25732 16772
rect 25676 16718 25678 16770
rect 25678 16718 25730 16770
rect 25730 16718 25732 16770
rect 25676 16716 25732 16718
rect 25676 16156 25732 16212
rect 26012 16828 26068 16884
rect 26348 21586 26404 21588
rect 26348 21534 26350 21586
rect 26350 21534 26402 21586
rect 26402 21534 26404 21586
rect 26348 21532 26404 21534
rect 26796 24050 26852 24052
rect 26796 23998 26798 24050
rect 26798 23998 26850 24050
rect 26850 23998 26852 24050
rect 26796 23996 26852 23998
rect 26796 23772 26852 23828
rect 26572 23378 26628 23380
rect 26572 23326 26574 23378
rect 26574 23326 26626 23378
rect 26626 23326 26628 23378
rect 26572 23324 26628 23326
rect 26684 21420 26740 21476
rect 26908 23436 26964 23492
rect 26908 22988 26964 23044
rect 26908 20524 26964 20580
rect 26796 20412 26852 20468
rect 27468 25900 27524 25956
rect 27580 24834 27636 24836
rect 27580 24782 27582 24834
rect 27582 24782 27634 24834
rect 27634 24782 27636 24834
rect 27580 24780 27636 24782
rect 27356 23436 27412 23492
rect 27356 23212 27412 23268
rect 27468 23154 27524 23156
rect 27468 23102 27470 23154
rect 27470 23102 27522 23154
rect 27522 23102 27524 23154
rect 27468 23100 27524 23102
rect 29372 31164 29428 31220
rect 29260 30156 29316 30212
rect 29148 29538 29204 29540
rect 29148 29486 29150 29538
rect 29150 29486 29202 29538
rect 29202 29486 29204 29538
rect 29148 29484 29204 29486
rect 28476 26178 28532 26180
rect 28476 26126 28478 26178
rect 28478 26126 28530 26178
rect 28530 26126 28532 26178
rect 28476 26124 28532 26126
rect 28364 25900 28420 25956
rect 28476 25452 28532 25508
rect 28252 25004 28308 25060
rect 28028 24444 28084 24500
rect 27580 22204 27636 22260
rect 27916 22258 27972 22260
rect 27916 22206 27918 22258
rect 27918 22206 27970 22258
rect 27970 22206 27972 22258
rect 27916 22204 27972 22206
rect 27468 21644 27524 21700
rect 28588 24498 28644 24500
rect 28588 24446 28590 24498
rect 28590 24446 28642 24498
rect 28642 24446 28644 24498
rect 28588 24444 28644 24446
rect 28476 23884 28532 23940
rect 27132 20972 27188 21028
rect 27356 20802 27412 20804
rect 27356 20750 27358 20802
rect 27358 20750 27410 20802
rect 27410 20750 27412 20802
rect 27356 20748 27412 20750
rect 27132 20690 27188 20692
rect 27132 20638 27134 20690
rect 27134 20638 27186 20690
rect 27186 20638 27188 20690
rect 27132 20636 27188 20638
rect 26908 20300 26964 20356
rect 26460 19740 26516 19796
rect 26348 19516 26404 19572
rect 26460 19180 26516 19236
rect 26572 18956 26628 19012
rect 27244 20300 27300 20356
rect 27244 20130 27300 20132
rect 27244 20078 27246 20130
rect 27246 20078 27298 20130
rect 27298 20078 27300 20130
rect 27244 20076 27300 20078
rect 27020 19180 27076 19236
rect 26572 18620 26628 18676
rect 26348 18450 26404 18452
rect 26348 18398 26350 18450
rect 26350 18398 26402 18450
rect 26402 18398 26404 18450
rect 26348 18396 26404 18398
rect 27244 18956 27300 19012
rect 27020 18674 27076 18676
rect 27020 18622 27022 18674
rect 27022 18622 27074 18674
rect 27074 18622 27076 18674
rect 27020 18620 27076 18622
rect 26908 18562 26964 18564
rect 26908 18510 26910 18562
rect 26910 18510 26962 18562
rect 26962 18510 26964 18562
rect 26908 18508 26964 18510
rect 27468 18508 27524 18564
rect 26124 16716 26180 16772
rect 25900 15484 25956 15540
rect 25676 15314 25732 15316
rect 25676 15262 25678 15314
rect 25678 15262 25730 15314
rect 25730 15262 25732 15314
rect 25676 15260 25732 15262
rect 24220 15036 24276 15092
rect 26236 15538 26292 15540
rect 26236 15486 26238 15538
rect 26238 15486 26290 15538
rect 26290 15486 26292 15538
rect 26236 15484 26292 15486
rect 24220 13468 24276 13524
rect 24780 13692 24836 13748
rect 25564 14364 25620 14420
rect 24892 13468 24948 13524
rect 24780 12850 24836 12852
rect 24780 12798 24782 12850
rect 24782 12798 24834 12850
rect 24834 12798 24836 12850
rect 24780 12796 24836 12798
rect 24220 12348 24276 12404
rect 24332 12290 24388 12292
rect 24332 12238 24334 12290
rect 24334 12238 24386 12290
rect 24386 12238 24388 12290
rect 24332 12236 24388 12238
rect 24444 10892 24500 10948
rect 24780 11170 24836 11172
rect 24780 11118 24782 11170
rect 24782 11118 24834 11170
rect 24834 11118 24836 11170
rect 24780 11116 24836 11118
rect 24332 10498 24388 10500
rect 24332 10446 24334 10498
rect 24334 10446 24386 10498
rect 24386 10446 24388 10498
rect 24332 10444 24388 10446
rect 25004 9884 25060 9940
rect 24668 9212 24724 9268
rect 25116 9212 25172 9268
rect 24668 7586 24724 7588
rect 24668 7534 24670 7586
rect 24670 7534 24722 7586
rect 24722 7534 24724 7586
rect 24668 7532 24724 7534
rect 24892 7980 24948 8036
rect 24220 6412 24276 6468
rect 24220 5964 24276 6020
rect 24444 7474 24500 7476
rect 24444 7422 24446 7474
rect 24446 7422 24498 7474
rect 24498 7422 24500 7474
rect 24444 7420 24500 7422
rect 24668 6690 24724 6692
rect 24668 6638 24670 6690
rect 24670 6638 24722 6690
rect 24722 6638 24724 6690
rect 24668 6636 24724 6638
rect 24780 6524 24836 6580
rect 24108 4844 24164 4900
rect 24556 5292 24612 5348
rect 25452 13468 25508 13524
rect 25340 11394 25396 11396
rect 25340 11342 25342 11394
rect 25342 11342 25394 11394
rect 25394 11342 25396 11394
rect 25340 11340 25396 11342
rect 26124 14364 26180 14420
rect 25900 14306 25956 14308
rect 25900 14254 25902 14306
rect 25902 14254 25954 14306
rect 25954 14254 25956 14306
rect 25900 14252 25956 14254
rect 26124 13468 26180 13524
rect 26572 17500 26628 17556
rect 26684 16882 26740 16884
rect 26684 16830 26686 16882
rect 26686 16830 26738 16882
rect 26738 16830 26740 16882
rect 26684 16828 26740 16830
rect 27132 17612 27188 17668
rect 27020 17052 27076 17108
rect 26908 15484 26964 15540
rect 27020 15596 27076 15652
rect 27020 15372 27076 15428
rect 27580 18450 27636 18452
rect 27580 18398 27582 18450
rect 27582 18398 27634 18450
rect 27634 18398 27636 18450
rect 27580 18396 27636 18398
rect 29148 26124 29204 26180
rect 29148 25564 29204 25620
rect 28812 22146 28868 22148
rect 28812 22094 28814 22146
rect 28814 22094 28866 22146
rect 28866 22094 28868 22146
rect 28812 22092 28868 22094
rect 27804 20972 27860 21028
rect 27804 20130 27860 20132
rect 27804 20078 27806 20130
rect 27806 20078 27858 20130
rect 27858 20078 27860 20130
rect 27804 20076 27860 20078
rect 27804 19516 27860 19572
rect 28700 20972 28756 21028
rect 28140 20300 28196 20356
rect 28028 20130 28084 20132
rect 28028 20078 28030 20130
rect 28030 20078 28082 20130
rect 28082 20078 28084 20130
rect 28028 20076 28084 20078
rect 28028 19852 28084 19908
rect 28364 20578 28420 20580
rect 28364 20526 28366 20578
rect 28366 20526 28418 20578
rect 28418 20526 28420 20578
rect 28364 20524 28420 20526
rect 28364 20300 28420 20356
rect 28588 20802 28644 20804
rect 28588 20750 28590 20802
rect 28590 20750 28642 20802
rect 28642 20750 28644 20802
rect 28588 20748 28644 20750
rect 29932 34076 29988 34132
rect 29820 33852 29876 33908
rect 29596 32508 29652 32564
rect 29932 32396 29988 32452
rect 30380 33740 30436 33796
rect 30380 33180 30436 33236
rect 30156 31052 30212 31108
rect 29596 29986 29652 29988
rect 29596 29934 29598 29986
rect 29598 29934 29650 29986
rect 29650 29934 29652 29986
rect 29596 29932 29652 29934
rect 29820 29596 29876 29652
rect 29932 30716 29988 30772
rect 29820 29314 29876 29316
rect 29820 29262 29822 29314
rect 29822 29262 29874 29314
rect 29874 29262 29876 29314
rect 29820 29260 29876 29262
rect 30156 29484 30212 29540
rect 30044 29260 30100 29316
rect 30044 29036 30100 29092
rect 29372 28082 29428 28084
rect 29372 28030 29374 28082
rect 29374 28030 29426 28082
rect 29426 28030 29428 28082
rect 29372 28028 29428 28030
rect 29484 27244 29540 27300
rect 29484 26402 29540 26404
rect 29484 26350 29486 26402
rect 29486 26350 29538 26402
rect 29538 26350 29540 26402
rect 29484 26348 29540 26350
rect 29372 26236 29428 26292
rect 29148 21810 29204 21812
rect 29148 21758 29150 21810
rect 29150 21758 29202 21810
rect 29202 21758 29204 21810
rect 29148 21756 29204 21758
rect 29260 21644 29316 21700
rect 29372 25900 29428 25956
rect 29708 26290 29764 26292
rect 29708 26238 29710 26290
rect 29710 26238 29762 26290
rect 29762 26238 29764 26290
rect 29708 26236 29764 26238
rect 29596 25900 29652 25956
rect 29932 28530 29988 28532
rect 29932 28478 29934 28530
rect 29934 28478 29986 28530
rect 29986 28478 29988 28530
rect 29932 28476 29988 28478
rect 30828 35810 30884 35812
rect 30828 35758 30830 35810
rect 30830 35758 30882 35810
rect 30882 35758 30884 35810
rect 30828 35756 30884 35758
rect 30604 33852 30660 33908
rect 30828 32508 30884 32564
rect 31052 35644 31108 35700
rect 31052 34914 31108 34916
rect 31052 34862 31054 34914
rect 31054 34862 31106 34914
rect 31106 34862 31108 34914
rect 31052 34860 31108 34862
rect 31500 38722 31556 38724
rect 31500 38670 31502 38722
rect 31502 38670 31554 38722
rect 31554 38670 31556 38722
rect 31500 38668 31556 38670
rect 31388 37548 31444 37604
rect 31276 37100 31332 37156
rect 31276 34972 31332 35028
rect 31164 34748 31220 34804
rect 32956 44994 33012 44996
rect 32956 44942 32958 44994
rect 32958 44942 33010 44994
rect 33010 44942 33012 44994
rect 32956 44940 33012 44942
rect 32956 43372 33012 43428
rect 32508 43314 32564 43316
rect 32508 43262 32510 43314
rect 32510 43262 32562 43314
rect 32562 43262 32564 43314
rect 32508 43260 32564 43262
rect 32844 43314 32900 43316
rect 32844 43262 32846 43314
rect 32846 43262 32898 43314
rect 32898 43262 32900 43314
rect 32844 43260 32900 43262
rect 37436 57036 37492 57092
rect 37548 57372 37604 57428
rect 36428 56754 36484 56756
rect 36428 56702 36430 56754
rect 36430 56702 36482 56754
rect 36482 56702 36484 56754
rect 36428 56700 36484 56702
rect 36316 56252 36372 56308
rect 37212 56588 37268 56644
rect 36092 55916 36148 55972
rect 36316 55186 36372 55188
rect 36316 55134 36318 55186
rect 36318 55134 36370 55186
rect 36370 55134 36372 55186
rect 36316 55132 36372 55134
rect 36092 53564 36148 53620
rect 36652 53452 36708 53508
rect 36540 51548 36596 51604
rect 35868 50652 35924 50708
rect 34076 50092 34132 50148
rect 34188 50428 34244 50484
rect 33852 49980 33908 50036
rect 33964 49868 34020 49924
rect 33628 48748 33684 48804
rect 33852 48748 33908 48804
rect 33292 47068 33348 47124
rect 34300 48412 34356 48468
rect 34412 48300 34468 48356
rect 34076 48242 34132 48244
rect 34076 48190 34078 48242
rect 34078 48190 34130 48242
rect 34130 48190 34132 48242
rect 34076 48188 34132 48190
rect 34076 47458 34132 47460
rect 34076 47406 34078 47458
rect 34078 47406 34130 47458
rect 34130 47406 34132 47458
rect 34076 47404 34132 47406
rect 33964 46172 34020 46228
rect 33516 46060 33572 46116
rect 33740 45948 33796 46004
rect 33180 43932 33236 43988
rect 31948 42754 32004 42756
rect 31948 42702 31950 42754
rect 31950 42702 32002 42754
rect 32002 42702 32004 42754
rect 31948 42700 32004 42702
rect 33292 45666 33348 45668
rect 33292 45614 33294 45666
rect 33294 45614 33346 45666
rect 33346 45614 33348 45666
rect 33292 45612 33348 45614
rect 33628 44994 33684 44996
rect 33628 44942 33630 44994
rect 33630 44942 33682 44994
rect 33682 44942 33684 44994
rect 33628 44940 33684 44942
rect 33292 42924 33348 42980
rect 33516 43426 33572 43428
rect 33516 43374 33518 43426
rect 33518 43374 33570 43426
rect 33570 43374 33572 43426
rect 33516 43372 33572 43374
rect 31724 41858 31780 41860
rect 31724 41806 31726 41858
rect 31726 41806 31778 41858
rect 31778 41806 31780 41858
rect 31724 41804 31780 41806
rect 32284 41692 32340 41748
rect 32508 41804 32564 41860
rect 32284 40796 32340 40852
rect 32284 40626 32340 40628
rect 32284 40574 32286 40626
rect 32286 40574 32338 40626
rect 32338 40574 32340 40626
rect 32284 40572 32340 40574
rect 32396 40348 32452 40404
rect 31724 40290 31780 40292
rect 31724 40238 31726 40290
rect 31726 40238 31778 40290
rect 31778 40238 31780 40290
rect 31724 40236 31780 40238
rect 31836 39900 31892 39956
rect 31724 39340 31780 39396
rect 31612 37772 31668 37828
rect 32172 39618 32228 39620
rect 32172 39566 32174 39618
rect 32174 39566 32226 39618
rect 32226 39566 32228 39618
rect 32172 39564 32228 39566
rect 31836 38668 31892 38724
rect 31724 37436 31780 37492
rect 32060 37884 32116 37940
rect 33068 40348 33124 40404
rect 32844 40236 32900 40292
rect 33516 41692 33572 41748
rect 33292 39340 33348 39396
rect 33404 40796 33460 40852
rect 32620 37826 32676 37828
rect 32620 37774 32622 37826
rect 32622 37774 32674 37826
rect 32674 37774 32676 37826
rect 32620 37772 32676 37774
rect 32396 37436 32452 37492
rect 31836 36988 31892 37044
rect 32172 36988 32228 37044
rect 33628 40908 33684 40964
rect 33516 40572 33572 40628
rect 33516 40236 33572 40292
rect 35308 49756 35364 49812
rect 35980 50204 36036 50260
rect 34636 49698 34692 49700
rect 34636 49646 34638 49698
rect 34638 49646 34690 49698
rect 34690 49646 34692 49698
rect 34636 49644 34692 49646
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 34524 48636 34580 48692
rect 34412 47404 34468 47460
rect 34412 47180 34468 47236
rect 34300 47068 34356 47124
rect 34300 46844 34356 46900
rect 34524 45948 34580 46004
rect 34748 47068 34804 47124
rect 35756 49698 35812 49700
rect 35756 49646 35758 49698
rect 35758 49646 35810 49698
rect 35810 49646 35812 49698
rect 35756 49644 35812 49646
rect 35532 48972 35588 49028
rect 36316 51324 36372 51380
rect 36428 50988 36484 51044
rect 36764 50594 36820 50596
rect 36764 50542 36766 50594
rect 36766 50542 36818 50594
rect 36818 50542 36820 50594
rect 36764 50540 36820 50542
rect 36876 50652 36932 50708
rect 36092 49026 36148 49028
rect 36092 48974 36094 49026
rect 36094 48974 36146 49026
rect 36146 48974 36148 49026
rect 36092 48972 36148 48974
rect 35644 48636 35700 48692
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 35644 46956 35700 47012
rect 35756 46674 35812 46676
rect 35756 46622 35758 46674
rect 35758 46622 35810 46674
rect 35810 46622 35812 46674
rect 35756 46620 35812 46622
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 35868 46562 35924 46564
rect 35868 46510 35870 46562
rect 35870 46510 35922 46562
rect 35922 46510 35924 46562
rect 35868 46508 35924 46510
rect 36540 49698 36596 49700
rect 36540 49646 36542 49698
rect 36542 49646 36594 49698
rect 36594 49646 36596 49698
rect 36540 49644 36596 49646
rect 36764 49644 36820 49700
rect 36428 48242 36484 48244
rect 36428 48190 36430 48242
rect 36430 48190 36482 48242
rect 36482 48190 36484 48242
rect 36428 48188 36484 48190
rect 36540 46956 36596 47012
rect 35532 45666 35588 45668
rect 35532 45614 35534 45666
rect 35534 45614 35586 45666
rect 35586 45614 35588 45666
rect 35532 45612 35588 45614
rect 35756 45612 35812 45668
rect 34860 45500 34916 45556
rect 34748 45388 34804 45444
rect 34636 45330 34692 45332
rect 34636 45278 34638 45330
rect 34638 45278 34690 45330
rect 34690 45278 34692 45330
rect 34636 45276 34692 45278
rect 34412 44716 34468 44772
rect 35084 45106 35140 45108
rect 35084 45054 35086 45106
rect 35086 45054 35138 45106
rect 35138 45054 35140 45106
rect 35084 45052 35140 45054
rect 35532 45052 35588 45108
rect 34860 44940 34916 44996
rect 34748 44156 34804 44212
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 34860 44044 34916 44100
rect 34076 43484 34132 43540
rect 33852 43148 33908 43204
rect 34188 43260 34244 43316
rect 34188 42252 34244 42308
rect 34300 41580 34356 41636
rect 34412 42028 34468 42084
rect 34188 40236 34244 40292
rect 33852 39116 33908 39172
rect 33628 38946 33684 38948
rect 33628 38894 33630 38946
rect 33630 38894 33682 38946
rect 33682 38894 33684 38946
rect 33628 38892 33684 38894
rect 34076 39058 34132 39060
rect 34076 39006 34078 39058
rect 34078 39006 34130 39058
rect 34130 39006 34132 39058
rect 34076 39004 34132 39006
rect 34300 40124 34356 40180
rect 34524 41916 34580 41972
rect 34524 41410 34580 41412
rect 34524 41358 34526 41410
rect 34526 41358 34578 41410
rect 34578 41358 34580 41410
rect 34524 41356 34580 41358
rect 34524 39564 34580 39620
rect 34748 40348 34804 40404
rect 35756 45106 35812 45108
rect 35756 45054 35758 45106
rect 35758 45054 35810 45106
rect 35810 45054 35812 45106
rect 35756 45052 35812 45054
rect 35756 44156 35812 44212
rect 35308 43596 35364 43652
rect 35084 43538 35140 43540
rect 35084 43486 35086 43538
rect 35086 43486 35138 43538
rect 35138 43486 35140 43538
rect 35084 43484 35140 43486
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 36092 45948 36148 46004
rect 35980 44940 36036 44996
rect 36204 45890 36260 45892
rect 36204 45838 36206 45890
rect 36206 45838 36258 45890
rect 36258 45838 36260 45890
rect 36204 45836 36260 45838
rect 37100 48636 37156 48692
rect 36988 47292 37044 47348
rect 36876 46620 36932 46676
rect 36988 46508 37044 46564
rect 36540 46060 36596 46116
rect 36764 45836 36820 45892
rect 36652 45218 36708 45220
rect 36652 45166 36654 45218
rect 36654 45166 36706 45218
rect 36706 45166 36708 45218
rect 36652 45164 36708 45166
rect 36316 44044 36372 44100
rect 35980 43538 36036 43540
rect 35980 43486 35982 43538
rect 35982 43486 36034 43538
rect 36034 43486 36036 43538
rect 35980 43484 36036 43486
rect 35532 42364 35588 42420
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35196 40962 35252 40964
rect 35196 40910 35198 40962
rect 35198 40910 35250 40962
rect 35250 40910 35252 40962
rect 35196 40908 35252 40910
rect 35644 41356 35700 41412
rect 35532 40460 35588 40516
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 34636 39452 34692 39508
rect 34188 38668 34244 38724
rect 34524 39116 34580 39172
rect 34636 39004 34692 39060
rect 34972 39564 35028 39620
rect 33404 38220 33460 38276
rect 33068 37884 33124 37940
rect 32732 36988 32788 37044
rect 32172 36652 32228 36708
rect 31948 36594 32004 36596
rect 31948 36542 31950 36594
rect 31950 36542 32002 36594
rect 32002 36542 32004 36594
rect 31948 36540 32004 36542
rect 31612 35196 31668 35252
rect 31500 34860 31556 34916
rect 32060 36370 32116 36372
rect 32060 36318 32062 36370
rect 32062 36318 32114 36370
rect 32114 36318 32116 36370
rect 32060 36316 32116 36318
rect 31836 35698 31892 35700
rect 31836 35646 31838 35698
rect 31838 35646 31890 35698
rect 31890 35646 31892 35698
rect 31836 35644 31892 35646
rect 32396 36204 32452 36260
rect 32620 36258 32676 36260
rect 32620 36206 32622 36258
rect 32622 36206 32674 36258
rect 32674 36206 32676 36258
rect 32620 36204 32676 36206
rect 32396 35756 32452 35812
rect 32620 35868 32676 35924
rect 32396 34972 32452 35028
rect 31724 34130 31780 34132
rect 31724 34078 31726 34130
rect 31726 34078 31778 34130
rect 31778 34078 31780 34130
rect 31724 34076 31780 34078
rect 32508 34748 32564 34804
rect 32060 34524 32116 34580
rect 30828 31612 30884 31668
rect 31276 33068 31332 33124
rect 30492 31500 30548 31556
rect 30380 30492 30436 30548
rect 30268 29148 30324 29204
rect 30156 28418 30212 28420
rect 30156 28366 30158 28418
rect 30158 28366 30210 28418
rect 30210 28366 30212 28418
rect 30156 28364 30212 28366
rect 30268 27692 30324 27748
rect 29820 25116 29876 25172
rect 29484 24834 29540 24836
rect 29484 24782 29486 24834
rect 29486 24782 29538 24834
rect 29538 24782 29540 24834
rect 29484 24780 29540 24782
rect 29372 22092 29428 22148
rect 29036 20860 29092 20916
rect 29260 20748 29316 20804
rect 28924 20188 28980 20244
rect 28476 20076 28532 20132
rect 27916 18620 27972 18676
rect 27132 15260 27188 15316
rect 27356 16604 27412 16660
rect 27356 15596 27412 15652
rect 26348 13692 26404 13748
rect 26460 13804 26516 13860
rect 26348 13468 26404 13524
rect 26460 13074 26516 13076
rect 26460 13022 26462 13074
rect 26462 13022 26514 13074
rect 26514 13022 26516 13074
rect 26460 13020 26516 13022
rect 26124 11340 26180 11396
rect 25900 11116 25956 11172
rect 26012 11004 26068 11060
rect 25900 10834 25956 10836
rect 25900 10782 25902 10834
rect 25902 10782 25954 10834
rect 25954 10782 25956 10834
rect 25900 10780 25956 10782
rect 25788 9826 25844 9828
rect 25788 9774 25790 9826
rect 25790 9774 25842 9826
rect 25842 9774 25844 9826
rect 25788 9772 25844 9774
rect 25676 9266 25732 9268
rect 25676 9214 25678 9266
rect 25678 9214 25730 9266
rect 25730 9214 25732 9266
rect 25676 9212 25732 9214
rect 26124 10722 26180 10724
rect 26124 10670 26126 10722
rect 26126 10670 26178 10722
rect 26178 10670 26180 10722
rect 26124 10668 26180 10670
rect 26348 11004 26404 11060
rect 27468 15036 27524 15092
rect 26796 14252 26852 14308
rect 27244 14364 27300 14420
rect 26684 13132 26740 13188
rect 27244 14140 27300 14196
rect 27356 14252 27412 14308
rect 27132 11788 27188 11844
rect 26460 10780 26516 10836
rect 26684 10050 26740 10052
rect 26684 9998 26686 10050
rect 26686 9998 26738 10050
rect 26738 9998 26740 10050
rect 26684 9996 26740 9998
rect 27244 11170 27300 11172
rect 27244 11118 27246 11170
rect 27246 11118 27298 11170
rect 27298 11118 27300 11170
rect 27244 11116 27300 11118
rect 27132 10668 27188 10724
rect 27020 9996 27076 10052
rect 27692 14140 27748 14196
rect 27580 13804 27636 13860
rect 27692 13746 27748 13748
rect 27692 13694 27694 13746
rect 27694 13694 27746 13746
rect 27746 13694 27748 13746
rect 27692 13692 27748 13694
rect 27580 12066 27636 12068
rect 27580 12014 27582 12066
rect 27582 12014 27634 12066
rect 27634 12014 27636 12066
rect 27580 12012 27636 12014
rect 28140 17442 28196 17444
rect 28140 17390 28142 17442
rect 28142 17390 28194 17442
rect 28194 17390 28196 17442
rect 28140 17388 28196 17390
rect 28476 18732 28532 18788
rect 28364 18450 28420 18452
rect 28364 18398 28366 18450
rect 28366 18398 28418 18450
rect 28418 18398 28420 18450
rect 28364 18396 28420 18398
rect 28476 17388 28532 17444
rect 28700 20018 28756 20020
rect 28700 19966 28702 20018
rect 28702 19966 28754 20018
rect 28754 19966 28756 20018
rect 28700 19964 28756 19966
rect 28812 19346 28868 19348
rect 28812 19294 28814 19346
rect 28814 19294 28866 19346
rect 28866 19294 28868 19346
rect 28812 19292 28868 19294
rect 28812 18172 28868 18228
rect 28364 17106 28420 17108
rect 28364 17054 28366 17106
rect 28366 17054 28418 17106
rect 28418 17054 28420 17106
rect 28364 17052 28420 17054
rect 28476 16658 28532 16660
rect 28476 16606 28478 16658
rect 28478 16606 28530 16658
rect 28530 16606 28532 16658
rect 28476 16604 28532 16606
rect 28700 17276 28756 17332
rect 28476 15820 28532 15876
rect 28588 15708 28644 15764
rect 28588 15260 28644 15316
rect 27916 14700 27972 14756
rect 28812 16380 28868 16436
rect 28812 15708 28868 15764
rect 28028 13468 28084 13524
rect 28588 15036 28644 15092
rect 29036 18396 29092 18452
rect 29260 19794 29316 19796
rect 29260 19742 29262 19794
rect 29262 19742 29314 19794
rect 29314 19742 29316 19794
rect 29260 19740 29316 19742
rect 29932 24834 29988 24836
rect 29932 24782 29934 24834
rect 29934 24782 29986 24834
rect 29986 24782 29988 24834
rect 29932 24780 29988 24782
rect 29596 23938 29652 23940
rect 29596 23886 29598 23938
rect 29598 23886 29650 23938
rect 29650 23886 29652 23938
rect 29596 23884 29652 23886
rect 30156 26236 30212 26292
rect 31164 31554 31220 31556
rect 31164 31502 31166 31554
rect 31166 31502 31218 31554
rect 31218 31502 31220 31554
rect 31164 31500 31220 31502
rect 30828 30156 30884 30212
rect 30940 30940 30996 30996
rect 30604 29484 30660 29540
rect 30492 28476 30548 28532
rect 30604 29148 30660 29204
rect 30380 27132 30436 27188
rect 30492 28252 30548 28308
rect 30380 25900 30436 25956
rect 30268 25452 30324 25508
rect 30380 25394 30436 25396
rect 30380 25342 30382 25394
rect 30382 25342 30434 25394
rect 30434 25342 30436 25394
rect 30380 25340 30436 25342
rect 30604 27692 30660 27748
rect 30828 29260 30884 29316
rect 30828 28588 30884 28644
rect 31052 30770 31108 30772
rect 31052 30718 31054 30770
rect 31054 30718 31106 30770
rect 31106 30718 31108 30770
rect 31052 30716 31108 30718
rect 31388 32620 31444 32676
rect 31388 31836 31444 31892
rect 31836 33628 31892 33684
rect 32284 33964 32340 34020
rect 31836 31778 31892 31780
rect 31836 31726 31838 31778
rect 31838 31726 31890 31778
rect 31890 31726 31892 31778
rect 31836 31724 31892 31726
rect 31724 31666 31780 31668
rect 31724 31614 31726 31666
rect 31726 31614 31778 31666
rect 31778 31614 31780 31666
rect 31724 31612 31780 31614
rect 31948 31554 32004 31556
rect 31948 31502 31950 31554
rect 31950 31502 32002 31554
rect 32002 31502 32004 31554
rect 31948 31500 32004 31502
rect 32172 33740 32228 33796
rect 31836 30994 31892 30996
rect 31836 30942 31838 30994
rect 31838 30942 31890 30994
rect 31890 30942 31892 30994
rect 31836 30940 31892 30942
rect 30940 28364 30996 28420
rect 31388 29372 31444 29428
rect 30716 27244 30772 27300
rect 30828 27132 30884 27188
rect 30940 27074 30996 27076
rect 30940 27022 30942 27074
rect 30942 27022 30994 27074
rect 30994 27022 30996 27074
rect 30940 27020 30996 27022
rect 31948 29426 32004 29428
rect 31948 29374 31950 29426
rect 31950 29374 32002 29426
rect 32002 29374 32004 29426
rect 31948 29372 32004 29374
rect 31388 28924 31444 28980
rect 31388 28028 31444 28084
rect 31164 27244 31220 27300
rect 31612 27020 31668 27076
rect 32508 33906 32564 33908
rect 32508 33854 32510 33906
rect 32510 33854 32562 33906
rect 32562 33854 32564 33906
rect 32508 33852 32564 33854
rect 32396 33628 32452 33684
rect 32956 36652 33012 36708
rect 32844 36316 32900 36372
rect 32844 34914 32900 34916
rect 32844 34862 32846 34914
rect 32846 34862 32898 34914
rect 32898 34862 32900 34914
rect 32844 34860 32900 34862
rect 32732 33740 32788 33796
rect 32620 33292 32676 33348
rect 32508 32956 32564 33012
rect 32620 32396 32676 32452
rect 32284 31164 32340 31220
rect 32284 28924 32340 28980
rect 31948 26236 32004 26292
rect 31164 25282 31220 25284
rect 31164 25230 31166 25282
rect 31166 25230 31218 25282
rect 31218 25230 31220 25282
rect 31164 25228 31220 25230
rect 31052 25116 31108 25172
rect 30940 23938 30996 23940
rect 30940 23886 30942 23938
rect 30942 23886 30994 23938
rect 30994 23886 30996 23938
rect 30940 23884 30996 23886
rect 30156 23660 30212 23716
rect 30940 23548 30996 23604
rect 30380 23436 30436 23492
rect 30156 22988 30212 23044
rect 30604 23212 30660 23268
rect 30716 23154 30772 23156
rect 30716 23102 30718 23154
rect 30718 23102 30770 23154
rect 30770 23102 30772 23154
rect 30716 23100 30772 23102
rect 30044 21308 30100 21364
rect 30604 22652 30660 22708
rect 30828 22370 30884 22372
rect 30828 22318 30830 22370
rect 30830 22318 30882 22370
rect 30882 22318 30884 22370
rect 30828 22316 30884 22318
rect 30828 21810 30884 21812
rect 30828 21758 30830 21810
rect 30830 21758 30882 21810
rect 30882 21758 30884 21810
rect 30828 21756 30884 21758
rect 30604 21698 30660 21700
rect 30604 21646 30606 21698
rect 30606 21646 30658 21698
rect 30658 21646 30660 21698
rect 30604 21644 30660 21646
rect 30492 21308 30548 21364
rect 29484 19292 29540 19348
rect 29708 20860 29764 20916
rect 29596 19068 29652 19124
rect 29372 18956 29428 19012
rect 29484 18620 29540 18676
rect 29596 18562 29652 18564
rect 29596 18510 29598 18562
rect 29598 18510 29650 18562
rect 29650 18510 29652 18562
rect 29596 18508 29652 18510
rect 29036 16828 29092 16884
rect 29148 17276 29204 17332
rect 28924 15820 28980 15876
rect 29036 16604 29092 16660
rect 28812 14140 28868 14196
rect 29372 17106 29428 17108
rect 29372 17054 29374 17106
rect 29374 17054 29426 17106
rect 29426 17054 29428 17106
rect 29372 17052 29428 17054
rect 29820 20188 29876 20244
rect 30156 19964 30212 20020
rect 29820 19740 29876 19796
rect 30268 19292 30324 19348
rect 30268 18732 30324 18788
rect 29932 18284 29988 18340
rect 30492 18956 30548 19012
rect 31276 24722 31332 24724
rect 31276 24670 31278 24722
rect 31278 24670 31330 24722
rect 31330 24670 31332 24722
rect 31276 24668 31332 24670
rect 32284 28642 32340 28644
rect 32284 28590 32286 28642
rect 32286 28590 32338 28642
rect 32338 28590 32340 28642
rect 32284 28588 32340 28590
rect 32620 31164 32676 31220
rect 32732 31106 32788 31108
rect 32732 31054 32734 31106
rect 32734 31054 32786 31106
rect 32786 31054 32788 31106
rect 32732 31052 32788 31054
rect 32844 30940 32900 30996
rect 32732 30770 32788 30772
rect 32732 30718 32734 30770
rect 32734 30718 32786 30770
rect 32786 30718 32788 30770
rect 32732 30716 32788 30718
rect 32956 30492 33012 30548
rect 32620 28476 32676 28532
rect 32732 28924 32788 28980
rect 32508 28418 32564 28420
rect 32508 28366 32510 28418
rect 32510 28366 32562 28418
rect 32562 28366 32564 28418
rect 32508 28364 32564 28366
rect 32396 28028 32452 28084
rect 33292 37938 33348 37940
rect 33292 37886 33294 37938
rect 33294 37886 33346 37938
rect 33346 37886 33348 37938
rect 33292 37884 33348 37886
rect 33292 37436 33348 37492
rect 33180 34914 33236 34916
rect 33180 34862 33182 34914
rect 33182 34862 33234 34914
rect 33234 34862 33236 34914
rect 33180 34860 33236 34862
rect 33852 38220 33908 38276
rect 33628 37938 33684 37940
rect 33628 37886 33630 37938
rect 33630 37886 33682 37938
rect 33682 37886 33684 37938
rect 33628 37884 33684 37886
rect 33404 36652 33460 36708
rect 33404 35644 33460 35700
rect 33740 37212 33796 37268
rect 33628 35474 33684 35476
rect 33628 35422 33630 35474
rect 33630 35422 33682 35474
rect 33682 35422 33684 35474
rect 33628 35420 33684 35422
rect 33404 33122 33460 33124
rect 33404 33070 33406 33122
rect 33406 33070 33458 33122
rect 33458 33070 33460 33122
rect 33404 33068 33460 33070
rect 33516 35196 33572 35252
rect 33628 34860 33684 34916
rect 34412 38220 34468 38276
rect 34188 38050 34244 38052
rect 34188 37998 34190 38050
rect 34190 37998 34242 38050
rect 34242 37998 34244 38050
rect 34188 37996 34244 37998
rect 34300 37826 34356 37828
rect 34300 37774 34302 37826
rect 34302 37774 34354 37826
rect 34354 37774 34356 37826
rect 34300 37772 34356 37774
rect 34188 37548 34244 37604
rect 34524 37938 34580 37940
rect 34524 37886 34526 37938
rect 34526 37886 34578 37938
rect 34578 37886 34580 37938
rect 34524 37884 34580 37886
rect 34300 36652 34356 36708
rect 33852 35922 33908 35924
rect 33852 35870 33854 35922
rect 33854 35870 33906 35922
rect 33906 35870 33908 35922
rect 33852 35868 33908 35870
rect 33964 35644 34020 35700
rect 33628 32450 33684 32452
rect 33628 32398 33630 32450
rect 33630 32398 33682 32450
rect 33682 32398 33684 32450
rect 33628 32396 33684 32398
rect 33516 32284 33572 32340
rect 33404 32172 33460 32228
rect 33404 31164 33460 31220
rect 33516 31500 33572 31556
rect 33292 30492 33348 30548
rect 32956 28588 33012 28644
rect 33068 29708 33124 29764
rect 32508 27468 32564 27524
rect 32508 27074 32564 27076
rect 32508 27022 32510 27074
rect 32510 27022 32562 27074
rect 32562 27022 32564 27074
rect 32508 27020 32564 27022
rect 32508 26850 32564 26852
rect 32508 26798 32510 26850
rect 32510 26798 32562 26850
rect 32562 26798 32564 26850
rect 32508 26796 32564 26798
rect 32844 28530 32900 28532
rect 32844 28478 32846 28530
rect 32846 28478 32898 28530
rect 32898 28478 32900 28530
rect 32844 28476 32900 28478
rect 33404 29708 33460 29764
rect 33180 28924 33236 28980
rect 32844 27244 32900 27300
rect 31724 24668 31780 24724
rect 31388 24556 31444 24612
rect 31276 23884 31332 23940
rect 31164 22652 31220 22708
rect 30604 18732 30660 18788
rect 30716 19010 30772 19012
rect 30716 18958 30718 19010
rect 30718 18958 30770 19010
rect 30770 18958 30772 19010
rect 30716 18956 30772 18958
rect 30268 17500 30324 17556
rect 29708 16604 29764 16660
rect 29596 16210 29652 16212
rect 29596 16158 29598 16210
rect 29598 16158 29650 16210
rect 29650 16158 29652 16210
rect 29596 16156 29652 16158
rect 29372 15820 29428 15876
rect 29596 15036 29652 15092
rect 29484 14364 29540 14420
rect 28364 12738 28420 12740
rect 28364 12686 28366 12738
rect 28366 12686 28418 12738
rect 28418 12686 28420 12738
rect 28364 12684 28420 12686
rect 29036 12908 29092 12964
rect 28588 12572 28644 12628
rect 28812 12572 28868 12628
rect 29596 14028 29652 14084
rect 29932 14418 29988 14420
rect 29932 14366 29934 14418
rect 29934 14366 29986 14418
rect 29986 14366 29988 14418
rect 29932 14364 29988 14366
rect 30268 15036 30324 15092
rect 30380 16716 30436 16772
rect 30604 18396 30660 18452
rect 30604 17554 30660 17556
rect 30604 17502 30606 17554
rect 30606 17502 30658 17554
rect 30658 17502 30660 17554
rect 30604 17500 30660 17502
rect 30492 16380 30548 16436
rect 30604 16492 30660 16548
rect 30828 17500 30884 17556
rect 30940 19292 30996 19348
rect 31164 19404 31220 19460
rect 31052 18508 31108 18564
rect 31164 18732 31220 18788
rect 32060 25394 32116 25396
rect 32060 25342 32062 25394
rect 32062 25342 32114 25394
rect 32114 25342 32116 25394
rect 32060 25340 32116 25342
rect 32284 25228 32340 25284
rect 32844 27020 32900 27076
rect 33068 28140 33124 28196
rect 31948 25116 32004 25172
rect 32844 25506 32900 25508
rect 32844 25454 32846 25506
rect 32846 25454 32898 25506
rect 32898 25454 32900 25506
rect 32844 25452 32900 25454
rect 32172 25004 32228 25060
rect 32508 25228 32564 25284
rect 32060 24946 32116 24948
rect 32060 24894 32062 24946
rect 32062 24894 32114 24946
rect 32114 24894 32116 24946
rect 32060 24892 32116 24894
rect 31388 22316 31444 22372
rect 31276 18620 31332 18676
rect 31388 20076 31444 20132
rect 31164 17442 31220 17444
rect 31164 17390 31166 17442
rect 31166 17390 31218 17442
rect 31218 17390 31220 17442
rect 31164 17388 31220 17390
rect 31612 21026 31668 21028
rect 31612 20974 31614 21026
rect 31614 20974 31666 21026
rect 31666 20974 31668 21026
rect 31612 20972 31668 20974
rect 33180 28028 33236 28084
rect 33180 25618 33236 25620
rect 33180 25566 33182 25618
rect 33182 25566 33234 25618
rect 33234 25566 33236 25618
rect 33180 25564 33236 25566
rect 33068 25452 33124 25508
rect 32956 25116 33012 25172
rect 32396 23996 32452 24052
rect 32060 23436 32116 23492
rect 32172 23266 32228 23268
rect 32172 23214 32174 23266
rect 32174 23214 32226 23266
rect 32226 23214 32228 23266
rect 32172 23212 32228 23214
rect 32060 22428 32116 22484
rect 32396 23660 32452 23716
rect 32396 23436 32452 23492
rect 32284 22764 32340 22820
rect 32172 21756 32228 21812
rect 31948 21644 32004 21700
rect 31836 20412 31892 20468
rect 31836 20076 31892 20132
rect 31724 20018 31780 20020
rect 31724 19966 31726 20018
rect 31726 19966 31778 20018
rect 31778 19966 31780 20018
rect 31724 19964 31780 19966
rect 32060 19740 32116 19796
rect 32732 25004 32788 25060
rect 32732 23324 32788 23380
rect 32844 24780 32900 24836
rect 32620 22876 32676 22932
rect 32844 22764 32900 22820
rect 33740 31164 33796 31220
rect 33628 30210 33684 30212
rect 33628 30158 33630 30210
rect 33630 30158 33682 30210
rect 33682 30158 33684 30210
rect 33628 30156 33684 30158
rect 34524 35868 34580 35924
rect 34636 35698 34692 35700
rect 34636 35646 34638 35698
rect 34638 35646 34690 35698
rect 34690 35646 34692 35698
rect 34636 35644 34692 35646
rect 34524 34914 34580 34916
rect 34524 34862 34526 34914
rect 34526 34862 34578 34914
rect 34578 34862 34580 34914
rect 34524 34860 34580 34862
rect 34300 34412 34356 34468
rect 34524 34636 34580 34692
rect 34076 32060 34132 32116
rect 35868 41970 35924 41972
rect 35868 41918 35870 41970
rect 35870 41918 35922 41970
rect 35922 41918 35924 41970
rect 35868 41916 35924 41918
rect 35980 41186 36036 41188
rect 35980 41134 35982 41186
rect 35982 41134 36034 41186
rect 36034 41134 36036 41186
rect 35980 41132 36036 41134
rect 35980 40626 36036 40628
rect 35980 40574 35982 40626
rect 35982 40574 36034 40626
rect 36034 40574 36036 40626
rect 35980 40572 36036 40574
rect 36204 43596 36260 43652
rect 36092 40236 36148 40292
rect 36204 42700 36260 42756
rect 36652 42700 36708 42756
rect 36428 42476 36484 42532
rect 36540 42082 36596 42084
rect 36540 42030 36542 42082
rect 36542 42030 36594 42082
rect 36594 42030 36596 42082
rect 36540 42028 36596 42030
rect 36428 41244 36484 41300
rect 36876 45612 36932 45668
rect 37100 45724 37156 45780
rect 36876 41692 36932 41748
rect 37100 45500 37156 45556
rect 36316 40684 36372 40740
rect 36092 39618 36148 39620
rect 36092 39566 36094 39618
rect 36094 39566 36146 39618
rect 36146 39566 36148 39618
rect 36092 39564 36148 39566
rect 35868 39506 35924 39508
rect 35868 39454 35870 39506
rect 35870 39454 35922 39506
rect 35922 39454 35924 39506
rect 35868 39452 35924 39454
rect 37100 41356 37156 41412
rect 36428 40236 36484 40292
rect 36428 40012 36484 40068
rect 36652 40236 36708 40292
rect 36988 40908 37044 40964
rect 36540 39004 36596 39060
rect 34972 37884 35028 37940
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35196 37884 35252 37940
rect 35308 37548 35364 37604
rect 35084 37212 35140 37268
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 36316 38162 36372 38164
rect 36316 38110 36318 38162
rect 36318 38110 36370 38162
rect 36370 38110 36372 38162
rect 36316 38108 36372 38110
rect 36204 37772 36260 37828
rect 36540 37772 36596 37828
rect 36204 36988 36260 37044
rect 34860 36428 34916 36484
rect 35308 36482 35364 36484
rect 35308 36430 35310 36482
rect 35310 36430 35362 36482
rect 35362 36430 35364 36482
rect 35308 36428 35364 36430
rect 35980 36258 36036 36260
rect 35980 36206 35982 36258
rect 35982 36206 36034 36258
rect 36034 36206 36036 36258
rect 35980 36204 36036 36206
rect 35756 35980 35812 36036
rect 34972 35922 35028 35924
rect 34972 35870 34974 35922
rect 34974 35870 35026 35922
rect 35026 35870 35028 35922
rect 34972 35868 35028 35870
rect 36428 36652 36484 36708
rect 36652 36204 36708 36260
rect 35084 35532 35140 35588
rect 34860 34860 34916 34916
rect 34076 31052 34132 31108
rect 34860 34412 34916 34468
rect 35532 35420 35588 35476
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35084 34636 35140 34692
rect 35196 34412 35252 34468
rect 35084 34076 35140 34132
rect 34412 32172 34468 32228
rect 34524 32284 34580 32340
rect 34412 31778 34468 31780
rect 34412 31726 34414 31778
rect 34414 31726 34466 31778
rect 34466 31726 34468 31778
rect 34412 31724 34468 31726
rect 34300 30828 34356 30884
rect 34300 30156 34356 30212
rect 33628 29538 33684 29540
rect 33628 29486 33630 29538
rect 33630 29486 33682 29538
rect 33682 29486 33684 29538
rect 33628 29484 33684 29486
rect 33852 29708 33908 29764
rect 33852 28700 33908 28756
rect 33852 28028 33908 28084
rect 33852 27356 33908 27412
rect 33292 25340 33348 25396
rect 33852 27020 33908 27076
rect 33740 26290 33796 26292
rect 33740 26238 33742 26290
rect 33742 26238 33794 26290
rect 33794 26238 33796 26290
rect 33740 26236 33796 26238
rect 33404 23212 33460 23268
rect 33516 25452 33572 25508
rect 34188 28252 34244 28308
rect 34188 28082 34244 28084
rect 34188 28030 34190 28082
rect 34190 28030 34242 28082
rect 34242 28030 34244 28082
rect 34188 28028 34244 28030
rect 34524 30044 34580 30100
rect 34636 32060 34692 32116
rect 34972 31612 35028 31668
rect 34972 30492 35028 30548
rect 34748 30380 34804 30436
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35756 35308 35812 35364
rect 35868 34914 35924 34916
rect 35868 34862 35870 34914
rect 35870 34862 35922 34914
rect 35922 34862 35924 34914
rect 35868 34860 35924 34862
rect 35756 34130 35812 34132
rect 35756 34078 35758 34130
rect 35758 34078 35810 34130
rect 35810 34078 35812 34130
rect 35756 34076 35812 34078
rect 36204 35586 36260 35588
rect 36204 35534 36206 35586
rect 36206 35534 36258 35586
rect 36258 35534 36260 35586
rect 36204 35532 36260 35534
rect 36876 38556 36932 38612
rect 36876 37100 36932 37156
rect 36876 35980 36932 36036
rect 37100 39058 37156 39060
rect 37100 39006 37102 39058
rect 37102 39006 37154 39058
rect 37154 39006 37156 39058
rect 37100 39004 37156 39006
rect 37100 38668 37156 38724
rect 37100 35586 37156 35588
rect 37100 35534 37102 35586
rect 37102 35534 37154 35586
rect 37154 35534 37156 35586
rect 37100 35532 37156 35534
rect 36988 35420 37044 35476
rect 36764 35084 36820 35140
rect 36092 34802 36148 34804
rect 36092 34750 36094 34802
rect 36094 34750 36146 34802
rect 36146 34750 36148 34802
rect 36092 34748 36148 34750
rect 36652 34354 36708 34356
rect 36652 34302 36654 34354
rect 36654 34302 36706 34354
rect 36706 34302 36708 34354
rect 36652 34300 36708 34302
rect 36204 34188 36260 34244
rect 36764 34076 36820 34132
rect 35980 33346 36036 33348
rect 35980 33294 35982 33346
rect 35982 33294 36034 33346
rect 36034 33294 36036 33346
rect 35980 33292 36036 33294
rect 36316 33234 36372 33236
rect 36316 33182 36318 33234
rect 36318 33182 36370 33234
rect 36370 33182 36372 33234
rect 36316 33180 36372 33182
rect 36428 33122 36484 33124
rect 36428 33070 36430 33122
rect 36430 33070 36482 33122
rect 36482 33070 36484 33122
rect 36428 33068 36484 33070
rect 35532 32732 35588 32788
rect 35308 32562 35364 32564
rect 35308 32510 35310 32562
rect 35310 32510 35362 32562
rect 35362 32510 35364 32562
rect 35308 32508 35364 32510
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35532 31948 35588 32004
rect 35644 32396 35700 32452
rect 35196 31836 35252 31892
rect 35644 30716 35700 30772
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 34636 29932 34692 29988
rect 34972 29650 35028 29652
rect 34972 29598 34974 29650
rect 34974 29598 35026 29650
rect 35026 29598 35028 29650
rect 34972 29596 35028 29598
rect 35084 29708 35140 29764
rect 34524 29036 34580 29092
rect 34524 28700 34580 28756
rect 34972 29372 35028 29428
rect 34748 28924 34804 28980
rect 34636 28476 34692 28532
rect 33964 26684 34020 26740
rect 33964 26402 34020 26404
rect 33964 26350 33966 26402
rect 33966 26350 34018 26402
rect 34018 26350 34020 26402
rect 33964 26348 34020 26350
rect 33964 25618 34020 25620
rect 33964 25566 33966 25618
rect 33966 25566 34018 25618
rect 34018 25566 34020 25618
rect 33964 25564 34020 25566
rect 34748 27692 34804 27748
rect 34748 27132 34804 27188
rect 34300 25564 34356 25620
rect 34412 26908 34468 26964
rect 33964 25116 34020 25172
rect 34300 25116 34356 25172
rect 34188 24722 34244 24724
rect 34188 24670 34190 24722
rect 34190 24670 34242 24722
rect 34242 24670 34244 24722
rect 34188 24668 34244 24670
rect 34076 23660 34132 23716
rect 32732 22092 32788 22148
rect 32284 19964 32340 20020
rect 31612 19010 31668 19012
rect 31612 18958 31614 19010
rect 31614 18958 31666 19010
rect 31666 18958 31668 19010
rect 31612 18956 31668 18958
rect 31500 18732 31556 18788
rect 31612 18620 31668 18676
rect 31500 18450 31556 18452
rect 31500 18398 31502 18450
rect 31502 18398 31554 18450
rect 31554 18398 31556 18450
rect 31500 18396 31556 18398
rect 31500 17388 31556 17444
rect 32060 18732 32116 18788
rect 32172 18562 32228 18564
rect 32172 18510 32174 18562
rect 32174 18510 32226 18562
rect 32226 18510 32228 18562
rect 32172 18508 32228 18510
rect 31724 17612 31780 17668
rect 31836 18172 31892 18228
rect 30716 16156 30772 16212
rect 30156 14754 30212 14756
rect 30156 14702 30158 14754
rect 30158 14702 30210 14754
rect 30210 14702 30212 14754
rect 30156 14700 30212 14702
rect 31276 16044 31332 16100
rect 31052 15708 31108 15764
rect 30828 15036 30884 15092
rect 30380 14364 30436 14420
rect 30492 14588 30548 14644
rect 29484 12572 29540 12628
rect 28588 12012 28644 12068
rect 29820 12962 29876 12964
rect 29820 12910 29822 12962
rect 29822 12910 29874 12962
rect 29874 12910 29876 12962
rect 29820 12908 29876 12910
rect 28364 11506 28420 11508
rect 28364 11454 28366 11506
rect 28366 11454 28418 11506
rect 28418 11454 28420 11506
rect 28364 11452 28420 11454
rect 27804 11004 27860 11060
rect 26908 9826 26964 9828
rect 26908 9774 26910 9826
rect 26910 9774 26962 9826
rect 26962 9774 26964 9826
rect 26908 9772 26964 9774
rect 26908 9548 26964 9604
rect 27132 9660 27188 9716
rect 25676 7980 25732 8036
rect 26012 8316 26068 8372
rect 25788 7586 25844 7588
rect 25788 7534 25790 7586
rect 25790 7534 25842 7586
rect 25842 7534 25844 7586
rect 25788 7532 25844 7534
rect 25788 6690 25844 6692
rect 25788 6638 25790 6690
rect 25790 6638 25842 6690
rect 25842 6638 25844 6690
rect 25788 6636 25844 6638
rect 25452 6466 25508 6468
rect 25452 6414 25454 6466
rect 25454 6414 25506 6466
rect 25506 6414 25508 6466
rect 25452 6412 25508 6414
rect 27692 9714 27748 9716
rect 27692 9662 27694 9714
rect 27694 9662 27746 9714
rect 27746 9662 27748 9714
rect 27692 9660 27748 9662
rect 27468 9602 27524 9604
rect 27468 9550 27470 9602
rect 27470 9550 27522 9602
rect 27522 9550 27524 9602
rect 27468 9548 27524 9550
rect 27580 9042 27636 9044
rect 27580 8990 27582 9042
rect 27582 8990 27634 9042
rect 27634 8990 27636 9042
rect 27580 8988 27636 8990
rect 28028 11116 28084 11172
rect 28924 11170 28980 11172
rect 28924 11118 28926 11170
rect 28926 11118 28978 11170
rect 28978 11118 28980 11170
rect 28924 11116 28980 11118
rect 27916 9548 27972 9604
rect 28588 9938 28644 9940
rect 28588 9886 28590 9938
rect 28590 9886 28642 9938
rect 28642 9886 28644 9938
rect 28588 9884 28644 9886
rect 28476 9714 28532 9716
rect 28476 9662 28478 9714
rect 28478 9662 28530 9714
rect 28530 9662 28532 9714
rect 28476 9660 28532 9662
rect 28140 8818 28196 8820
rect 28140 8766 28142 8818
rect 28142 8766 28194 8818
rect 28194 8766 28196 8818
rect 28140 8764 28196 8766
rect 27244 8034 27300 8036
rect 27244 7982 27246 8034
rect 27246 7982 27298 8034
rect 27298 7982 27300 8034
rect 27244 7980 27300 7982
rect 27132 7756 27188 7812
rect 26684 7644 26740 7700
rect 27468 7698 27524 7700
rect 27468 7646 27470 7698
rect 27470 7646 27522 7698
rect 27522 7646 27524 7698
rect 27468 7644 27524 7646
rect 27692 7644 27748 7700
rect 27356 7586 27412 7588
rect 27356 7534 27358 7586
rect 27358 7534 27410 7586
rect 27410 7534 27412 7586
rect 27356 7532 27412 7534
rect 26796 7196 26852 7252
rect 28700 9602 28756 9604
rect 28700 9550 28702 9602
rect 28702 9550 28754 9602
rect 28754 9550 28756 9602
rect 28700 9548 28756 9550
rect 30156 12850 30212 12852
rect 30156 12798 30158 12850
rect 30158 12798 30210 12850
rect 30210 12798 30212 12850
rect 30156 12796 30212 12798
rect 29932 11116 29988 11172
rect 30044 12684 30100 12740
rect 31388 15538 31444 15540
rect 31388 15486 31390 15538
rect 31390 15486 31442 15538
rect 31442 15486 31444 15538
rect 31388 15484 31444 15486
rect 31388 15260 31444 15316
rect 31836 17164 31892 17220
rect 32508 20860 32564 20916
rect 32508 19794 32564 19796
rect 32508 19742 32510 19794
rect 32510 19742 32562 19794
rect 32562 19742 32564 19794
rect 32508 19740 32564 19742
rect 33068 22092 33124 22148
rect 32732 21698 32788 21700
rect 32732 21646 32734 21698
rect 32734 21646 32786 21698
rect 32786 21646 32788 21698
rect 32732 21644 32788 21646
rect 32956 21532 33012 21588
rect 32732 20188 32788 20244
rect 32956 20076 33012 20132
rect 32844 19964 32900 20020
rect 32396 19292 32452 19348
rect 33740 22764 33796 22820
rect 33292 21868 33348 21924
rect 32732 18338 32788 18340
rect 32732 18286 32734 18338
rect 32734 18286 32786 18338
rect 32786 18286 32788 18338
rect 32732 18284 32788 18286
rect 32284 18172 32340 18228
rect 32284 17612 32340 17668
rect 32620 17612 32676 17668
rect 32732 17554 32788 17556
rect 32732 17502 32734 17554
rect 32734 17502 32786 17554
rect 32786 17502 32788 17554
rect 32732 17500 32788 17502
rect 32396 16156 32452 16212
rect 32172 15708 32228 15764
rect 32732 16210 32788 16212
rect 32732 16158 32734 16210
rect 32734 16158 32786 16210
rect 32786 16158 32788 16210
rect 32732 16156 32788 16158
rect 33068 18844 33124 18900
rect 32956 16882 33012 16884
rect 32956 16830 32958 16882
rect 32958 16830 33010 16882
rect 33010 16830 33012 16882
rect 32956 16828 33012 16830
rect 33404 20412 33460 20468
rect 33852 22370 33908 22372
rect 33852 22318 33854 22370
rect 33854 22318 33906 22370
rect 33906 22318 33908 22370
rect 33852 22316 33908 22318
rect 34188 22876 34244 22932
rect 33740 21644 33796 21700
rect 33516 20188 33572 20244
rect 33628 20802 33684 20804
rect 33628 20750 33630 20802
rect 33630 20750 33682 20802
rect 33682 20750 33684 20802
rect 33628 20748 33684 20750
rect 33516 18674 33572 18676
rect 33516 18622 33518 18674
rect 33518 18622 33570 18674
rect 33570 18622 33572 18674
rect 33516 18620 33572 18622
rect 33628 18396 33684 18452
rect 33292 18284 33348 18340
rect 33068 16156 33124 16212
rect 33180 17500 33236 17556
rect 33180 16940 33236 16996
rect 32844 15932 32900 15988
rect 32620 15372 32676 15428
rect 31724 15036 31780 15092
rect 31500 14476 31556 14532
rect 32172 15260 32228 15316
rect 31500 13970 31556 13972
rect 31500 13918 31502 13970
rect 31502 13918 31554 13970
rect 31554 13918 31556 13970
rect 31500 13916 31556 13918
rect 30828 13858 30884 13860
rect 30828 13806 30830 13858
rect 30830 13806 30882 13858
rect 30882 13806 30884 13858
rect 30828 13804 30884 13806
rect 31164 13692 31220 13748
rect 30716 12850 30772 12852
rect 30716 12798 30718 12850
rect 30718 12798 30770 12850
rect 30770 12798 30772 12850
rect 30716 12796 30772 12798
rect 29596 9884 29652 9940
rect 29708 9602 29764 9604
rect 29708 9550 29710 9602
rect 29710 9550 29762 9602
rect 29762 9550 29764 9602
rect 29708 9548 29764 9550
rect 28588 8428 28644 8484
rect 28476 8316 28532 8372
rect 28252 7586 28308 7588
rect 28252 7534 28254 7586
rect 28254 7534 28306 7586
rect 28306 7534 28308 7586
rect 28252 7532 28308 7534
rect 28812 8146 28868 8148
rect 28812 8094 28814 8146
rect 28814 8094 28866 8146
rect 28866 8094 28868 8146
rect 28812 8092 28868 8094
rect 26348 6412 26404 6468
rect 26012 6130 26068 6132
rect 26012 6078 26014 6130
rect 26014 6078 26066 6130
rect 26066 6078 26068 6130
rect 26012 6076 26068 6078
rect 25900 5964 25956 6020
rect 26572 6076 26628 6132
rect 27020 6524 27076 6580
rect 27580 6578 27636 6580
rect 27580 6526 27582 6578
rect 27582 6526 27634 6578
rect 27634 6526 27636 6578
rect 27580 6524 27636 6526
rect 26460 6018 26516 6020
rect 26460 5966 26462 6018
rect 26462 5966 26514 6018
rect 26514 5966 26516 6018
rect 26460 5964 26516 5966
rect 26236 5628 26292 5684
rect 25900 5404 25956 5460
rect 24668 4956 24724 5012
rect 24668 4508 24724 4564
rect 25004 4844 25060 4900
rect 25452 5122 25508 5124
rect 25452 5070 25454 5122
rect 25454 5070 25506 5122
rect 25506 5070 25508 5122
rect 25452 5068 25508 5070
rect 25788 4562 25844 4564
rect 25788 4510 25790 4562
rect 25790 4510 25842 4562
rect 25842 4510 25844 4562
rect 25788 4508 25844 4510
rect 24220 3666 24276 3668
rect 24220 3614 24222 3666
rect 24222 3614 24274 3666
rect 24274 3614 24276 3666
rect 24220 3612 24276 3614
rect 24668 3666 24724 3668
rect 24668 3614 24670 3666
rect 24670 3614 24722 3666
rect 24722 3614 24724 3666
rect 24668 3612 24724 3614
rect 25564 3612 25620 3668
rect 26012 5068 26068 5124
rect 26348 5404 26404 5460
rect 26908 5628 26964 5684
rect 27580 5682 27636 5684
rect 27580 5630 27582 5682
rect 27582 5630 27634 5682
rect 27634 5630 27636 5682
rect 27580 5628 27636 5630
rect 27020 5404 27076 5460
rect 27468 5404 27524 5460
rect 27132 5292 27188 5348
rect 26460 4284 26516 4340
rect 26796 4284 26852 4340
rect 26348 4060 26404 4116
rect 26908 4226 26964 4228
rect 26908 4174 26910 4226
rect 26910 4174 26962 4226
rect 26962 4174 26964 4226
rect 26908 4172 26964 4174
rect 30156 12236 30212 12292
rect 30492 12290 30548 12292
rect 30492 12238 30494 12290
rect 30494 12238 30546 12290
rect 30546 12238 30548 12290
rect 30492 12236 30548 12238
rect 31500 13692 31556 13748
rect 30940 12348 30996 12404
rect 30268 11452 30324 11508
rect 30380 12012 30436 12068
rect 30156 10332 30212 10388
rect 30268 9548 30324 9604
rect 29932 8988 29988 9044
rect 29148 8930 29204 8932
rect 29148 8878 29150 8930
rect 29150 8878 29202 8930
rect 29202 8878 29204 8930
rect 29148 8876 29204 8878
rect 28924 7980 28980 8036
rect 29036 8428 29092 8484
rect 28812 7196 28868 7252
rect 28028 6636 28084 6692
rect 28588 6690 28644 6692
rect 28588 6638 28590 6690
rect 28590 6638 28642 6690
rect 28642 6638 28644 6690
rect 28588 6636 28644 6638
rect 27804 5292 27860 5348
rect 28476 5404 28532 5460
rect 27692 5068 27748 5124
rect 27580 4844 27636 4900
rect 28252 4732 28308 4788
rect 28476 4396 28532 4452
rect 28364 4338 28420 4340
rect 28364 4286 28366 4338
rect 28366 4286 28418 4338
rect 28418 4286 28420 4338
rect 28364 4284 28420 4286
rect 28140 4226 28196 4228
rect 28140 4174 28142 4226
rect 28142 4174 28194 4226
rect 28194 4174 28196 4226
rect 28140 4172 28196 4174
rect 28140 3554 28196 3556
rect 28140 3502 28142 3554
rect 28142 3502 28194 3554
rect 28194 3502 28196 3554
rect 28140 3500 28196 3502
rect 29932 8428 29988 8484
rect 29708 8316 29764 8372
rect 29708 8034 29764 8036
rect 29708 7982 29710 8034
rect 29710 7982 29762 8034
rect 29762 7982 29764 8034
rect 29708 7980 29764 7982
rect 29820 7644 29876 7700
rect 30268 8316 30324 8372
rect 30268 7644 30324 7700
rect 30604 11564 30660 11620
rect 30828 11452 30884 11508
rect 30492 11394 30548 11396
rect 30492 11342 30494 11394
rect 30494 11342 30546 11394
rect 30546 11342 30548 11394
rect 30492 11340 30548 11342
rect 30716 9548 30772 9604
rect 30380 7420 30436 7476
rect 30492 8034 30548 8036
rect 30492 7982 30494 8034
rect 30494 7982 30546 8034
rect 30546 7982 30548 8034
rect 30492 7980 30548 7982
rect 30268 7362 30324 7364
rect 30268 7310 30270 7362
rect 30270 7310 30322 7362
rect 30322 7310 30324 7362
rect 30268 7308 30324 7310
rect 30156 7250 30212 7252
rect 30156 7198 30158 7250
rect 30158 7198 30210 7250
rect 30210 7198 30212 7250
rect 30156 7196 30212 7198
rect 29596 6524 29652 6580
rect 28924 5068 28980 5124
rect 28812 4844 28868 4900
rect 29372 6300 29428 6356
rect 29372 6076 29428 6132
rect 29036 4284 29092 4340
rect 28700 3500 28756 3556
rect 29932 6524 29988 6580
rect 29708 6300 29764 6356
rect 29708 5122 29764 5124
rect 29708 5070 29710 5122
rect 29710 5070 29762 5122
rect 29762 5070 29764 5122
rect 29708 5068 29764 5070
rect 30268 5516 30324 5572
rect 30604 6300 30660 6356
rect 30604 6130 30660 6132
rect 30604 6078 30606 6130
rect 30606 6078 30658 6130
rect 30658 6078 30660 6130
rect 30604 6076 30660 6078
rect 31052 12124 31108 12180
rect 31276 11564 31332 11620
rect 31388 11340 31444 11396
rect 31052 11228 31108 11284
rect 32508 15036 32564 15092
rect 31724 13468 31780 13524
rect 32284 14476 32340 14532
rect 33404 17666 33460 17668
rect 33404 17614 33406 17666
rect 33406 17614 33458 17666
rect 33458 17614 33460 17666
rect 33404 17612 33460 17614
rect 33852 20524 33908 20580
rect 33852 20076 33908 20132
rect 34188 21644 34244 21700
rect 34076 21308 34132 21364
rect 34188 20972 34244 21028
rect 34636 26460 34692 26516
rect 34524 24556 34580 24612
rect 35532 30434 35588 30436
rect 35532 30382 35534 30434
rect 35534 30382 35586 30434
rect 35586 30382 35588 30434
rect 35532 30380 35588 30382
rect 35196 29372 35252 29428
rect 35420 29820 35476 29876
rect 35084 29148 35140 29204
rect 35420 29148 35476 29204
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35084 28476 35140 28532
rect 36316 32396 36372 32452
rect 36092 32338 36148 32340
rect 36092 32286 36094 32338
rect 36094 32286 36146 32338
rect 36146 32286 36148 32338
rect 36092 32284 36148 32286
rect 35868 31666 35924 31668
rect 35868 31614 35870 31666
rect 35870 31614 35922 31666
rect 35922 31614 35924 31666
rect 35868 31612 35924 31614
rect 36092 31388 36148 31444
rect 35868 30940 35924 30996
rect 36204 30716 36260 30772
rect 36092 30210 36148 30212
rect 36092 30158 36094 30210
rect 36094 30158 36146 30210
rect 36146 30158 36148 30210
rect 36092 30156 36148 30158
rect 35980 29820 36036 29876
rect 36428 31052 36484 31108
rect 36540 31500 36596 31556
rect 35756 29426 35812 29428
rect 35756 29374 35758 29426
rect 35758 29374 35810 29426
rect 35810 29374 35812 29426
rect 35756 29372 35812 29374
rect 35868 28754 35924 28756
rect 35868 28702 35870 28754
rect 35870 28702 35922 28754
rect 35922 28702 35924 28754
rect 35868 28700 35924 28702
rect 36092 29148 36148 29204
rect 35756 28588 35812 28644
rect 35980 28642 36036 28644
rect 35980 28590 35982 28642
rect 35982 28590 36034 28642
rect 36034 28590 36036 28642
rect 35980 28588 36036 28590
rect 36092 28530 36148 28532
rect 36092 28478 36094 28530
rect 36094 28478 36146 28530
rect 36146 28478 36148 28530
rect 36092 28476 36148 28478
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35644 27468 35700 27524
rect 35308 27244 35364 27300
rect 34972 26684 35028 26740
rect 34972 26124 35028 26180
rect 34860 26012 34916 26068
rect 34748 25564 34804 25620
rect 34636 23660 34692 23716
rect 34860 24780 34916 24836
rect 35196 26514 35252 26516
rect 35196 26462 35198 26514
rect 35198 26462 35250 26514
rect 35250 26462 35252 26514
rect 35196 26460 35252 26462
rect 35532 26796 35588 26852
rect 35420 26290 35476 26292
rect 35420 26238 35422 26290
rect 35422 26238 35474 26290
rect 35474 26238 35476 26290
rect 35420 26236 35476 26238
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35084 25116 35140 25172
rect 35308 25228 35364 25284
rect 34972 24668 35028 24724
rect 34748 23548 34804 23604
rect 34636 23154 34692 23156
rect 34636 23102 34638 23154
rect 34638 23102 34690 23154
rect 34690 23102 34692 23154
rect 34636 23100 34692 23102
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35196 23436 35252 23492
rect 35084 23266 35140 23268
rect 35084 23214 35086 23266
rect 35086 23214 35138 23266
rect 35138 23214 35140 23266
rect 35084 23212 35140 23214
rect 36316 28028 36372 28084
rect 36988 32562 37044 32564
rect 36988 32510 36990 32562
rect 36990 32510 37042 32562
rect 37042 32510 37044 32562
rect 36988 32508 37044 32510
rect 36876 31612 36932 31668
rect 36764 30994 36820 30996
rect 36764 30942 36766 30994
rect 36766 30942 36818 30994
rect 36818 30942 36820 30994
rect 36764 30940 36820 30942
rect 36652 30828 36708 30884
rect 36876 31052 36932 31108
rect 36652 27916 36708 27972
rect 36764 28028 36820 28084
rect 36540 27356 36596 27412
rect 36540 26796 36596 26852
rect 35868 25788 35924 25844
rect 35756 25282 35812 25284
rect 35756 25230 35758 25282
rect 35758 25230 35810 25282
rect 35810 25230 35812 25282
rect 35756 25228 35812 25230
rect 35532 23436 35588 23492
rect 35644 23212 35700 23268
rect 35532 23100 35588 23156
rect 34972 22988 35028 23044
rect 34636 22876 34692 22932
rect 35644 23042 35700 23044
rect 35644 22990 35646 23042
rect 35646 22990 35698 23042
rect 35698 22990 35700 23042
rect 35644 22988 35700 22990
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35644 22482 35700 22484
rect 35644 22430 35646 22482
rect 35646 22430 35698 22482
rect 35698 22430 35700 22482
rect 35644 22428 35700 22430
rect 35196 22146 35252 22148
rect 35196 22094 35198 22146
rect 35198 22094 35250 22146
rect 35250 22094 35252 22146
rect 35196 22092 35252 22094
rect 35644 21980 35700 22036
rect 34972 21868 35028 21924
rect 35308 21868 35364 21924
rect 35532 21756 35588 21812
rect 34188 20802 34244 20804
rect 34188 20750 34190 20802
rect 34190 20750 34242 20802
rect 34242 20750 34244 20802
rect 34188 20748 34244 20750
rect 34076 20412 34132 20468
rect 33964 19292 34020 19348
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 34748 21026 34804 21028
rect 34748 20974 34750 21026
rect 34750 20974 34802 21026
rect 34802 20974 34804 21026
rect 34748 20972 34804 20974
rect 34860 20860 34916 20916
rect 34636 20748 34692 20804
rect 34636 20300 34692 20356
rect 34412 19516 34468 19572
rect 34524 19740 34580 19796
rect 34188 18450 34244 18452
rect 34188 18398 34190 18450
rect 34190 18398 34242 18450
rect 34242 18398 34244 18450
rect 34188 18396 34244 18398
rect 33852 17612 33908 17668
rect 34188 17666 34244 17668
rect 34188 17614 34190 17666
rect 34190 17614 34242 17666
rect 34242 17614 34244 17666
rect 34188 17612 34244 17614
rect 33964 17164 34020 17220
rect 34076 17106 34132 17108
rect 34076 17054 34078 17106
rect 34078 17054 34130 17106
rect 34130 17054 34132 17106
rect 34076 17052 34132 17054
rect 34188 16994 34244 16996
rect 34188 16942 34190 16994
rect 34190 16942 34242 16994
rect 34242 16942 34244 16994
rect 34188 16940 34244 16942
rect 34188 16604 34244 16660
rect 34076 16098 34132 16100
rect 34076 16046 34078 16098
rect 34078 16046 34130 16098
rect 34130 16046 34132 16098
rect 34076 16044 34132 16046
rect 33628 15932 33684 15988
rect 34188 15986 34244 15988
rect 34188 15934 34190 15986
rect 34190 15934 34242 15986
rect 34242 15934 34244 15986
rect 34188 15932 34244 15934
rect 33516 15260 33572 15316
rect 32732 14530 32788 14532
rect 32732 14478 32734 14530
rect 32734 14478 32786 14530
rect 32786 14478 32788 14530
rect 32732 14476 32788 14478
rect 32508 13916 32564 13972
rect 32396 13746 32452 13748
rect 32396 13694 32398 13746
rect 32398 13694 32450 13746
rect 32450 13694 32452 13746
rect 32396 13692 32452 13694
rect 32396 13468 32452 13524
rect 31500 11228 31556 11284
rect 32172 11282 32228 11284
rect 32172 11230 32174 11282
rect 32174 11230 32226 11282
rect 32226 11230 32228 11282
rect 32172 11228 32228 11230
rect 32620 13468 32676 13524
rect 32844 13580 32900 13636
rect 32956 13468 33012 13524
rect 32956 12572 33012 12628
rect 32396 10780 32452 10836
rect 32172 10668 32228 10724
rect 32620 10722 32676 10724
rect 32620 10670 32622 10722
rect 32622 10670 32674 10722
rect 32674 10670 32676 10722
rect 32620 10668 32676 10670
rect 31388 9772 31444 9828
rect 31500 10556 31556 10612
rect 30940 8876 30996 8932
rect 32508 10610 32564 10612
rect 32508 10558 32510 10610
rect 32510 10558 32562 10610
rect 32562 10558 32564 10610
rect 32508 10556 32564 10558
rect 33964 15314 34020 15316
rect 33964 15262 33966 15314
rect 33966 15262 34018 15314
rect 34018 15262 34020 15314
rect 33964 15260 34020 15262
rect 34412 18562 34468 18564
rect 34412 18510 34414 18562
rect 34414 18510 34466 18562
rect 34466 18510 34468 18562
rect 34412 18508 34468 18510
rect 36092 25116 36148 25172
rect 36428 25788 36484 25844
rect 36316 24722 36372 24724
rect 36316 24670 36318 24722
rect 36318 24670 36370 24722
rect 36370 24670 36372 24722
rect 36316 24668 36372 24670
rect 35868 23548 35924 23604
rect 36092 23996 36148 24052
rect 36204 23884 36260 23940
rect 36316 21868 36372 21924
rect 36204 21756 36260 21812
rect 35532 20188 35588 20244
rect 35084 20076 35140 20132
rect 34972 19794 35028 19796
rect 34972 19742 34974 19794
rect 34974 19742 35026 19794
rect 35026 19742 35028 19794
rect 34972 19740 35028 19742
rect 34748 19346 34804 19348
rect 34748 19294 34750 19346
rect 34750 19294 34802 19346
rect 34802 19294 34804 19346
rect 34748 19292 34804 19294
rect 34860 19180 34916 19236
rect 34636 18620 34692 18676
rect 34748 18844 34804 18900
rect 34636 17612 34692 17668
rect 34748 18284 34804 18340
rect 34524 17052 34580 17108
rect 33516 12572 33572 12628
rect 33628 14028 33684 14084
rect 33740 13746 33796 13748
rect 33740 13694 33742 13746
rect 33742 13694 33794 13746
rect 33794 13694 33796 13746
rect 33740 13692 33796 13694
rect 33852 13580 33908 13636
rect 33964 13804 34020 13860
rect 32956 10780 33012 10836
rect 32172 9826 32228 9828
rect 32172 9774 32174 9826
rect 32174 9774 32226 9826
rect 32226 9774 32228 9826
rect 32172 9772 32228 9774
rect 31612 9154 31668 9156
rect 31612 9102 31614 9154
rect 31614 9102 31666 9154
rect 31666 9102 31668 9154
rect 31612 9100 31668 9102
rect 31164 8316 31220 8372
rect 32844 9548 32900 9604
rect 32396 8652 32452 8708
rect 31612 7474 31668 7476
rect 31612 7422 31614 7474
rect 31614 7422 31666 7474
rect 31666 7422 31668 7474
rect 31612 7420 31668 7422
rect 31276 7362 31332 7364
rect 31276 7310 31278 7362
rect 31278 7310 31330 7362
rect 31330 7310 31332 7362
rect 31276 7308 31332 7310
rect 31164 7196 31220 7252
rect 30380 4732 30436 4788
rect 31836 7308 31892 7364
rect 30828 5740 30884 5796
rect 30380 4562 30436 4564
rect 30380 4510 30382 4562
rect 30382 4510 30434 4562
rect 30434 4510 30436 4562
rect 30380 4508 30436 4510
rect 32620 7474 32676 7476
rect 32620 7422 32622 7474
rect 32622 7422 32674 7474
rect 32674 7422 32676 7474
rect 32620 7420 32676 7422
rect 32844 8034 32900 8036
rect 32844 7982 32846 8034
rect 32846 7982 32898 8034
rect 32898 7982 32900 8034
rect 32844 7980 32900 7982
rect 33628 11116 33684 11172
rect 34300 14028 34356 14084
rect 34076 13634 34132 13636
rect 34076 13582 34078 13634
rect 34078 13582 34130 13634
rect 34130 13582 34132 13634
rect 34076 13580 34132 13582
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35868 21586 35924 21588
rect 35868 21534 35870 21586
rect 35870 21534 35922 21586
rect 35922 21534 35924 21586
rect 35868 21532 35924 21534
rect 35756 20972 35812 21028
rect 36092 20914 36148 20916
rect 36092 20862 36094 20914
rect 36094 20862 36146 20914
rect 36146 20862 36148 20914
rect 36092 20860 36148 20862
rect 35868 20524 35924 20580
rect 35980 20076 36036 20132
rect 36652 26684 36708 26740
rect 36652 26124 36708 26180
rect 36988 30044 37044 30100
rect 36988 27804 37044 27860
rect 37100 27580 37156 27636
rect 36876 27468 36932 27524
rect 36876 27132 36932 27188
rect 38892 57820 38948 57876
rect 38108 57148 38164 57204
rect 38220 57036 38276 57092
rect 37772 56924 37828 56980
rect 38668 57260 38724 57316
rect 38444 57036 38500 57092
rect 40796 59500 40852 59556
rect 40572 59276 40628 59332
rect 40348 58994 40404 58996
rect 40348 58942 40350 58994
rect 40350 58942 40402 58994
rect 40402 58942 40404 58994
rect 40348 58940 40404 58942
rect 40572 58828 40628 58884
rect 42028 59330 42084 59332
rect 42028 59278 42030 59330
rect 42030 59278 42082 59330
rect 42082 59278 42084 59330
rect 42028 59276 42084 59278
rect 41468 59218 41524 59220
rect 41468 59166 41470 59218
rect 41470 59166 41522 59218
rect 41522 59166 41524 59218
rect 41468 59164 41524 59166
rect 41804 58940 41860 58996
rect 41580 58716 41636 58772
rect 40796 58492 40852 58548
rect 41244 58604 41300 58660
rect 40348 58380 40404 58436
rect 40236 58322 40292 58324
rect 40236 58270 40238 58322
rect 40238 58270 40290 58322
rect 40290 58270 40292 58322
rect 40236 58268 40292 58270
rect 38780 57596 38836 57652
rect 38556 56924 38612 56980
rect 38332 56812 38388 56868
rect 38780 56866 38836 56868
rect 38780 56814 38782 56866
rect 38782 56814 38834 56866
rect 38834 56814 38836 56866
rect 38780 56812 38836 56814
rect 38556 56754 38612 56756
rect 38556 56702 38558 56754
rect 38558 56702 38610 56754
rect 38610 56702 38612 56754
rect 38556 56700 38612 56702
rect 37548 53564 37604 53620
rect 37548 51602 37604 51604
rect 37548 51550 37550 51602
rect 37550 51550 37602 51602
rect 37602 51550 37604 51602
rect 37548 51548 37604 51550
rect 37324 51378 37380 51380
rect 37324 51326 37326 51378
rect 37326 51326 37378 51378
rect 37378 51326 37380 51378
rect 37324 51324 37380 51326
rect 37660 50988 37716 51044
rect 37660 50706 37716 50708
rect 37660 50654 37662 50706
rect 37662 50654 37714 50706
rect 37714 50654 37716 50706
rect 37660 50652 37716 50654
rect 37548 49084 37604 49140
rect 37436 47458 37492 47460
rect 37436 47406 37438 47458
rect 37438 47406 37490 47458
rect 37490 47406 37492 47458
rect 37436 47404 37492 47406
rect 37548 47292 37604 47348
rect 38220 56364 38276 56420
rect 38668 55916 38724 55972
rect 38556 55468 38612 55524
rect 39116 56700 39172 56756
rect 39004 56476 39060 56532
rect 39452 57650 39508 57652
rect 39452 57598 39454 57650
rect 39454 57598 39506 57650
rect 39506 57598 39508 57650
rect 39452 57596 39508 57598
rect 39340 56866 39396 56868
rect 39340 56814 39342 56866
rect 39342 56814 39394 56866
rect 39394 56814 39396 56866
rect 39340 56812 39396 56814
rect 42364 59164 42420 59220
rect 42476 58828 42532 58884
rect 42812 58546 42868 58548
rect 42812 58494 42814 58546
rect 42814 58494 42866 58546
rect 42866 58494 42868 58546
rect 42812 58492 42868 58494
rect 43148 58492 43204 58548
rect 43036 58156 43092 58212
rect 43708 58716 43764 58772
rect 43596 58492 43652 58548
rect 43484 58156 43540 58212
rect 43260 57874 43316 57876
rect 43260 57822 43262 57874
rect 43262 57822 43314 57874
rect 43314 57822 43316 57874
rect 43260 57820 43316 57822
rect 43484 57874 43540 57876
rect 43484 57822 43486 57874
rect 43486 57822 43538 57874
rect 43538 57822 43540 57874
rect 43484 57820 43540 57822
rect 40684 57484 40740 57540
rect 40348 56812 40404 56868
rect 39788 56364 39844 56420
rect 40236 56642 40292 56644
rect 40236 56590 40238 56642
rect 40238 56590 40290 56642
rect 40290 56590 40292 56642
rect 40236 56588 40292 56590
rect 39228 55916 39284 55972
rect 41020 56642 41076 56644
rect 41020 56590 41022 56642
rect 41022 56590 41074 56642
rect 41074 56590 41076 56642
rect 41020 56588 41076 56590
rect 39564 55858 39620 55860
rect 39564 55806 39566 55858
rect 39566 55806 39618 55858
rect 39618 55806 39620 55858
rect 39564 55804 39620 55806
rect 40348 55692 40404 55748
rect 42588 57260 42644 57316
rect 43372 57538 43428 57540
rect 43372 57486 43374 57538
rect 43374 57486 43426 57538
rect 43426 57486 43428 57538
rect 43372 57484 43428 57486
rect 44492 58604 44548 58660
rect 44940 59218 44996 59220
rect 44940 59166 44942 59218
rect 44942 59166 44994 59218
rect 44994 59166 44996 59218
rect 44940 59164 44996 59166
rect 49868 59778 49924 59780
rect 49868 59726 49870 59778
rect 49870 59726 49922 59778
rect 49922 59726 49924 59778
rect 49868 59724 49924 59726
rect 50428 59724 50484 59780
rect 50556 59610 50612 59612
rect 50556 59558 50558 59610
rect 50558 59558 50610 59610
rect 50610 59558 50612 59610
rect 50556 59556 50612 59558
rect 50660 59610 50716 59612
rect 50660 59558 50662 59610
rect 50662 59558 50714 59610
rect 50714 59558 50716 59610
rect 50660 59556 50716 59558
rect 50764 59610 50820 59612
rect 50764 59558 50766 59610
rect 50766 59558 50818 59610
rect 50818 59558 50820 59610
rect 50764 59556 50820 59558
rect 45500 59330 45556 59332
rect 45500 59278 45502 59330
rect 45502 59278 45554 59330
rect 45554 59278 45556 59330
rect 45500 59276 45556 59278
rect 45388 59218 45444 59220
rect 45388 59166 45390 59218
rect 45390 59166 45442 59218
rect 45442 59166 45444 59218
rect 45388 59164 45444 59166
rect 45052 58492 45108 58548
rect 44380 57932 44436 57988
rect 44492 58268 44548 58324
rect 44268 57820 44324 57876
rect 44604 57932 44660 57988
rect 45388 57820 45444 57876
rect 43820 57090 43876 57092
rect 43820 57038 43822 57090
rect 43822 57038 43874 57090
rect 43874 57038 43876 57090
rect 43820 57036 43876 57038
rect 44156 57036 44212 57092
rect 42812 56306 42868 56308
rect 42812 56254 42814 56306
rect 42814 56254 42866 56306
rect 42866 56254 42868 56306
rect 42812 56252 42868 56254
rect 43932 56306 43988 56308
rect 43932 56254 43934 56306
rect 43934 56254 43986 56306
rect 43986 56254 43988 56306
rect 43932 56252 43988 56254
rect 45500 57036 45556 57092
rect 46396 58546 46452 58548
rect 46396 58494 46398 58546
rect 46398 58494 46450 58546
rect 46450 58494 46452 58546
rect 46396 58492 46452 58494
rect 46732 58492 46788 58548
rect 46620 58434 46676 58436
rect 46620 58382 46622 58434
rect 46622 58382 46674 58434
rect 46674 58382 46676 58434
rect 46620 58380 46676 58382
rect 46060 57932 46116 57988
rect 47180 58546 47236 58548
rect 47180 58494 47182 58546
rect 47182 58494 47234 58546
rect 47234 58494 47236 58546
rect 47180 58492 47236 58494
rect 47516 58434 47572 58436
rect 47516 58382 47518 58434
rect 47518 58382 47570 58434
rect 47570 58382 47572 58434
rect 47516 58380 47572 58382
rect 50092 58434 50148 58436
rect 50092 58382 50094 58434
rect 50094 58382 50146 58434
rect 50146 58382 50148 58434
rect 50092 58380 50148 58382
rect 47292 58210 47348 58212
rect 47292 58158 47294 58210
rect 47294 58158 47346 58210
rect 47346 58158 47348 58210
rect 47292 58156 47348 58158
rect 50556 58042 50612 58044
rect 50556 57990 50558 58042
rect 50558 57990 50610 58042
rect 50610 57990 50612 58042
rect 50556 57988 50612 57990
rect 50660 58042 50716 58044
rect 50660 57990 50662 58042
rect 50662 57990 50714 58042
rect 50714 57990 50716 58042
rect 50660 57988 50716 57990
rect 50764 58042 50820 58044
rect 50764 57990 50766 58042
rect 50766 57990 50818 58042
rect 50818 57990 50820 58042
rect 50764 57988 50820 57990
rect 45948 57036 46004 57092
rect 44604 56082 44660 56084
rect 44604 56030 44606 56082
rect 44606 56030 44658 56082
rect 44658 56030 44660 56082
rect 44604 56028 44660 56030
rect 43372 55970 43428 55972
rect 43372 55918 43374 55970
rect 43374 55918 43426 55970
rect 43426 55918 43428 55970
rect 43372 55916 43428 55918
rect 43260 55522 43316 55524
rect 43260 55470 43262 55522
rect 43262 55470 43314 55522
rect 43314 55470 43316 55522
rect 43260 55468 43316 55470
rect 38108 55298 38164 55300
rect 38108 55246 38110 55298
rect 38110 55246 38162 55298
rect 38162 55246 38164 55298
rect 38108 55244 38164 55246
rect 39452 55298 39508 55300
rect 39452 55246 39454 55298
rect 39454 55246 39506 55298
rect 39506 55246 39508 55298
rect 39452 55244 39508 55246
rect 37884 55132 37940 55188
rect 38668 55186 38724 55188
rect 38668 55134 38670 55186
rect 38670 55134 38722 55186
rect 38722 55134 38724 55186
rect 38668 55132 38724 55134
rect 38780 54684 38836 54740
rect 39676 55298 39732 55300
rect 39676 55246 39678 55298
rect 39678 55246 39730 55298
rect 39730 55246 39732 55298
rect 39676 55244 39732 55246
rect 40460 55298 40516 55300
rect 40460 55246 40462 55298
rect 40462 55246 40514 55298
rect 40514 55246 40516 55298
rect 40460 55244 40516 55246
rect 40684 55132 40740 55188
rect 41580 55244 41636 55300
rect 39788 54684 39844 54740
rect 40460 55020 40516 55076
rect 38332 53676 38388 53732
rect 39564 53730 39620 53732
rect 39564 53678 39566 53730
rect 39566 53678 39618 53730
rect 39618 53678 39620 53730
rect 39564 53676 39620 53678
rect 40348 53954 40404 53956
rect 40348 53902 40350 53954
rect 40350 53902 40402 53954
rect 40402 53902 40404 53954
rect 40348 53900 40404 53902
rect 39340 52220 39396 52276
rect 39228 52108 39284 52164
rect 38556 50706 38612 50708
rect 38556 50654 38558 50706
rect 38558 50654 38610 50706
rect 38610 50654 38612 50706
rect 38556 50652 38612 50654
rect 37884 50594 37940 50596
rect 37884 50542 37886 50594
rect 37886 50542 37938 50594
rect 37938 50542 37940 50594
rect 37884 50540 37940 50542
rect 38556 50428 38612 50484
rect 38332 49138 38388 49140
rect 38332 49086 38334 49138
rect 38334 49086 38386 49138
rect 38386 49086 38388 49138
rect 38332 49084 38388 49086
rect 37884 48636 37940 48692
rect 37884 48242 37940 48244
rect 37884 48190 37886 48242
rect 37886 48190 37938 48242
rect 37938 48190 37940 48242
rect 37884 48188 37940 48190
rect 37772 47180 37828 47236
rect 37996 47068 38052 47124
rect 38444 48188 38500 48244
rect 39116 50428 39172 50484
rect 39564 52780 39620 52836
rect 40348 52834 40404 52836
rect 40348 52782 40350 52834
rect 40350 52782 40402 52834
rect 40402 52782 40404 52834
rect 40348 52780 40404 52782
rect 39564 52108 39620 52164
rect 39900 52274 39956 52276
rect 39900 52222 39902 52274
rect 39902 52222 39954 52274
rect 39954 52222 39956 52274
rect 39900 52220 39956 52222
rect 39788 52162 39844 52164
rect 39788 52110 39790 52162
rect 39790 52110 39842 52162
rect 39842 52110 39844 52162
rect 39788 52108 39844 52110
rect 39788 50988 39844 51044
rect 39340 50652 39396 50708
rect 38780 48130 38836 48132
rect 38780 48078 38782 48130
rect 38782 48078 38834 48130
rect 38834 48078 38836 48130
rect 38780 48076 38836 48078
rect 38108 47180 38164 47236
rect 38668 47234 38724 47236
rect 38668 47182 38670 47234
rect 38670 47182 38722 47234
rect 38722 47182 38724 47234
rect 38668 47180 38724 47182
rect 38444 46898 38500 46900
rect 38444 46846 38446 46898
rect 38446 46846 38498 46898
rect 38498 46846 38500 46898
rect 38444 46844 38500 46846
rect 37772 46060 37828 46116
rect 38556 46114 38612 46116
rect 38556 46062 38558 46114
rect 38558 46062 38610 46114
rect 38610 46062 38612 46114
rect 38556 46060 38612 46062
rect 37996 46002 38052 46004
rect 37996 45950 37998 46002
rect 37998 45950 38050 46002
rect 38050 45950 38052 46002
rect 37996 45948 38052 45950
rect 37772 45890 37828 45892
rect 37772 45838 37774 45890
rect 37774 45838 37826 45890
rect 37826 45838 37828 45890
rect 37772 45836 37828 45838
rect 38668 45724 38724 45780
rect 38444 45612 38500 45668
rect 38220 45218 38276 45220
rect 38220 45166 38222 45218
rect 38222 45166 38274 45218
rect 38274 45166 38276 45218
rect 38220 45164 38276 45166
rect 37548 44994 37604 44996
rect 37548 44942 37550 44994
rect 37550 44942 37602 44994
rect 37602 44942 37604 44994
rect 37548 44940 37604 44942
rect 37548 43708 37604 43764
rect 37884 43596 37940 43652
rect 38108 44156 38164 44212
rect 37324 43538 37380 43540
rect 37324 43486 37326 43538
rect 37326 43486 37378 43538
rect 37378 43486 37380 43538
rect 37324 43484 37380 43486
rect 38220 43762 38276 43764
rect 38220 43710 38222 43762
rect 38222 43710 38274 43762
rect 38274 43710 38276 43762
rect 38220 43708 38276 43710
rect 37548 42364 37604 42420
rect 37436 42194 37492 42196
rect 37436 42142 37438 42194
rect 37438 42142 37490 42194
rect 37490 42142 37492 42194
rect 37436 42140 37492 42142
rect 37660 42252 37716 42308
rect 37324 41916 37380 41972
rect 37996 42588 38052 42644
rect 37884 42028 37940 42084
rect 37660 40348 37716 40404
rect 37772 41132 37828 41188
rect 38780 45330 38836 45332
rect 38780 45278 38782 45330
rect 38782 45278 38834 45330
rect 38834 45278 38836 45330
rect 38780 45276 38836 45278
rect 38780 44380 38836 44436
rect 39900 50764 39956 50820
rect 40348 50764 40404 50820
rect 40348 50482 40404 50484
rect 40348 50430 40350 50482
rect 40350 50430 40402 50482
rect 40402 50430 40404 50482
rect 40348 50428 40404 50430
rect 42476 55298 42532 55300
rect 42476 55246 42478 55298
rect 42478 55246 42530 55298
rect 42530 55246 42532 55298
rect 42476 55244 42532 55246
rect 41804 54738 41860 54740
rect 41804 54686 41806 54738
rect 41806 54686 41858 54738
rect 41858 54686 41860 54738
rect 41804 54684 41860 54686
rect 41916 54626 41972 54628
rect 41916 54574 41918 54626
rect 41918 54574 41970 54626
rect 41970 54574 41972 54626
rect 41916 54572 41972 54574
rect 44380 55970 44436 55972
rect 44380 55918 44382 55970
rect 44382 55918 44434 55970
rect 44434 55918 44436 55970
rect 44380 55916 44436 55918
rect 44828 55970 44884 55972
rect 44828 55918 44830 55970
rect 44830 55918 44882 55970
rect 44882 55918 44884 55970
rect 44828 55916 44884 55918
rect 44044 55804 44100 55860
rect 46284 55468 46340 55524
rect 46956 57650 47012 57652
rect 46956 57598 46958 57650
rect 46958 57598 47010 57650
rect 47010 57598 47012 57650
rect 46956 57596 47012 57598
rect 47068 57372 47124 57428
rect 47740 57650 47796 57652
rect 47740 57598 47742 57650
rect 47742 57598 47794 57650
rect 47794 57598 47796 57650
rect 47740 57596 47796 57598
rect 47516 57372 47572 57428
rect 43372 55020 43428 55076
rect 46508 56588 46564 56644
rect 47740 56642 47796 56644
rect 47740 56590 47742 56642
rect 47742 56590 47794 56642
rect 47794 56590 47796 56642
rect 47740 56588 47796 56590
rect 46508 56028 46564 56084
rect 46732 56082 46788 56084
rect 46732 56030 46734 56082
rect 46734 56030 46786 56082
rect 46786 56030 46788 56082
rect 46732 56028 46788 56030
rect 48412 57596 48468 57652
rect 48188 56866 48244 56868
rect 48188 56814 48190 56866
rect 48190 56814 48242 56866
rect 48242 56814 48244 56866
rect 48188 56812 48244 56814
rect 48300 57372 48356 57428
rect 49980 57484 50036 57540
rect 50092 56866 50148 56868
rect 50092 56814 50094 56866
rect 50094 56814 50146 56866
rect 50146 56814 50148 56866
rect 50092 56812 50148 56814
rect 47852 56028 47908 56084
rect 46508 55804 46564 55860
rect 47852 55692 47908 55748
rect 47740 55298 47796 55300
rect 47740 55246 47742 55298
rect 47742 55246 47794 55298
rect 47794 55246 47796 55298
rect 47740 55244 47796 55246
rect 47964 54684 48020 54740
rect 48076 55132 48132 55188
rect 42588 54572 42644 54628
rect 41580 53900 41636 53956
rect 41692 54236 41748 54292
rect 40572 53788 40628 53844
rect 41692 53788 41748 53844
rect 42140 53228 42196 53284
rect 41132 52162 41188 52164
rect 41132 52110 41134 52162
rect 41134 52110 41186 52162
rect 41186 52110 41188 52162
rect 41132 52108 41188 52110
rect 42700 53228 42756 53284
rect 43148 54290 43204 54292
rect 43148 54238 43150 54290
rect 43150 54238 43202 54290
rect 43202 54238 43204 54290
rect 43148 54236 43204 54238
rect 44044 54236 44100 54292
rect 42924 53228 42980 53284
rect 44716 53842 44772 53844
rect 44716 53790 44718 53842
rect 44718 53790 44770 53842
rect 44770 53790 44772 53842
rect 44716 53788 44772 53790
rect 45948 53842 46004 53844
rect 45948 53790 45950 53842
rect 45950 53790 46002 53842
rect 46002 53790 46004 53842
rect 45948 53788 46004 53790
rect 46844 53730 46900 53732
rect 46844 53678 46846 53730
rect 46846 53678 46898 53730
rect 46898 53678 46900 53730
rect 46844 53676 46900 53678
rect 45276 53340 45332 53396
rect 41916 50818 41972 50820
rect 41916 50766 41918 50818
rect 41918 50766 41970 50818
rect 41970 50766 41972 50818
rect 41916 50764 41972 50766
rect 39676 49922 39732 49924
rect 39676 49870 39678 49922
rect 39678 49870 39730 49922
rect 39730 49870 39732 49922
rect 39676 49868 39732 49870
rect 40348 49922 40404 49924
rect 40348 49870 40350 49922
rect 40350 49870 40402 49922
rect 40402 49870 40404 49922
rect 40348 49868 40404 49870
rect 39452 47346 39508 47348
rect 39452 47294 39454 47346
rect 39454 47294 39506 47346
rect 39506 47294 39508 47346
rect 39452 47292 39508 47294
rect 40460 48860 40516 48916
rect 40908 50372 40964 50428
rect 41580 50594 41636 50596
rect 41580 50542 41582 50594
rect 41582 50542 41634 50594
rect 41634 50542 41636 50594
rect 41580 50540 41636 50542
rect 40684 48300 40740 48356
rect 40796 48748 40852 48804
rect 39676 48130 39732 48132
rect 39676 48078 39678 48130
rect 39678 48078 39730 48130
rect 39730 48078 39732 48130
rect 39676 48076 39732 48078
rect 40012 47404 40068 47460
rect 39676 47292 39732 47348
rect 39228 46060 39284 46116
rect 39452 45948 39508 46004
rect 38444 42476 38500 42532
rect 38668 41970 38724 41972
rect 38668 41918 38670 41970
rect 38670 41918 38722 41970
rect 38722 41918 38724 41970
rect 38668 41916 38724 41918
rect 37996 41580 38052 41636
rect 37324 40236 37380 40292
rect 37548 39116 37604 39172
rect 37324 38892 37380 38948
rect 37436 37266 37492 37268
rect 37436 37214 37438 37266
rect 37438 37214 37490 37266
rect 37490 37214 37492 37266
rect 37436 37212 37492 37214
rect 37436 36258 37492 36260
rect 37436 36206 37438 36258
rect 37438 36206 37490 36258
rect 37490 36206 37492 36258
rect 37436 36204 37492 36206
rect 37324 35698 37380 35700
rect 37324 35646 37326 35698
rect 37326 35646 37378 35698
rect 37378 35646 37380 35698
rect 37324 35644 37380 35646
rect 37548 35084 37604 35140
rect 37324 34300 37380 34356
rect 37548 34188 37604 34244
rect 37548 33628 37604 33684
rect 37436 33346 37492 33348
rect 37436 33294 37438 33346
rect 37438 33294 37490 33346
rect 37490 33294 37492 33346
rect 37436 33292 37492 33294
rect 37436 32284 37492 32340
rect 38556 41074 38612 41076
rect 38556 41022 38558 41074
rect 38558 41022 38610 41074
rect 38610 41022 38612 41074
rect 38556 41020 38612 41022
rect 37996 40348 38052 40404
rect 38444 40514 38500 40516
rect 38444 40462 38446 40514
rect 38446 40462 38498 40514
rect 38498 40462 38500 40514
rect 38444 40460 38500 40462
rect 38556 40348 38612 40404
rect 37772 38556 37828 38612
rect 37884 36482 37940 36484
rect 37884 36430 37886 36482
rect 37886 36430 37938 36482
rect 37938 36430 37940 36482
rect 37884 36428 37940 36430
rect 37772 35308 37828 35364
rect 37324 31612 37380 31668
rect 37436 31554 37492 31556
rect 37436 31502 37438 31554
rect 37438 31502 37490 31554
rect 37490 31502 37492 31554
rect 37436 31500 37492 31502
rect 38332 38050 38388 38052
rect 38332 37998 38334 38050
rect 38334 37998 38386 38050
rect 38386 37998 38388 38050
rect 38332 37996 38388 37998
rect 38108 37772 38164 37828
rect 38444 37548 38500 37604
rect 38332 37436 38388 37492
rect 38332 35980 38388 36036
rect 38892 41916 38948 41972
rect 38892 41132 38948 41188
rect 38892 40402 38948 40404
rect 38892 40350 38894 40402
rect 38894 40350 38946 40402
rect 38946 40350 38948 40402
rect 38892 40348 38948 40350
rect 38780 38668 38836 38724
rect 39116 41804 39172 41860
rect 40348 47346 40404 47348
rect 40348 47294 40350 47346
rect 40350 47294 40402 47346
rect 40402 47294 40404 47346
rect 40348 47292 40404 47294
rect 40572 47346 40628 47348
rect 40572 47294 40574 47346
rect 40574 47294 40626 47346
rect 40626 47294 40628 47346
rect 40572 47292 40628 47294
rect 40460 47068 40516 47124
rect 40236 45778 40292 45780
rect 40236 45726 40238 45778
rect 40238 45726 40290 45778
rect 40290 45726 40292 45778
rect 40236 45724 40292 45726
rect 39564 45666 39620 45668
rect 39564 45614 39566 45666
rect 39566 45614 39618 45666
rect 39618 45614 39620 45666
rect 39564 45612 39620 45614
rect 39676 44380 39732 44436
rect 39900 44434 39956 44436
rect 39900 44382 39902 44434
rect 39902 44382 39954 44434
rect 39954 44382 39956 44434
rect 39900 44380 39956 44382
rect 40348 44994 40404 44996
rect 40348 44942 40350 44994
rect 40350 44942 40402 44994
rect 40402 44942 40404 44994
rect 40348 44940 40404 44942
rect 40236 44434 40292 44436
rect 40236 44382 40238 44434
rect 40238 44382 40290 44434
rect 40290 44382 40292 44434
rect 40236 44380 40292 44382
rect 40012 44268 40068 44324
rect 39676 44210 39732 44212
rect 39676 44158 39678 44210
rect 39678 44158 39730 44210
rect 39730 44158 39732 44210
rect 39676 44156 39732 44158
rect 39564 44044 39620 44100
rect 39676 43650 39732 43652
rect 39676 43598 39678 43650
rect 39678 43598 39730 43650
rect 39730 43598 39732 43650
rect 39676 43596 39732 43598
rect 40348 43650 40404 43652
rect 40348 43598 40350 43650
rect 40350 43598 40402 43650
rect 40402 43598 40404 43650
rect 40348 43596 40404 43598
rect 40572 45666 40628 45668
rect 40572 45614 40574 45666
rect 40574 45614 40626 45666
rect 40626 45614 40628 45666
rect 40572 45612 40628 45614
rect 40572 44604 40628 44660
rect 40572 43538 40628 43540
rect 40572 43486 40574 43538
rect 40574 43486 40626 43538
rect 40626 43486 40628 43538
rect 40572 43484 40628 43486
rect 40460 43372 40516 43428
rect 39788 42642 39844 42644
rect 39788 42590 39790 42642
rect 39790 42590 39842 42642
rect 39842 42590 39844 42642
rect 39788 42588 39844 42590
rect 39676 41804 39732 41860
rect 39452 41186 39508 41188
rect 39452 41134 39454 41186
rect 39454 41134 39506 41186
rect 39506 41134 39508 41186
rect 39452 41132 39508 41134
rect 39788 41468 39844 41524
rect 39004 40236 39060 40292
rect 39228 40796 39284 40852
rect 38668 37548 38724 37604
rect 38780 37490 38836 37492
rect 38780 37438 38782 37490
rect 38782 37438 38834 37490
rect 38834 37438 38836 37490
rect 38780 37436 38836 37438
rect 38780 36988 38836 37044
rect 38668 36876 38724 36932
rect 38108 35084 38164 35140
rect 37884 34914 37940 34916
rect 37884 34862 37886 34914
rect 37886 34862 37938 34914
rect 37938 34862 37940 34914
rect 37884 34860 37940 34862
rect 38220 34188 38276 34244
rect 38556 34524 38612 34580
rect 38332 34076 38388 34132
rect 38108 33628 38164 33684
rect 38556 33404 38612 33460
rect 39004 38050 39060 38052
rect 39004 37998 39006 38050
rect 39006 37998 39058 38050
rect 39058 37998 39060 38050
rect 39004 37996 39060 37998
rect 39004 37548 39060 37604
rect 38892 34972 38948 35028
rect 39004 35532 39060 35588
rect 40348 42642 40404 42644
rect 40348 42590 40350 42642
rect 40350 42590 40402 42642
rect 40402 42590 40404 42642
rect 40348 42588 40404 42590
rect 40796 43426 40852 43428
rect 40796 43374 40798 43426
rect 40798 43374 40850 43426
rect 40850 43374 40852 43426
rect 40796 43372 40852 43374
rect 40796 42530 40852 42532
rect 40796 42478 40798 42530
rect 40798 42478 40850 42530
rect 40850 42478 40852 42530
rect 40796 42476 40852 42478
rect 41020 47458 41076 47460
rect 41020 47406 41022 47458
rect 41022 47406 41074 47458
rect 41074 47406 41076 47458
rect 41020 47404 41076 47406
rect 41804 48914 41860 48916
rect 41804 48862 41806 48914
rect 41806 48862 41858 48914
rect 41858 48862 41860 48914
rect 41804 48860 41860 48862
rect 42924 51324 42980 51380
rect 42588 50764 42644 50820
rect 42924 50540 42980 50596
rect 47516 54290 47572 54292
rect 47516 54238 47518 54290
rect 47518 54238 47570 54290
rect 47570 54238 47572 54290
rect 47516 54236 47572 54238
rect 50204 56252 50260 56308
rect 50204 56082 50260 56084
rect 50204 56030 50206 56082
rect 50206 56030 50258 56082
rect 50258 56030 50260 56082
rect 50204 56028 50260 56030
rect 48300 55244 48356 55300
rect 48524 55916 48580 55972
rect 48412 55186 48468 55188
rect 48412 55134 48414 55186
rect 48414 55134 48466 55186
rect 48466 55134 48468 55186
rect 48412 55132 48468 55134
rect 49532 55970 49588 55972
rect 49532 55918 49534 55970
rect 49534 55918 49586 55970
rect 49586 55918 49588 55970
rect 49532 55916 49588 55918
rect 48412 54738 48468 54740
rect 48412 54686 48414 54738
rect 48414 54686 48466 54738
rect 48466 54686 48468 54738
rect 48412 54684 48468 54686
rect 48524 54626 48580 54628
rect 48524 54574 48526 54626
rect 48526 54574 48578 54626
rect 48578 54574 48580 54626
rect 48524 54572 48580 54574
rect 50540 57538 50596 57540
rect 50540 57486 50542 57538
rect 50542 57486 50594 57538
rect 50594 57486 50596 57538
rect 50540 57484 50596 57486
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 53788 57820 53844 57876
rect 51884 57650 51940 57652
rect 51884 57598 51886 57650
rect 51886 57598 51938 57650
rect 51938 57598 51940 57650
rect 51884 57596 51940 57598
rect 51996 57538 52052 57540
rect 51996 57486 51998 57538
rect 51998 57486 52050 57538
rect 52050 57486 52052 57538
rect 51996 57484 52052 57486
rect 51548 57372 51604 57428
rect 51660 56924 51716 56980
rect 51324 56028 51380 56084
rect 51436 56252 51492 56308
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 51996 57036 52052 57092
rect 52108 56812 52164 56868
rect 52220 57596 52276 57652
rect 52332 56924 52388 56980
rect 52332 56754 52388 56756
rect 52332 56702 52334 56754
rect 52334 56702 52386 56754
rect 52386 56702 52388 56754
rect 52332 56700 52388 56702
rect 52220 56588 52276 56644
rect 52892 56588 52948 56644
rect 52220 56082 52276 56084
rect 52220 56030 52222 56082
rect 52222 56030 52274 56082
rect 52274 56030 52276 56082
rect 52220 56028 52276 56030
rect 53564 56588 53620 56644
rect 53900 56700 53956 56756
rect 53900 55970 53956 55972
rect 53900 55918 53902 55970
rect 53902 55918 53954 55970
rect 53954 55918 53956 55970
rect 53900 55916 53956 55918
rect 52892 55804 52948 55860
rect 54460 55970 54516 55972
rect 54460 55918 54462 55970
rect 54462 55918 54514 55970
rect 54514 55918 54516 55970
rect 54460 55916 54516 55918
rect 55132 55916 55188 55972
rect 51996 55244 52052 55300
rect 48300 54236 48356 54292
rect 48636 54348 48692 54404
rect 48524 53730 48580 53732
rect 48524 53678 48526 53730
rect 48526 53678 48578 53730
rect 48578 53678 48580 53730
rect 48524 53676 48580 53678
rect 48188 53618 48244 53620
rect 48188 53566 48190 53618
rect 48190 53566 48242 53618
rect 48242 53566 48244 53618
rect 48188 53564 48244 53566
rect 47292 53004 47348 53060
rect 47964 53506 48020 53508
rect 47964 53454 47966 53506
rect 47966 53454 48018 53506
rect 48018 53454 48020 53506
rect 47964 53452 48020 53454
rect 47740 52834 47796 52836
rect 47740 52782 47742 52834
rect 47742 52782 47794 52834
rect 47794 52782 47796 52834
rect 47740 52780 47796 52782
rect 45724 52108 45780 52164
rect 46172 52162 46228 52164
rect 46172 52110 46174 52162
rect 46174 52110 46226 52162
rect 46226 52110 46228 52162
rect 46172 52108 46228 52110
rect 45276 51436 45332 51492
rect 43148 51378 43204 51380
rect 43148 51326 43150 51378
rect 43150 51326 43202 51378
rect 43202 51326 43204 51378
rect 43148 51324 43204 51326
rect 44044 51378 44100 51380
rect 44044 51326 44046 51378
rect 44046 51326 44098 51378
rect 44098 51326 44100 51378
rect 44044 51324 44100 51326
rect 44940 51378 44996 51380
rect 44940 51326 44942 51378
rect 44942 51326 44994 51378
rect 44994 51326 44996 51378
rect 44940 51324 44996 51326
rect 43260 50764 43316 50820
rect 44156 51100 44212 51156
rect 43596 49756 43652 49812
rect 43820 49698 43876 49700
rect 43820 49646 43822 49698
rect 43822 49646 43874 49698
rect 43874 49646 43876 49698
rect 43820 49644 43876 49646
rect 42028 48802 42084 48804
rect 42028 48750 42030 48802
rect 42030 48750 42082 48802
rect 42082 48750 42084 48802
rect 42028 48748 42084 48750
rect 42476 47570 42532 47572
rect 42476 47518 42478 47570
rect 42478 47518 42530 47570
rect 42530 47518 42532 47570
rect 42476 47516 42532 47518
rect 41580 47458 41636 47460
rect 41580 47406 41582 47458
rect 41582 47406 41634 47458
rect 41634 47406 41636 47458
rect 41580 47404 41636 47406
rect 41132 46396 41188 46452
rect 41244 47292 41300 47348
rect 41804 47292 41860 47348
rect 41804 46844 41860 46900
rect 41132 45612 41188 45668
rect 41692 45724 41748 45780
rect 41468 45388 41524 45444
rect 41356 45052 41412 45108
rect 41356 44380 41412 44436
rect 41244 44322 41300 44324
rect 41244 44270 41246 44322
rect 41246 44270 41298 44322
rect 41298 44270 41300 44322
rect 41244 44268 41300 44270
rect 41580 44322 41636 44324
rect 41580 44270 41582 44322
rect 41582 44270 41634 44322
rect 41634 44270 41636 44322
rect 41580 44268 41636 44270
rect 41580 43538 41636 43540
rect 41580 43486 41582 43538
rect 41582 43486 41634 43538
rect 41634 43486 41636 43538
rect 41580 43484 41636 43486
rect 41356 42530 41412 42532
rect 41356 42478 41358 42530
rect 41358 42478 41410 42530
rect 41410 42478 41412 42530
rect 41356 42476 41412 42478
rect 40908 41916 40964 41972
rect 39900 40908 39956 40964
rect 40684 40572 40740 40628
rect 40012 40460 40068 40516
rect 40236 40178 40292 40180
rect 40236 40126 40238 40178
rect 40238 40126 40290 40178
rect 40290 40126 40292 40178
rect 40236 40124 40292 40126
rect 40796 40124 40852 40180
rect 40460 39730 40516 39732
rect 40460 39678 40462 39730
rect 40462 39678 40514 39730
rect 40514 39678 40516 39730
rect 40460 39676 40516 39678
rect 40796 38946 40852 38948
rect 40796 38894 40798 38946
rect 40798 38894 40850 38946
rect 40850 38894 40852 38946
rect 40796 38892 40852 38894
rect 39676 37660 39732 37716
rect 39564 37548 39620 37604
rect 40124 38162 40180 38164
rect 40124 38110 40126 38162
rect 40126 38110 40178 38162
rect 40178 38110 40180 38162
rect 40124 38108 40180 38110
rect 41244 40962 41300 40964
rect 41244 40910 41246 40962
rect 41246 40910 41298 40962
rect 41298 40910 41300 40962
rect 41244 40908 41300 40910
rect 41468 40572 41524 40628
rect 41132 40124 41188 40180
rect 41580 39618 41636 39620
rect 41580 39566 41582 39618
rect 41582 39566 41634 39618
rect 41634 39566 41636 39618
rect 41580 39564 41636 39566
rect 41804 43260 41860 43316
rect 42140 45890 42196 45892
rect 42140 45838 42142 45890
rect 42142 45838 42194 45890
rect 42194 45838 42196 45890
rect 42140 45836 42196 45838
rect 41804 42530 41860 42532
rect 41804 42478 41806 42530
rect 41806 42478 41858 42530
rect 41858 42478 41860 42530
rect 41804 42476 41860 42478
rect 41804 40962 41860 40964
rect 41804 40910 41806 40962
rect 41806 40910 41858 40962
rect 41858 40910 41860 40962
rect 41804 40908 41860 40910
rect 42812 45890 42868 45892
rect 42812 45838 42814 45890
rect 42814 45838 42866 45890
rect 42866 45838 42868 45890
rect 42812 45836 42868 45838
rect 42588 45724 42644 45780
rect 42476 45612 42532 45668
rect 42252 45106 42308 45108
rect 42252 45054 42254 45106
rect 42254 45054 42306 45106
rect 42306 45054 42308 45106
rect 42252 45052 42308 45054
rect 42252 43538 42308 43540
rect 42252 43486 42254 43538
rect 42254 43486 42306 43538
rect 42306 43486 42308 43538
rect 42252 43484 42308 43486
rect 42028 41468 42084 41524
rect 42140 42364 42196 42420
rect 42252 42140 42308 42196
rect 42364 42476 42420 42532
rect 42140 40796 42196 40852
rect 43260 47516 43316 47572
rect 43820 48860 43876 48916
rect 43596 48802 43652 48804
rect 43596 48750 43598 48802
rect 43598 48750 43650 48802
rect 43650 48750 43652 48802
rect 43596 48748 43652 48750
rect 44044 47292 44100 47348
rect 43036 45778 43092 45780
rect 43036 45726 43038 45778
rect 43038 45726 43090 45778
rect 43090 45726 43092 45778
rect 43036 45724 43092 45726
rect 43596 45218 43652 45220
rect 43596 45166 43598 45218
rect 43598 45166 43650 45218
rect 43650 45166 43652 45218
rect 43596 45164 43652 45166
rect 42588 44322 42644 44324
rect 42588 44270 42590 44322
rect 42590 44270 42642 44322
rect 42642 44270 42644 44322
rect 42588 44268 42644 44270
rect 42924 44268 42980 44324
rect 43484 44210 43540 44212
rect 43484 44158 43486 44210
rect 43486 44158 43538 44210
rect 43538 44158 43540 44210
rect 43484 44156 43540 44158
rect 43596 43708 43652 43764
rect 43932 43484 43988 43540
rect 45052 51154 45108 51156
rect 45052 51102 45054 51154
rect 45054 51102 45106 51154
rect 45106 51102 45108 51154
rect 45052 51100 45108 51102
rect 44604 50316 44660 50372
rect 45164 49644 45220 49700
rect 44716 49026 44772 49028
rect 44716 48974 44718 49026
rect 44718 48974 44770 49026
rect 44770 48974 44772 49026
rect 44716 48972 44772 48974
rect 44604 48802 44660 48804
rect 44604 48750 44606 48802
rect 44606 48750 44658 48802
rect 44658 48750 44660 48802
rect 44604 48748 44660 48750
rect 44604 47458 44660 47460
rect 44604 47406 44606 47458
rect 44606 47406 44658 47458
rect 44658 47406 44660 47458
rect 44604 47404 44660 47406
rect 44716 46732 44772 46788
rect 44156 45666 44212 45668
rect 44156 45614 44158 45666
rect 44158 45614 44210 45666
rect 44210 45614 44212 45666
rect 44156 45612 44212 45614
rect 46284 51100 46340 51156
rect 47404 51436 47460 51492
rect 47180 51378 47236 51380
rect 47180 51326 47182 51378
rect 47182 51326 47234 51378
rect 47234 51326 47236 51378
rect 47180 51324 47236 51326
rect 47068 51100 47124 51156
rect 48748 53900 48804 53956
rect 50092 53676 50148 53732
rect 48636 52780 48692 52836
rect 47404 50540 47460 50596
rect 45836 50316 45892 50372
rect 46060 50370 46116 50372
rect 46060 50318 46062 50370
rect 46062 50318 46114 50370
rect 46114 50318 46116 50370
rect 46060 50316 46116 50318
rect 46956 50370 47012 50372
rect 46956 50318 46958 50370
rect 46958 50318 47010 50370
rect 47010 50318 47012 50370
rect 46956 50316 47012 50318
rect 45724 48972 45780 49028
rect 47180 49250 47236 49252
rect 47180 49198 47182 49250
rect 47182 49198 47234 49250
rect 47234 49198 47236 49250
rect 47180 49196 47236 49198
rect 46060 48860 46116 48916
rect 46732 48860 46788 48916
rect 46172 48242 46228 48244
rect 46172 48190 46174 48242
rect 46174 48190 46226 48242
rect 46226 48190 46228 48242
rect 46172 48188 46228 48190
rect 46060 47516 46116 47572
rect 45388 47458 45444 47460
rect 45388 47406 45390 47458
rect 45390 47406 45442 47458
rect 45442 47406 45444 47458
rect 45388 47404 45444 47406
rect 45164 45836 45220 45892
rect 44492 45724 44548 45780
rect 45052 45388 45108 45444
rect 45276 46956 45332 47012
rect 44268 45218 44324 45220
rect 44268 45166 44270 45218
rect 44270 45166 44322 45218
rect 44322 45166 44324 45218
rect 44268 45164 44324 45166
rect 44268 44434 44324 44436
rect 44268 44382 44270 44434
rect 44270 44382 44322 44434
rect 44322 44382 44324 44434
rect 44268 44380 44324 44382
rect 46844 48188 46900 48244
rect 46732 47570 46788 47572
rect 46732 47518 46734 47570
rect 46734 47518 46786 47570
rect 46786 47518 46788 47570
rect 46732 47516 46788 47518
rect 45836 47346 45892 47348
rect 45836 47294 45838 47346
rect 45838 47294 45890 47346
rect 45890 47294 45892 47346
rect 45836 47292 45892 47294
rect 45500 46786 45556 46788
rect 45500 46734 45502 46786
rect 45502 46734 45554 46786
rect 45554 46734 45556 46786
rect 45500 46732 45556 46734
rect 47180 47068 47236 47124
rect 45500 45778 45556 45780
rect 45500 45726 45502 45778
rect 45502 45726 45554 45778
rect 45554 45726 45556 45778
rect 45500 45724 45556 45726
rect 45948 45890 46004 45892
rect 45948 45838 45950 45890
rect 45950 45838 46002 45890
rect 46002 45838 46004 45890
rect 45948 45836 46004 45838
rect 45724 45388 45780 45444
rect 44604 44044 44660 44100
rect 42476 42364 42532 42420
rect 44716 43596 44772 43652
rect 42700 42364 42756 42420
rect 44716 42530 44772 42532
rect 44716 42478 44718 42530
rect 44718 42478 44770 42530
rect 44770 42478 44772 42530
rect 44716 42476 44772 42478
rect 43148 41858 43204 41860
rect 43148 41806 43150 41858
rect 43150 41806 43202 41858
rect 43202 41806 43204 41858
rect 43148 41804 43204 41806
rect 43372 41970 43428 41972
rect 43372 41918 43374 41970
rect 43374 41918 43426 41970
rect 43426 41918 43428 41970
rect 43372 41916 43428 41918
rect 43260 41468 43316 41524
rect 43820 41858 43876 41860
rect 43820 41806 43822 41858
rect 43822 41806 43874 41858
rect 43874 41806 43876 41858
rect 43820 41804 43876 41806
rect 43820 41244 43876 41300
rect 43596 41074 43652 41076
rect 43596 41022 43598 41074
rect 43598 41022 43650 41074
rect 43650 41022 43652 41074
rect 43596 41020 43652 41022
rect 42700 40684 42756 40740
rect 43036 40908 43092 40964
rect 42476 40572 42532 40628
rect 42140 39676 42196 39732
rect 40908 38108 40964 38164
rect 40236 38050 40292 38052
rect 40236 37998 40238 38050
rect 40238 37998 40290 38050
rect 40290 37998 40292 38050
rect 40236 37996 40292 37998
rect 39340 37436 39396 37492
rect 39900 37436 39956 37492
rect 39228 35532 39284 35588
rect 39116 34860 39172 34916
rect 39004 34636 39060 34692
rect 39676 36988 39732 37044
rect 39564 36316 39620 36372
rect 39900 36988 39956 37044
rect 40236 37660 40292 37716
rect 39900 36204 39956 36260
rect 39564 35474 39620 35476
rect 39564 35422 39566 35474
rect 39566 35422 39618 35474
rect 39618 35422 39620 35474
rect 39564 35420 39620 35422
rect 39452 34130 39508 34132
rect 39452 34078 39454 34130
rect 39454 34078 39506 34130
rect 39506 34078 39508 34130
rect 39452 34076 39508 34078
rect 39116 33570 39172 33572
rect 39116 33518 39118 33570
rect 39118 33518 39170 33570
rect 39170 33518 39172 33570
rect 39116 33516 39172 33518
rect 39340 33740 39396 33796
rect 39004 33180 39060 33236
rect 38332 32674 38388 32676
rect 38332 32622 38334 32674
rect 38334 32622 38386 32674
rect 38386 32622 38388 32674
rect 38332 32620 38388 32622
rect 37772 31666 37828 31668
rect 37772 31614 37774 31666
rect 37774 31614 37826 31666
rect 37826 31614 37828 31666
rect 37772 31612 37828 31614
rect 38108 31948 38164 32004
rect 37660 31388 37716 31444
rect 37324 29708 37380 29764
rect 37436 29484 37492 29540
rect 36988 26236 37044 26292
rect 36988 25564 37044 25620
rect 37324 28700 37380 28756
rect 36764 23826 36820 23828
rect 36764 23774 36766 23826
rect 36766 23774 36818 23826
rect 36818 23774 36820 23826
rect 36764 23772 36820 23774
rect 36876 23660 36932 23716
rect 36764 23548 36820 23604
rect 37212 26460 37268 26516
rect 36988 23266 37044 23268
rect 36988 23214 36990 23266
rect 36990 23214 37042 23266
rect 37042 23214 37044 23266
rect 36988 23212 37044 23214
rect 38556 32562 38612 32564
rect 38556 32510 38558 32562
rect 38558 32510 38610 32562
rect 38610 32510 38612 32562
rect 38556 32508 38612 32510
rect 38444 32396 38500 32452
rect 38220 31276 38276 31332
rect 38332 31388 38388 31444
rect 38108 31218 38164 31220
rect 38108 31166 38110 31218
rect 38110 31166 38162 31218
rect 38162 31166 38164 31218
rect 38108 31164 38164 31166
rect 38332 30268 38388 30324
rect 37884 29596 37940 29652
rect 38220 29260 38276 29316
rect 38332 29202 38388 29204
rect 38332 29150 38334 29202
rect 38334 29150 38386 29202
rect 38386 29150 38388 29202
rect 38332 29148 38388 29150
rect 38220 28588 38276 28644
rect 37548 28364 37604 28420
rect 38108 28476 38164 28532
rect 37660 27468 37716 27524
rect 37436 25618 37492 25620
rect 37436 25566 37438 25618
rect 37438 25566 37490 25618
rect 37490 25566 37492 25618
rect 37436 25564 37492 25566
rect 37884 25394 37940 25396
rect 37884 25342 37886 25394
rect 37886 25342 37938 25394
rect 37938 25342 37940 25394
rect 37884 25340 37940 25342
rect 37324 23436 37380 23492
rect 37772 24444 37828 24500
rect 37772 24050 37828 24052
rect 37772 23998 37774 24050
rect 37774 23998 37826 24050
rect 37826 23998 37828 24050
rect 37772 23996 37828 23998
rect 37548 23938 37604 23940
rect 37548 23886 37550 23938
rect 37550 23886 37602 23938
rect 37602 23886 37604 23938
rect 37548 23884 37604 23886
rect 36540 22316 36596 22372
rect 36764 21644 36820 21700
rect 35756 19740 35812 19796
rect 36092 19740 36148 19796
rect 36764 21084 36820 21140
rect 36652 20748 36708 20804
rect 36540 20524 36596 20580
rect 36540 20130 36596 20132
rect 36540 20078 36542 20130
rect 36542 20078 36594 20130
rect 36594 20078 36596 20130
rect 36540 20076 36596 20078
rect 36428 19740 36484 19796
rect 36764 20130 36820 20132
rect 36764 20078 36766 20130
rect 36766 20078 36818 20130
rect 36818 20078 36820 20130
rect 36764 20076 36820 20078
rect 36876 19964 36932 20020
rect 36204 19234 36260 19236
rect 36204 19182 36206 19234
rect 36206 19182 36258 19234
rect 36258 19182 36260 19234
rect 36204 19180 36260 19182
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35868 17666 35924 17668
rect 35868 17614 35870 17666
rect 35870 17614 35922 17666
rect 35922 17614 35924 17666
rect 35868 17612 35924 17614
rect 36092 18450 36148 18452
rect 36092 18398 36094 18450
rect 36094 18398 36146 18450
rect 36146 18398 36148 18450
rect 36092 18396 36148 18398
rect 36652 17836 36708 17892
rect 34860 17164 34916 17220
rect 34748 16210 34804 16212
rect 34748 16158 34750 16210
rect 34750 16158 34802 16210
rect 34802 16158 34804 16210
rect 34748 16156 34804 16158
rect 34860 15372 34916 15428
rect 35308 17500 35364 17556
rect 35084 17052 35140 17108
rect 35644 17554 35700 17556
rect 35644 17502 35646 17554
rect 35646 17502 35698 17554
rect 35698 17502 35700 17554
rect 35644 17500 35700 17502
rect 35980 17442 36036 17444
rect 35980 17390 35982 17442
rect 35982 17390 36034 17442
rect 36034 17390 36036 17442
rect 35980 17388 36036 17390
rect 36092 17052 36148 17108
rect 35532 16882 35588 16884
rect 35532 16830 35534 16882
rect 35534 16830 35586 16882
rect 35586 16830 35588 16882
rect 35532 16828 35588 16830
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35420 16156 35476 16212
rect 35756 16044 35812 16100
rect 35084 15260 35140 15316
rect 35644 15820 35700 15876
rect 35868 15372 35924 15428
rect 35980 15484 36036 15540
rect 36204 16604 36260 16660
rect 36764 17554 36820 17556
rect 36764 17502 36766 17554
rect 36766 17502 36818 17554
rect 36818 17502 36820 17554
rect 36764 17500 36820 17502
rect 36540 16994 36596 16996
rect 36540 16942 36542 16994
rect 36542 16942 36594 16994
rect 36594 16942 36596 16994
rect 36540 16940 36596 16942
rect 36428 15986 36484 15988
rect 36428 15934 36430 15986
rect 36430 15934 36482 15986
rect 36482 15934 36484 15986
rect 36428 15932 36484 15934
rect 36204 15484 36260 15540
rect 36204 15314 36260 15316
rect 36204 15262 36206 15314
rect 36206 15262 36258 15314
rect 36258 15262 36260 15314
rect 36204 15260 36260 15262
rect 35420 15036 35476 15092
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35756 14924 35812 14980
rect 34524 14530 34580 14532
rect 34524 14478 34526 14530
rect 34526 14478 34578 14530
rect 34578 14478 34580 14530
rect 34524 14476 34580 14478
rect 34636 13858 34692 13860
rect 34636 13806 34638 13858
rect 34638 13806 34690 13858
rect 34690 13806 34692 13858
rect 34636 13804 34692 13806
rect 34636 13580 34692 13636
rect 34188 11394 34244 11396
rect 34188 11342 34190 11394
rect 34190 11342 34242 11394
rect 34242 11342 34244 11394
rect 34188 11340 34244 11342
rect 33740 11004 33796 11060
rect 33516 10556 33572 10612
rect 34188 11004 34244 11060
rect 33516 9938 33572 9940
rect 33516 9886 33518 9938
rect 33518 9886 33570 9938
rect 33570 9886 33572 9938
rect 33516 9884 33572 9886
rect 33292 8428 33348 8484
rect 33628 8316 33684 8372
rect 33740 8204 33796 8260
rect 32956 6636 33012 6692
rect 32508 5906 32564 5908
rect 32508 5854 32510 5906
rect 32510 5854 32562 5906
rect 32562 5854 32564 5906
rect 32508 5852 32564 5854
rect 31612 5516 31668 5572
rect 30940 4844 30996 4900
rect 31836 4898 31892 4900
rect 31836 4846 31838 4898
rect 31838 4846 31890 4898
rect 31890 4846 31892 4898
rect 31836 4844 31892 4846
rect 30828 4508 30884 4564
rect 31500 4508 31556 4564
rect 29820 4396 29876 4452
rect 29708 4284 29764 4340
rect 33068 6412 33124 6468
rect 31948 4396 32004 4452
rect 32844 4562 32900 4564
rect 32844 4510 32846 4562
rect 32846 4510 32898 4562
rect 32898 4510 32900 4562
rect 32844 4508 32900 4510
rect 29708 3724 29764 3780
rect 30716 3724 30772 3780
rect 29260 3554 29316 3556
rect 29260 3502 29262 3554
rect 29262 3502 29314 3554
rect 29314 3502 29316 3554
rect 29260 3500 29316 3502
rect 27244 3442 27300 3444
rect 27244 3390 27246 3442
rect 27246 3390 27298 3442
rect 27298 3390 27300 3442
rect 27244 3388 27300 3390
rect 30156 3388 30212 3444
rect 14476 3276 14532 3332
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 30380 3442 30436 3444
rect 30380 3390 30382 3442
rect 30382 3390 30434 3442
rect 30434 3390 30436 3442
rect 30380 3388 30436 3390
rect 31612 3612 31668 3668
rect 33740 6466 33796 6468
rect 33740 6414 33742 6466
rect 33742 6414 33794 6466
rect 33794 6414 33796 6466
rect 33740 6412 33796 6414
rect 33180 6076 33236 6132
rect 33852 5906 33908 5908
rect 33852 5854 33854 5906
rect 33854 5854 33906 5906
rect 33906 5854 33908 5906
rect 33852 5852 33908 5854
rect 33628 5180 33684 5236
rect 33068 3724 33124 3780
rect 32284 3666 32340 3668
rect 32284 3614 32286 3666
rect 32286 3614 32338 3666
rect 32338 3614 32340 3666
rect 32284 3612 32340 3614
rect 34636 12178 34692 12180
rect 34636 12126 34638 12178
rect 34638 12126 34690 12178
rect 34690 12126 34692 12178
rect 34636 12124 34692 12126
rect 34748 11340 34804 11396
rect 34300 10722 34356 10724
rect 34300 10670 34302 10722
rect 34302 10670 34354 10722
rect 34354 10670 34356 10722
rect 34300 10668 34356 10670
rect 34076 9884 34132 9940
rect 34412 9772 34468 9828
rect 34076 8370 34132 8372
rect 34076 8318 34078 8370
rect 34078 8318 34130 8370
rect 34130 8318 34132 8370
rect 34076 8316 34132 8318
rect 34300 8258 34356 8260
rect 34300 8206 34302 8258
rect 34302 8206 34354 8258
rect 34354 8206 34356 8258
rect 34300 8204 34356 8206
rect 34188 6636 34244 6692
rect 34636 9884 34692 9940
rect 35084 14476 35140 14532
rect 35308 14700 35364 14756
rect 35420 13858 35476 13860
rect 35420 13806 35422 13858
rect 35422 13806 35474 13858
rect 35474 13806 35476 13858
rect 35420 13804 35476 13806
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35420 12402 35476 12404
rect 35420 12350 35422 12402
rect 35422 12350 35474 12402
rect 35474 12350 35476 12402
rect 35420 12348 35476 12350
rect 34972 12290 35028 12292
rect 34972 12238 34974 12290
rect 34974 12238 35026 12290
rect 35026 12238 35028 12290
rect 34972 12236 35028 12238
rect 35532 12236 35588 12292
rect 35644 12124 35700 12180
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35420 10668 35476 10724
rect 35308 10610 35364 10612
rect 35308 10558 35310 10610
rect 35310 10558 35362 10610
rect 35362 10558 35364 10610
rect 35308 10556 35364 10558
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35084 9884 35140 9940
rect 35308 9826 35364 9828
rect 35308 9774 35310 9826
rect 35310 9774 35362 9826
rect 35362 9774 35364 9826
rect 35308 9772 35364 9774
rect 34972 9714 35028 9716
rect 34972 9662 34974 9714
rect 34974 9662 35026 9714
rect 35026 9662 35028 9714
rect 34972 9660 35028 9662
rect 36316 14924 36372 14980
rect 36764 15484 36820 15540
rect 36764 14700 36820 14756
rect 36316 14418 36372 14420
rect 36316 14366 36318 14418
rect 36318 14366 36370 14418
rect 36370 14366 36372 14418
rect 36316 14364 36372 14366
rect 38668 32396 38724 32452
rect 38556 32284 38612 32340
rect 38780 31612 38836 31668
rect 38892 32844 38948 32900
rect 39116 32844 39172 32900
rect 39564 33180 39620 33236
rect 39900 35698 39956 35700
rect 39900 35646 39902 35698
rect 39902 35646 39954 35698
rect 39954 35646 39956 35698
rect 39900 35644 39956 35646
rect 40124 35420 40180 35476
rect 39900 34690 39956 34692
rect 39900 34638 39902 34690
rect 39902 34638 39954 34690
rect 39954 34638 39956 34690
rect 39900 34636 39956 34638
rect 39676 32844 39732 32900
rect 39900 34242 39956 34244
rect 39900 34190 39902 34242
rect 39902 34190 39954 34242
rect 39954 34190 39956 34242
rect 39900 34188 39956 34190
rect 39340 32732 39396 32788
rect 39228 32562 39284 32564
rect 39228 32510 39230 32562
rect 39230 32510 39282 32562
rect 39282 32510 39284 32562
rect 39228 32508 39284 32510
rect 39116 31388 39172 31444
rect 39116 31106 39172 31108
rect 39116 31054 39118 31106
rect 39118 31054 39170 31106
rect 39170 31054 39172 31106
rect 39116 31052 39172 31054
rect 39228 30882 39284 30884
rect 39228 30830 39230 30882
rect 39230 30830 39282 30882
rect 39282 30830 39284 30882
rect 39228 30828 39284 30830
rect 38780 30604 38836 30660
rect 38892 29932 38948 29988
rect 38892 29708 38948 29764
rect 38780 28364 38836 28420
rect 38556 27804 38612 27860
rect 38668 27580 38724 27636
rect 38668 27132 38724 27188
rect 38780 26684 38836 26740
rect 38556 26514 38612 26516
rect 38556 26462 38558 26514
rect 38558 26462 38610 26514
rect 38610 26462 38612 26514
rect 38556 26460 38612 26462
rect 38780 26460 38836 26516
rect 40012 33740 40068 33796
rect 40572 37154 40628 37156
rect 40572 37102 40574 37154
rect 40574 37102 40626 37154
rect 40626 37102 40628 37154
rect 40572 37100 40628 37102
rect 40460 35474 40516 35476
rect 40460 35422 40462 35474
rect 40462 35422 40514 35474
rect 40514 35422 40516 35474
rect 40460 35420 40516 35422
rect 40460 33740 40516 33796
rect 39900 33068 39956 33124
rect 40236 33404 40292 33460
rect 40124 33122 40180 33124
rect 40124 33070 40126 33122
rect 40126 33070 40178 33122
rect 40178 33070 40180 33122
rect 40124 33068 40180 33070
rect 40236 32732 40292 32788
rect 40012 32396 40068 32452
rect 39452 31388 39508 31444
rect 40796 35644 40852 35700
rect 41468 37490 41524 37492
rect 41468 37438 41470 37490
rect 41470 37438 41522 37490
rect 41522 37438 41524 37490
rect 41468 37436 41524 37438
rect 41356 36482 41412 36484
rect 41356 36430 41358 36482
rect 41358 36430 41410 36482
rect 41410 36430 41412 36482
rect 41356 36428 41412 36430
rect 42028 39058 42084 39060
rect 42028 39006 42030 39058
rect 42030 39006 42082 39058
rect 42082 39006 42084 39058
rect 42028 39004 42084 39006
rect 42140 36876 42196 36932
rect 41692 36594 41748 36596
rect 41692 36542 41694 36594
rect 41694 36542 41746 36594
rect 41746 36542 41748 36594
rect 41692 36540 41748 36542
rect 41132 35644 41188 35700
rect 41804 36428 41860 36484
rect 42252 36258 42308 36260
rect 42252 36206 42254 36258
rect 42254 36206 42306 36258
rect 42306 36206 42308 36258
rect 42252 36204 42308 36206
rect 43148 40684 43204 40740
rect 43708 40796 43764 40852
rect 43708 40348 43764 40404
rect 44604 41020 44660 41076
rect 44268 40402 44324 40404
rect 44268 40350 44270 40402
rect 44270 40350 44322 40402
rect 44322 40350 44324 40402
rect 44268 40348 44324 40350
rect 42588 39730 42644 39732
rect 42588 39678 42590 39730
rect 42590 39678 42642 39730
rect 42642 39678 42644 39730
rect 42588 39676 42644 39678
rect 42812 39004 42868 39060
rect 42924 39564 42980 39620
rect 43148 39564 43204 39620
rect 45052 40348 45108 40404
rect 44716 39506 44772 39508
rect 44716 39454 44718 39506
rect 44718 39454 44770 39506
rect 44770 39454 44772 39506
rect 44716 39452 44772 39454
rect 44268 38892 44324 38948
rect 44492 38780 44548 38836
rect 42924 38668 42980 38724
rect 43708 38668 43764 38724
rect 42700 37154 42756 37156
rect 42700 37102 42702 37154
rect 42702 37102 42754 37154
rect 42754 37102 42756 37154
rect 42700 37100 42756 37102
rect 42588 36876 42644 36932
rect 43372 37154 43428 37156
rect 43372 37102 43374 37154
rect 43374 37102 43426 37154
rect 43426 37102 43428 37154
rect 43372 37100 43428 37102
rect 42476 35980 42532 36036
rect 42700 35868 42756 35924
rect 41804 35756 41860 35812
rect 40796 35026 40852 35028
rect 40796 34974 40798 35026
rect 40798 34974 40850 35026
rect 40850 34974 40852 35026
rect 40796 34972 40852 34974
rect 40796 34242 40852 34244
rect 40796 34190 40798 34242
rect 40798 34190 40850 34242
rect 40850 34190 40852 34242
rect 40796 34188 40852 34190
rect 41244 34188 41300 34244
rect 40908 33234 40964 33236
rect 40908 33182 40910 33234
rect 40910 33182 40962 33234
rect 40962 33182 40964 33234
rect 40908 33180 40964 33182
rect 41020 33122 41076 33124
rect 41020 33070 41022 33122
rect 41022 33070 41074 33122
rect 41074 33070 41076 33122
rect 41020 33068 41076 33070
rect 40684 32284 40740 32340
rect 40012 31890 40068 31892
rect 40012 31838 40014 31890
rect 40014 31838 40066 31890
rect 40066 31838 40068 31890
rect 40012 31836 40068 31838
rect 40236 31836 40292 31892
rect 39788 31388 39844 31444
rect 40012 30828 40068 30884
rect 40012 30044 40068 30100
rect 40012 28866 40068 28868
rect 40012 28814 40014 28866
rect 40014 28814 40066 28866
rect 40066 28814 40068 28866
rect 40012 28812 40068 28814
rect 40572 31276 40628 31332
rect 40796 30828 40852 30884
rect 40348 30268 40404 30324
rect 40572 30098 40628 30100
rect 40572 30046 40574 30098
rect 40574 30046 40626 30098
rect 40626 30046 40628 30098
rect 40572 30044 40628 30046
rect 40460 29426 40516 29428
rect 40460 29374 40462 29426
rect 40462 29374 40514 29426
rect 40514 29374 40516 29426
rect 40460 29372 40516 29374
rect 40572 29036 40628 29092
rect 40684 28812 40740 28868
rect 40796 28754 40852 28756
rect 40796 28702 40798 28754
rect 40798 28702 40850 28754
rect 40850 28702 40852 28754
rect 40796 28700 40852 28702
rect 39676 28530 39732 28532
rect 39676 28478 39678 28530
rect 39678 28478 39730 28530
rect 39730 28478 39732 28530
rect 39676 28476 39732 28478
rect 39116 27244 39172 27300
rect 39452 27244 39508 27300
rect 39228 27132 39284 27188
rect 39004 26796 39060 26852
rect 39340 26908 39396 26964
rect 39564 27020 39620 27076
rect 39900 28140 39956 28196
rect 40236 28140 40292 28196
rect 40012 27580 40068 27636
rect 40236 27356 40292 27412
rect 38892 25900 38948 25956
rect 38780 24722 38836 24724
rect 38780 24670 38782 24722
rect 38782 24670 38834 24722
rect 38834 24670 38836 24722
rect 38780 24668 38836 24670
rect 38220 23996 38276 24052
rect 38332 23938 38388 23940
rect 38332 23886 38334 23938
rect 38334 23886 38386 23938
rect 38386 23886 38388 23938
rect 38332 23884 38388 23886
rect 38220 23826 38276 23828
rect 38220 23774 38222 23826
rect 38222 23774 38274 23826
rect 38274 23774 38276 23826
rect 38220 23772 38276 23774
rect 37324 22092 37380 22148
rect 37212 21810 37268 21812
rect 37212 21758 37214 21810
rect 37214 21758 37266 21810
rect 37266 21758 37268 21810
rect 37212 21756 37268 21758
rect 37100 21586 37156 21588
rect 37100 21534 37102 21586
rect 37102 21534 37154 21586
rect 37154 21534 37156 21586
rect 37100 21532 37156 21534
rect 37548 20802 37604 20804
rect 37548 20750 37550 20802
rect 37550 20750 37602 20802
rect 37602 20750 37604 20802
rect 37548 20748 37604 20750
rect 37548 20130 37604 20132
rect 37548 20078 37550 20130
rect 37550 20078 37602 20130
rect 37602 20078 37604 20130
rect 37548 20076 37604 20078
rect 37324 18620 37380 18676
rect 37436 18508 37492 18564
rect 38444 23714 38500 23716
rect 38444 23662 38446 23714
rect 38446 23662 38498 23714
rect 38498 23662 38500 23714
rect 38444 23660 38500 23662
rect 37996 22988 38052 23044
rect 37884 21868 37940 21924
rect 38220 21810 38276 21812
rect 38220 21758 38222 21810
rect 38222 21758 38274 21810
rect 38274 21758 38276 21810
rect 38220 21756 38276 21758
rect 38108 20860 38164 20916
rect 38780 23042 38836 23044
rect 38780 22990 38782 23042
rect 38782 22990 38834 23042
rect 38834 22990 38836 23042
rect 38780 22988 38836 22990
rect 38780 21756 38836 21812
rect 39004 26236 39060 26292
rect 39228 25676 39284 25732
rect 39228 25282 39284 25284
rect 39228 25230 39230 25282
rect 39230 25230 39282 25282
rect 39282 25230 39284 25282
rect 39228 25228 39284 25230
rect 39004 23772 39060 23828
rect 39452 24108 39508 24164
rect 39676 25788 39732 25844
rect 39340 22482 39396 22484
rect 39340 22430 39342 22482
rect 39342 22430 39394 22482
rect 39394 22430 39396 22482
rect 39340 22428 39396 22430
rect 39228 21980 39284 22036
rect 39116 21868 39172 21924
rect 38556 20578 38612 20580
rect 38556 20526 38558 20578
rect 38558 20526 38610 20578
rect 38610 20526 38612 20578
rect 38556 20524 38612 20526
rect 38668 20860 38724 20916
rect 37996 20188 38052 20244
rect 38892 21362 38948 21364
rect 38892 21310 38894 21362
rect 38894 21310 38946 21362
rect 38946 21310 38948 21362
rect 38892 21308 38948 21310
rect 39228 21586 39284 21588
rect 39228 21534 39230 21586
rect 39230 21534 39282 21586
rect 39282 21534 39284 21586
rect 39228 21532 39284 21534
rect 39004 20300 39060 20356
rect 37884 19234 37940 19236
rect 37884 19182 37886 19234
rect 37886 19182 37938 19234
rect 37938 19182 37940 19234
rect 37884 19180 37940 19182
rect 37436 17836 37492 17892
rect 37660 17890 37716 17892
rect 37660 17838 37662 17890
rect 37662 17838 37714 17890
rect 37714 17838 37716 17890
rect 37660 17836 37716 17838
rect 39228 21196 39284 21252
rect 39004 18562 39060 18564
rect 39004 18510 39006 18562
rect 39006 18510 39058 18562
rect 39058 18510 39060 18562
rect 39004 18508 39060 18510
rect 37772 17500 37828 17556
rect 38332 17724 38388 17780
rect 37884 17442 37940 17444
rect 37884 17390 37886 17442
rect 37886 17390 37938 17442
rect 37938 17390 37940 17442
rect 37884 17388 37940 17390
rect 38892 17778 38948 17780
rect 38892 17726 38894 17778
rect 38894 17726 38946 17778
rect 38946 17726 38948 17778
rect 38892 17724 38948 17726
rect 39116 17724 39172 17780
rect 39004 17164 39060 17220
rect 37548 16716 37604 16772
rect 39116 16380 39172 16436
rect 37436 16210 37492 16212
rect 37436 16158 37438 16210
rect 37438 16158 37490 16210
rect 37490 16158 37492 16210
rect 37436 16156 37492 16158
rect 37884 16210 37940 16212
rect 37884 16158 37886 16210
rect 37886 16158 37938 16210
rect 37938 16158 37940 16210
rect 37884 16156 37940 16158
rect 38444 16210 38500 16212
rect 38444 16158 38446 16210
rect 38446 16158 38498 16210
rect 38498 16158 38500 16210
rect 38444 16156 38500 16158
rect 38108 15484 38164 15540
rect 37436 15426 37492 15428
rect 37436 15374 37438 15426
rect 37438 15374 37490 15426
rect 37490 15374 37492 15426
rect 37436 15372 37492 15374
rect 37996 15426 38052 15428
rect 37996 15374 37998 15426
rect 37998 15374 38050 15426
rect 38050 15374 38052 15426
rect 37996 15372 38052 15374
rect 37212 15314 37268 15316
rect 37212 15262 37214 15314
rect 37214 15262 37266 15314
rect 37266 15262 37268 15314
rect 37212 15260 37268 15262
rect 37772 14924 37828 14980
rect 39116 16156 39172 16212
rect 39004 16098 39060 16100
rect 39004 16046 39006 16098
rect 39006 16046 39058 16098
rect 39058 16046 39060 16098
rect 39004 16044 39060 16046
rect 39676 23154 39732 23156
rect 39676 23102 39678 23154
rect 39678 23102 39730 23154
rect 39730 23102 39732 23154
rect 39676 23100 39732 23102
rect 40124 26290 40180 26292
rect 40124 26238 40126 26290
rect 40126 26238 40178 26290
rect 40178 26238 40180 26290
rect 40124 26236 40180 26238
rect 39900 26178 39956 26180
rect 39900 26126 39902 26178
rect 39902 26126 39954 26178
rect 39954 26126 39956 26178
rect 39900 26124 39956 26126
rect 40908 28476 40964 28532
rect 40572 27074 40628 27076
rect 40572 27022 40574 27074
rect 40574 27022 40626 27074
rect 40626 27022 40628 27074
rect 40572 27020 40628 27022
rect 41132 28252 41188 28308
rect 40908 26908 40964 26964
rect 41020 27580 41076 27636
rect 40460 26796 40516 26852
rect 40796 26850 40852 26852
rect 40796 26798 40798 26850
rect 40798 26798 40850 26850
rect 40850 26798 40852 26850
rect 40796 26796 40852 26798
rect 40348 26348 40404 26404
rect 40460 26514 40516 26516
rect 40460 26462 40462 26514
rect 40462 26462 40514 26514
rect 40514 26462 40516 26514
rect 40460 26460 40516 26462
rect 40236 25788 40292 25844
rect 40124 25676 40180 25732
rect 41020 26236 41076 26292
rect 40684 26012 40740 26068
rect 39900 24444 39956 24500
rect 41244 27692 41300 27748
rect 43484 35810 43540 35812
rect 43484 35758 43486 35810
rect 43486 35758 43538 35810
rect 43538 35758 43540 35810
rect 43484 35756 43540 35758
rect 42028 35698 42084 35700
rect 42028 35646 42030 35698
rect 42030 35646 42082 35698
rect 42082 35646 42084 35698
rect 42028 35644 42084 35646
rect 42476 35420 42532 35476
rect 41692 35138 41748 35140
rect 41692 35086 41694 35138
rect 41694 35086 41746 35138
rect 41746 35086 41748 35138
rect 41692 35084 41748 35086
rect 42028 34860 42084 34916
rect 41468 34130 41524 34132
rect 41468 34078 41470 34130
rect 41470 34078 41522 34130
rect 41522 34078 41524 34130
rect 41468 34076 41524 34078
rect 41916 33964 41972 34020
rect 42028 34636 42084 34692
rect 41468 33628 41524 33684
rect 41692 33516 41748 33572
rect 42364 34018 42420 34020
rect 42364 33966 42366 34018
rect 42366 33966 42418 34018
rect 42418 33966 42420 34018
rect 42364 33964 42420 33966
rect 43036 35420 43092 35476
rect 44156 38050 44212 38052
rect 44156 37998 44158 38050
rect 44158 37998 44210 38050
rect 44210 37998 44212 38050
rect 44156 37996 44212 37998
rect 44156 37154 44212 37156
rect 44156 37102 44158 37154
rect 44158 37102 44210 37154
rect 44210 37102 44212 37154
rect 44156 37100 44212 37102
rect 43820 36594 43876 36596
rect 43820 36542 43822 36594
rect 43822 36542 43874 36594
rect 43874 36542 43876 36594
rect 43820 36540 43876 36542
rect 44380 36540 44436 36596
rect 44156 36204 44212 36260
rect 43708 35308 43764 35364
rect 43932 35084 43988 35140
rect 42588 34914 42644 34916
rect 42588 34862 42590 34914
rect 42590 34862 42642 34914
rect 42642 34862 42644 34914
rect 42588 34860 42644 34862
rect 42700 34802 42756 34804
rect 42700 34750 42702 34802
rect 42702 34750 42754 34802
rect 42754 34750 42756 34802
rect 42700 34748 42756 34750
rect 42588 34242 42644 34244
rect 42588 34190 42590 34242
rect 42590 34190 42642 34242
rect 42642 34190 42644 34242
rect 42588 34188 42644 34190
rect 42812 34188 42868 34244
rect 43820 34690 43876 34692
rect 43820 34638 43822 34690
rect 43822 34638 43874 34690
rect 43874 34638 43876 34690
rect 43820 34636 43876 34638
rect 44044 34636 44100 34692
rect 43820 33964 43876 34020
rect 42140 32844 42196 32900
rect 41916 32562 41972 32564
rect 41916 32510 41918 32562
rect 41918 32510 41970 32562
rect 41970 32510 41972 32562
rect 41916 32508 41972 32510
rect 41916 31836 41972 31892
rect 41692 31612 41748 31668
rect 42252 31778 42308 31780
rect 42252 31726 42254 31778
rect 42254 31726 42306 31778
rect 42306 31726 42308 31778
rect 42252 31724 42308 31726
rect 42140 30882 42196 30884
rect 42140 30830 42142 30882
rect 42142 30830 42194 30882
rect 42194 30830 42196 30882
rect 42140 30828 42196 30830
rect 41804 30156 41860 30212
rect 42028 30044 42084 30100
rect 41692 29986 41748 29988
rect 41692 29934 41694 29986
rect 41694 29934 41746 29986
rect 41746 29934 41748 29986
rect 41692 29932 41748 29934
rect 41692 29426 41748 29428
rect 41692 29374 41694 29426
rect 41694 29374 41746 29426
rect 41746 29374 41748 29426
rect 41692 29372 41748 29374
rect 41580 29148 41636 29204
rect 41916 28812 41972 28868
rect 41916 28530 41972 28532
rect 41916 28478 41918 28530
rect 41918 28478 41970 28530
rect 41970 28478 41972 28530
rect 41916 28476 41972 28478
rect 43036 32620 43092 32676
rect 43820 32732 43876 32788
rect 42924 32562 42980 32564
rect 42924 32510 42926 32562
rect 42926 32510 42978 32562
rect 42978 32510 42980 32562
rect 42924 32508 42980 32510
rect 42588 31724 42644 31780
rect 42588 31052 42644 31108
rect 44044 32844 44100 32900
rect 43820 32284 43876 32340
rect 43596 31724 43652 31780
rect 43820 31948 43876 32004
rect 42700 31164 42756 31220
rect 42812 30828 42868 30884
rect 43820 31218 43876 31220
rect 43820 31166 43822 31218
rect 43822 31166 43874 31218
rect 43874 31166 43876 31218
rect 43820 31164 43876 31166
rect 43708 30882 43764 30884
rect 43708 30830 43710 30882
rect 43710 30830 43762 30882
rect 43762 30830 43764 30882
rect 43708 30828 43764 30830
rect 42924 30156 42980 30212
rect 43484 30098 43540 30100
rect 43484 30046 43486 30098
rect 43486 30046 43538 30098
rect 43538 30046 43540 30098
rect 43484 30044 43540 30046
rect 44380 35868 44436 35924
rect 44940 38834 44996 38836
rect 44940 38782 44942 38834
rect 44942 38782 44994 38834
rect 44994 38782 44996 38834
rect 44940 38780 44996 38782
rect 45724 44492 45780 44548
rect 46732 45052 46788 45108
rect 47068 45106 47124 45108
rect 47068 45054 47070 45106
rect 47070 45054 47122 45106
rect 47122 45054 47124 45106
rect 47068 45052 47124 45054
rect 45836 44434 45892 44436
rect 45836 44382 45838 44434
rect 45838 44382 45890 44434
rect 45890 44382 45892 44434
rect 45836 44380 45892 44382
rect 46172 44380 46228 44436
rect 47180 44604 47236 44660
rect 45276 43596 45332 43652
rect 45836 43372 45892 43428
rect 46060 43260 46116 43316
rect 46956 43426 47012 43428
rect 46956 43374 46958 43426
rect 46958 43374 47010 43426
rect 47010 43374 47012 43426
rect 46956 43372 47012 43374
rect 48412 50428 48468 50484
rect 48412 49868 48468 49924
rect 48188 49810 48244 49812
rect 48188 49758 48190 49810
rect 48190 49758 48242 49810
rect 48242 49758 48244 49810
rect 48188 49756 48244 49758
rect 48524 49644 48580 49700
rect 48412 49196 48468 49252
rect 49084 53618 49140 53620
rect 49084 53566 49086 53618
rect 49086 53566 49138 53618
rect 49138 53566 49140 53618
rect 49084 53564 49140 53566
rect 49196 53506 49252 53508
rect 49196 53454 49198 53506
rect 49198 53454 49250 53506
rect 49250 53454 49252 53506
rect 49196 53452 49252 53454
rect 49868 53452 49924 53508
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 51772 54514 51828 54516
rect 51772 54462 51774 54514
rect 51774 54462 51826 54514
rect 51826 54462 51828 54514
rect 51772 54460 51828 54462
rect 49084 52780 49140 52836
rect 50092 52834 50148 52836
rect 50092 52782 50094 52834
rect 50094 52782 50146 52834
rect 50146 52782 50148 52834
rect 50092 52780 50148 52782
rect 49084 49756 49140 49812
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 49532 49810 49588 49812
rect 49532 49758 49534 49810
rect 49534 49758 49586 49810
rect 49586 49758 49588 49810
rect 49532 49756 49588 49758
rect 51772 50316 51828 50372
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 54012 55020 54068 55076
rect 54460 55074 54516 55076
rect 54460 55022 54462 55074
rect 54462 55022 54514 55074
rect 54514 55022 54516 55074
rect 54460 55020 54516 55022
rect 52444 54626 52500 54628
rect 52444 54574 52446 54626
rect 52446 54574 52498 54626
rect 52498 54574 52500 54626
rect 52444 54572 52500 54574
rect 53228 54572 53284 54628
rect 52108 53900 52164 53956
rect 50204 49756 50260 49812
rect 49756 49698 49812 49700
rect 49756 49646 49758 49698
rect 49758 49646 49810 49698
rect 49810 49646 49812 49698
rect 49756 49644 49812 49646
rect 48636 48748 48692 48804
rect 47852 47068 47908 47124
rect 48300 47068 48356 47124
rect 50876 49308 50932 49364
rect 48860 47068 48916 47124
rect 48636 46956 48692 47012
rect 48524 46844 48580 46900
rect 49980 46898 50036 46900
rect 49980 46846 49982 46898
rect 49982 46846 50034 46898
rect 50034 46846 50036 46898
rect 49980 46844 50036 46846
rect 48748 46674 48804 46676
rect 48748 46622 48750 46674
rect 48750 46622 48802 46674
rect 48802 46622 48804 46674
rect 48748 46620 48804 46622
rect 49532 46674 49588 46676
rect 49532 46622 49534 46674
rect 49534 46622 49586 46674
rect 49586 46622 49588 46674
rect 49532 46620 49588 46622
rect 47740 45052 47796 45108
rect 45836 42476 45892 42532
rect 46732 43260 46788 43316
rect 45724 41970 45780 41972
rect 45724 41918 45726 41970
rect 45726 41918 45778 41970
rect 45778 41918 45780 41970
rect 45724 41916 45780 41918
rect 45276 41692 45332 41748
rect 45612 41692 45668 41748
rect 45500 40124 45556 40180
rect 45724 40124 45780 40180
rect 44492 35756 44548 35812
rect 45724 38668 45780 38724
rect 46396 42028 46452 42084
rect 46172 41916 46228 41972
rect 47404 42700 47460 42756
rect 47628 43372 47684 43428
rect 46732 42028 46788 42084
rect 46172 40460 46228 40516
rect 46060 40348 46116 40404
rect 48748 45106 48804 45108
rect 48748 45054 48750 45106
rect 48750 45054 48802 45106
rect 48802 45054 48804 45106
rect 48748 45052 48804 45054
rect 48524 44994 48580 44996
rect 48524 44942 48526 44994
rect 48526 44942 48578 44994
rect 48578 44942 48580 44994
rect 48524 44940 48580 44942
rect 48188 44268 48244 44324
rect 48300 44156 48356 44212
rect 48412 44044 48468 44100
rect 47852 43426 47908 43428
rect 47852 43374 47854 43426
rect 47854 43374 47906 43426
rect 47906 43374 47908 43426
rect 47852 43372 47908 43374
rect 48188 42700 48244 42756
rect 47852 41916 47908 41972
rect 47628 41804 47684 41860
rect 46956 41298 47012 41300
rect 46956 41246 46958 41298
rect 46958 41246 47010 41298
rect 47010 41246 47012 41298
rect 46956 41244 47012 41246
rect 46844 41020 46900 41076
rect 47404 41074 47460 41076
rect 47404 41022 47406 41074
rect 47406 41022 47458 41074
rect 47458 41022 47460 41074
rect 47404 41020 47460 41022
rect 48412 42476 48468 42532
rect 49868 45106 49924 45108
rect 49868 45054 49870 45106
rect 49870 45054 49922 45106
rect 49922 45054 49924 45106
rect 49868 45052 49924 45054
rect 49084 44940 49140 44996
rect 49644 44994 49700 44996
rect 49644 44942 49646 44994
rect 49646 44942 49698 44994
rect 49698 44942 49700 44994
rect 49644 44940 49700 44942
rect 51436 49532 51492 49588
rect 51100 48802 51156 48804
rect 51100 48750 51102 48802
rect 51102 48750 51154 48802
rect 51154 48750 51156 48802
rect 51100 48748 51156 48750
rect 52220 53676 52276 53732
rect 52556 53676 52612 53732
rect 53004 54514 53060 54516
rect 53004 54462 53006 54514
rect 53006 54462 53058 54514
rect 53058 54462 53060 54514
rect 53004 54460 53060 54462
rect 52668 52220 52724 52276
rect 52444 52108 52500 52164
rect 52108 49980 52164 50036
rect 51884 49586 51940 49588
rect 51884 49534 51886 49586
rect 51886 49534 51938 49586
rect 51938 49534 51940 49586
rect 51884 49532 51940 49534
rect 52556 50204 52612 50260
rect 54348 54626 54404 54628
rect 54348 54574 54350 54626
rect 54350 54574 54402 54626
rect 54402 54574 54404 54626
rect 54348 54572 54404 54574
rect 53676 54514 53732 54516
rect 53676 54462 53678 54514
rect 53678 54462 53730 54514
rect 53730 54462 53732 54514
rect 53676 54460 53732 54462
rect 54236 54514 54292 54516
rect 54236 54462 54238 54514
rect 54238 54462 54290 54514
rect 54290 54462 54292 54514
rect 54236 54460 54292 54462
rect 53452 53900 53508 53956
rect 53900 53730 53956 53732
rect 53900 53678 53902 53730
rect 53902 53678 53954 53730
rect 53954 53678 53956 53730
rect 53900 53676 53956 53678
rect 53900 52220 53956 52276
rect 53564 52162 53620 52164
rect 53564 52110 53566 52162
rect 53566 52110 53618 52162
rect 53618 52110 53620 52162
rect 53564 52108 53620 52110
rect 57148 55804 57204 55860
rect 55244 55020 55300 55076
rect 57036 55020 57092 55076
rect 53788 50540 53844 50596
rect 54236 50594 54292 50596
rect 54236 50542 54238 50594
rect 54238 50542 54290 50594
rect 54290 50542 54292 50594
rect 54236 50540 54292 50542
rect 53900 50428 53956 50484
rect 53116 50204 53172 50260
rect 53452 50316 53508 50372
rect 51660 48860 51716 48916
rect 51436 48748 51492 48804
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 52332 49308 52388 49364
rect 52332 48914 52388 48916
rect 52332 48862 52334 48914
rect 52334 48862 52386 48914
rect 52386 48862 52388 48914
rect 52332 48860 52388 48862
rect 52668 48412 52724 48468
rect 52444 48242 52500 48244
rect 52444 48190 52446 48242
rect 52446 48190 52498 48242
rect 52498 48190 52500 48242
rect 52444 48188 52500 48190
rect 50876 47404 50932 47460
rect 50204 47180 50260 47236
rect 49644 44210 49700 44212
rect 49644 44158 49646 44210
rect 49646 44158 49698 44210
rect 49698 44158 49700 44210
rect 49644 44156 49700 44158
rect 50092 44322 50148 44324
rect 50092 44270 50094 44322
rect 50094 44270 50146 44322
rect 50146 44270 50148 44322
rect 50092 44268 50148 44270
rect 49868 44044 49924 44100
rect 51100 47234 51156 47236
rect 51100 47182 51102 47234
rect 51102 47182 51154 47234
rect 51154 47182 51156 47234
rect 51100 47180 51156 47182
rect 51660 47180 51716 47236
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 50540 44994 50596 44996
rect 50540 44942 50542 44994
rect 50542 44942 50594 44994
rect 50594 44942 50596 44994
rect 50540 44940 50596 44942
rect 51100 44940 51156 44996
rect 50876 44828 50932 44884
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 49084 42530 49140 42532
rect 49084 42478 49086 42530
rect 49086 42478 49138 42530
rect 49138 42478 49140 42530
rect 49084 42476 49140 42478
rect 49532 42476 49588 42532
rect 48300 41804 48356 41860
rect 48636 41970 48692 41972
rect 48636 41918 48638 41970
rect 48638 41918 48690 41970
rect 48690 41918 48692 41970
rect 48636 41916 48692 41918
rect 49084 41244 49140 41300
rect 49196 40908 49252 40964
rect 46844 40514 46900 40516
rect 46844 40462 46846 40514
rect 46846 40462 46898 40514
rect 46898 40462 46900 40514
rect 46844 40460 46900 40462
rect 47180 40460 47236 40516
rect 46732 40236 46788 40292
rect 46732 39564 46788 39620
rect 44380 34690 44436 34692
rect 44380 34638 44382 34690
rect 44382 34638 44434 34690
rect 44434 34638 44436 34690
rect 44380 34636 44436 34638
rect 44492 34018 44548 34020
rect 44492 33966 44494 34018
rect 44494 33966 44546 34018
rect 44546 33966 44548 34018
rect 44492 33964 44548 33966
rect 44380 32956 44436 33012
rect 44268 31612 44324 31668
rect 44492 32620 44548 32676
rect 44156 29708 44212 29764
rect 42364 28588 42420 28644
rect 41356 27580 41412 27636
rect 41468 27468 41524 27524
rect 41356 27356 41412 27412
rect 41356 27186 41412 27188
rect 41356 27134 41358 27186
rect 41358 27134 41410 27186
rect 41410 27134 41412 27186
rect 41356 27132 41412 27134
rect 41692 28252 41748 28308
rect 42924 28642 42980 28644
rect 42924 28590 42926 28642
rect 42926 28590 42978 28642
rect 42978 28590 42980 28642
rect 42924 28588 42980 28590
rect 42588 28364 42644 28420
rect 42364 28028 42420 28084
rect 41804 27468 41860 27524
rect 41132 25116 41188 25172
rect 41244 26796 41300 26852
rect 41132 24162 41188 24164
rect 41132 24110 41134 24162
rect 41134 24110 41186 24162
rect 41186 24110 41188 24162
rect 41132 24108 41188 24110
rect 40908 23938 40964 23940
rect 40908 23886 40910 23938
rect 40910 23886 40962 23938
rect 40962 23886 40964 23938
rect 40908 23884 40964 23886
rect 39788 22876 39844 22932
rect 40572 23772 40628 23828
rect 40012 23378 40068 23380
rect 40012 23326 40014 23378
rect 40014 23326 40066 23378
rect 40066 23326 40068 23378
rect 40012 23324 40068 23326
rect 40124 22876 40180 22932
rect 39900 22428 39956 22484
rect 39452 20578 39508 20580
rect 39452 20526 39454 20578
rect 39454 20526 39506 20578
rect 39506 20526 39508 20578
rect 39452 20524 39508 20526
rect 39452 19404 39508 19460
rect 39340 19346 39396 19348
rect 39340 19294 39342 19346
rect 39342 19294 39394 19346
rect 39394 19294 39396 19346
rect 39340 19292 39396 19294
rect 39452 18956 39508 19012
rect 39452 16268 39508 16324
rect 40124 21756 40180 21812
rect 39788 21420 39844 21476
rect 39788 20972 39844 21028
rect 40012 20972 40068 21028
rect 40348 23100 40404 23156
rect 40796 22876 40852 22932
rect 40460 22092 40516 22148
rect 40236 20972 40292 21028
rect 40348 21308 40404 21364
rect 40124 20076 40180 20132
rect 39676 19292 39732 19348
rect 40572 21810 40628 21812
rect 40572 21758 40574 21810
rect 40574 21758 40626 21810
rect 40626 21758 40628 21810
rect 40572 21756 40628 21758
rect 40684 21308 40740 21364
rect 40684 21026 40740 21028
rect 40684 20974 40686 21026
rect 40686 20974 40738 21026
rect 40738 20974 40740 21026
rect 40684 20972 40740 20974
rect 40572 20300 40628 20356
rect 40796 20300 40852 20356
rect 40460 20076 40516 20132
rect 40348 19180 40404 19236
rect 40236 19010 40292 19012
rect 40236 18958 40238 19010
rect 40238 18958 40290 19010
rect 40290 18958 40292 19010
rect 40236 18956 40292 18958
rect 39788 18396 39844 18452
rect 40236 18450 40292 18452
rect 40236 18398 40238 18450
rect 40238 18398 40290 18450
rect 40290 18398 40292 18450
rect 40236 18396 40292 18398
rect 41020 20802 41076 20804
rect 41020 20750 41022 20802
rect 41022 20750 41074 20802
rect 41074 20750 41076 20802
rect 41020 20748 41076 20750
rect 40908 19180 40964 19236
rect 41020 19292 41076 19348
rect 40908 18844 40964 18900
rect 40460 18172 40516 18228
rect 40796 18732 40852 18788
rect 39564 17106 39620 17108
rect 39564 17054 39566 17106
rect 39566 17054 39618 17106
rect 39618 17054 39620 17106
rect 39564 17052 39620 17054
rect 39564 16156 39620 16212
rect 38332 15314 38388 15316
rect 38332 15262 38334 15314
rect 38334 15262 38386 15314
rect 38386 15262 38388 15314
rect 38332 15260 38388 15262
rect 38332 13858 38388 13860
rect 38332 13806 38334 13858
rect 38334 13806 38386 13858
rect 38386 13806 38388 13858
rect 38332 13804 38388 13806
rect 38220 13634 38276 13636
rect 38220 13582 38222 13634
rect 38222 13582 38274 13634
rect 38274 13582 38276 13634
rect 38220 13580 38276 13582
rect 37772 13356 37828 13412
rect 37324 12684 37380 12740
rect 35868 12236 35924 12292
rect 36652 12178 36708 12180
rect 36652 12126 36654 12178
rect 36654 12126 36706 12178
rect 36706 12126 36708 12178
rect 36652 12124 36708 12126
rect 36988 12290 37044 12292
rect 36988 12238 36990 12290
rect 36990 12238 37042 12290
rect 37042 12238 37044 12290
rect 36988 12236 37044 12238
rect 36876 11900 36932 11956
rect 36540 10610 36596 10612
rect 36540 10558 36542 10610
rect 36542 10558 36594 10610
rect 36594 10558 36596 10610
rect 36540 10556 36596 10558
rect 34860 9212 34916 9268
rect 35644 9324 35700 9380
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 36316 10108 36372 10164
rect 36204 9324 36260 9380
rect 37548 12124 37604 12180
rect 38892 13356 38948 13412
rect 37884 11900 37940 11956
rect 38556 12684 38612 12740
rect 38332 11900 38388 11956
rect 37100 10108 37156 10164
rect 38108 9996 38164 10052
rect 35980 8428 36036 8484
rect 34972 8316 35028 8372
rect 35308 8316 35364 8372
rect 35532 8258 35588 8260
rect 35532 8206 35534 8258
rect 35534 8206 35586 8258
rect 35586 8206 35588 8258
rect 35532 8204 35588 8206
rect 35980 8258 36036 8260
rect 35980 8206 35982 8258
rect 35982 8206 36034 8258
rect 36034 8206 36036 8258
rect 35980 8204 36036 8206
rect 37436 9884 37492 9940
rect 37884 9884 37940 9940
rect 37996 9826 38052 9828
rect 37996 9774 37998 9826
rect 37998 9774 38050 9826
rect 38050 9774 38052 9826
rect 37996 9772 38052 9774
rect 37548 9714 37604 9716
rect 37548 9662 37550 9714
rect 37550 9662 37602 9714
rect 37602 9662 37604 9714
rect 37548 9660 37604 9662
rect 36316 8092 36372 8148
rect 37324 8428 37380 8484
rect 37884 9042 37940 9044
rect 37884 8990 37886 9042
rect 37886 8990 37938 9042
rect 37938 8990 37940 9042
rect 37884 8988 37940 8990
rect 38108 8428 38164 8484
rect 34860 6690 34916 6692
rect 34860 6638 34862 6690
rect 34862 6638 34914 6690
rect 34914 6638 34916 6690
rect 34860 6636 34916 6638
rect 34748 5852 34804 5908
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35084 6636 35140 6692
rect 35980 6690 36036 6692
rect 35980 6638 35982 6690
rect 35982 6638 36034 6690
rect 36034 6638 36036 6690
rect 35980 6636 36036 6638
rect 35532 6018 35588 6020
rect 35532 5966 35534 6018
rect 35534 5966 35586 6018
rect 35586 5966 35588 6018
rect 35532 5964 35588 5966
rect 35308 5906 35364 5908
rect 35308 5854 35310 5906
rect 35310 5854 35362 5906
rect 35362 5854 35364 5906
rect 35308 5852 35364 5854
rect 36988 5964 37044 6020
rect 37660 5852 37716 5908
rect 35644 5794 35700 5796
rect 35644 5742 35646 5794
rect 35646 5742 35698 5794
rect 35698 5742 35700 5794
rect 35644 5740 35700 5742
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 33964 4956 34020 5012
rect 34412 4732 34468 4788
rect 33516 3388 33572 3444
rect 34076 4396 34132 4452
rect 33852 3612 33908 3668
rect 36652 5180 36708 5236
rect 35644 5122 35700 5124
rect 35644 5070 35646 5122
rect 35646 5070 35698 5122
rect 35698 5070 35700 5122
rect 35644 5068 35700 5070
rect 36428 5122 36484 5124
rect 36428 5070 36430 5122
rect 36430 5070 36482 5122
rect 36482 5070 36484 5122
rect 36428 5068 36484 5070
rect 34972 4956 35028 5012
rect 35308 4956 35364 5012
rect 34412 3724 34468 3780
rect 36540 4284 36596 4340
rect 37212 4338 37268 4340
rect 37212 4286 37214 4338
rect 37214 4286 37266 4338
rect 37266 4286 37268 4338
rect 37212 4284 37268 4286
rect 35420 4226 35476 4228
rect 35420 4174 35422 4226
rect 35422 4174 35474 4226
rect 35474 4174 35476 4226
rect 35420 4172 35476 4174
rect 35308 4060 35364 4116
rect 35532 4060 35588 4116
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 34524 3666 34580 3668
rect 34524 3614 34526 3666
rect 34526 3614 34578 3666
rect 34578 3614 34580 3666
rect 34524 3612 34580 3614
rect 36988 4226 37044 4228
rect 36988 4174 36990 4226
rect 36990 4174 37042 4226
rect 37042 4174 37044 4226
rect 36988 4172 37044 4174
rect 36204 4060 36260 4116
rect 35756 3666 35812 3668
rect 35756 3614 35758 3666
rect 35758 3614 35810 3666
rect 35810 3614 35812 3666
rect 35756 3612 35812 3614
rect 39228 15426 39284 15428
rect 39228 15374 39230 15426
rect 39230 15374 39282 15426
rect 39282 15374 39284 15426
rect 39228 15372 39284 15374
rect 39340 15260 39396 15316
rect 39900 15314 39956 15316
rect 39900 15262 39902 15314
rect 39902 15262 39954 15314
rect 39954 15262 39956 15314
rect 39900 15260 39956 15262
rect 39564 13804 39620 13860
rect 39788 13970 39844 13972
rect 39788 13918 39790 13970
rect 39790 13918 39842 13970
rect 39842 13918 39844 13970
rect 39788 13916 39844 13918
rect 40348 17442 40404 17444
rect 40348 17390 40350 17442
rect 40350 17390 40402 17442
rect 40402 17390 40404 17442
rect 40348 17388 40404 17390
rect 40348 17164 40404 17220
rect 40124 16044 40180 16100
rect 40236 16380 40292 16436
rect 40236 15372 40292 15428
rect 40572 17106 40628 17108
rect 40572 17054 40574 17106
rect 40574 17054 40626 17106
rect 40626 17054 40628 17106
rect 40572 17052 40628 17054
rect 40684 16658 40740 16660
rect 40684 16606 40686 16658
rect 40686 16606 40738 16658
rect 40738 16606 40740 16658
rect 40684 16604 40740 16606
rect 40908 17388 40964 17444
rect 40460 14924 40516 14980
rect 40012 14028 40068 14084
rect 39676 13020 39732 13076
rect 40124 13916 40180 13972
rect 39788 12908 39844 12964
rect 39452 12738 39508 12740
rect 39452 12686 39454 12738
rect 39454 12686 39506 12738
rect 39506 12686 39508 12738
rect 39452 12684 39508 12686
rect 38780 11676 38836 11732
rect 39452 12290 39508 12292
rect 39452 12238 39454 12290
rect 39454 12238 39506 12290
rect 39506 12238 39508 12290
rect 39452 12236 39508 12238
rect 39228 11900 39284 11956
rect 39340 11676 39396 11732
rect 40012 11676 40068 11732
rect 40236 12236 40292 12292
rect 40796 15260 40852 15316
rect 41916 27020 41972 27076
rect 42252 26962 42308 26964
rect 42252 26910 42254 26962
rect 42254 26910 42306 26962
rect 42306 26910 42308 26962
rect 42252 26908 42308 26910
rect 44044 29314 44100 29316
rect 44044 29262 44046 29314
rect 44046 29262 44098 29314
rect 44098 29262 44100 29314
rect 44044 29260 44100 29262
rect 43036 28252 43092 28308
rect 43148 29202 43204 29204
rect 43148 29150 43150 29202
rect 43150 29150 43202 29202
rect 43202 29150 43204 29202
rect 43148 29148 43204 29150
rect 43372 29148 43428 29204
rect 42700 27186 42756 27188
rect 42700 27134 42702 27186
rect 42702 27134 42754 27186
rect 42754 27134 42756 27186
rect 42700 27132 42756 27134
rect 42924 27580 42980 27636
rect 41916 26290 41972 26292
rect 41916 26238 41918 26290
rect 41918 26238 41970 26290
rect 41970 26238 41972 26290
rect 41916 26236 41972 26238
rect 41692 26012 41748 26068
rect 41468 25618 41524 25620
rect 41468 25566 41470 25618
rect 41470 25566 41522 25618
rect 41522 25566 41524 25618
rect 41468 25564 41524 25566
rect 42140 25228 42196 25284
rect 42364 26178 42420 26180
rect 42364 26126 42366 26178
rect 42366 26126 42418 26178
rect 42418 26126 42420 26178
rect 42364 26124 42420 26126
rect 42364 25618 42420 25620
rect 42364 25566 42366 25618
rect 42366 25566 42418 25618
rect 42418 25566 42420 25618
rect 42364 25564 42420 25566
rect 42812 25506 42868 25508
rect 42812 25454 42814 25506
rect 42814 25454 42866 25506
rect 42866 25454 42868 25506
rect 42812 25452 42868 25454
rect 42252 25004 42308 25060
rect 42364 25228 42420 25284
rect 41692 24108 41748 24164
rect 41468 23826 41524 23828
rect 41468 23774 41470 23826
rect 41470 23774 41522 23826
rect 41522 23774 41524 23826
rect 41468 23772 41524 23774
rect 42028 23884 42084 23940
rect 41692 22876 41748 22932
rect 41468 22146 41524 22148
rect 41468 22094 41470 22146
rect 41470 22094 41522 22146
rect 41522 22094 41524 22146
rect 41468 22092 41524 22094
rect 41468 21586 41524 21588
rect 41468 21534 41470 21586
rect 41470 21534 41522 21586
rect 41522 21534 41524 21586
rect 41468 21532 41524 21534
rect 41244 19292 41300 19348
rect 41468 19234 41524 19236
rect 41468 19182 41470 19234
rect 41470 19182 41522 19234
rect 41522 19182 41524 19234
rect 41468 19180 41524 19182
rect 41356 18620 41412 18676
rect 41356 17778 41412 17780
rect 41356 17726 41358 17778
rect 41358 17726 41410 17778
rect 41410 17726 41412 17778
rect 41356 17724 41412 17726
rect 41916 21196 41972 21252
rect 42028 21308 42084 21364
rect 43148 26962 43204 26964
rect 43148 26910 43150 26962
rect 43150 26910 43202 26962
rect 43202 26910 43204 26962
rect 43148 26908 43204 26910
rect 43036 26124 43092 26180
rect 43148 25900 43204 25956
rect 42476 23826 42532 23828
rect 42476 23774 42478 23826
rect 42478 23774 42530 23826
rect 42530 23774 42532 23826
rect 42476 23772 42532 23774
rect 42588 23154 42644 23156
rect 42588 23102 42590 23154
rect 42590 23102 42642 23154
rect 42642 23102 42644 23154
rect 42588 23100 42644 23102
rect 42924 23938 42980 23940
rect 42924 23886 42926 23938
rect 42926 23886 42978 23938
rect 42978 23886 42980 23938
rect 42924 23884 42980 23886
rect 43260 25228 43316 25284
rect 42364 22146 42420 22148
rect 42364 22094 42366 22146
rect 42366 22094 42418 22146
rect 42418 22094 42420 22146
rect 42364 22092 42420 22094
rect 43932 28924 43988 28980
rect 43708 28530 43764 28532
rect 43708 28478 43710 28530
rect 43710 28478 43762 28530
rect 43762 28478 43764 28530
rect 43708 28476 43764 28478
rect 43596 28028 43652 28084
rect 44044 28364 44100 28420
rect 43596 27580 43652 27636
rect 44044 26962 44100 26964
rect 44044 26910 44046 26962
rect 44046 26910 44098 26962
rect 44098 26910 44100 26962
rect 44044 26908 44100 26910
rect 45724 37826 45780 37828
rect 45724 37774 45726 37826
rect 45726 37774 45778 37826
rect 45778 37774 45780 37826
rect 45724 37772 45780 37774
rect 45052 37378 45108 37380
rect 45052 37326 45054 37378
rect 45054 37326 45106 37378
rect 45106 37326 45108 37378
rect 45052 37324 45108 37326
rect 45052 36540 45108 36596
rect 44940 35810 44996 35812
rect 44940 35758 44942 35810
rect 44942 35758 44994 35810
rect 44994 35758 44996 35810
rect 44940 35756 44996 35758
rect 44940 34636 44996 34692
rect 44828 32956 44884 33012
rect 44940 32396 44996 32452
rect 44828 31948 44884 32004
rect 44716 31666 44772 31668
rect 44716 31614 44718 31666
rect 44718 31614 44770 31666
rect 44770 31614 44772 31666
rect 44716 31612 44772 31614
rect 44268 26908 44324 26964
rect 43708 26514 43764 26516
rect 43708 26462 43710 26514
rect 43710 26462 43762 26514
rect 43762 26462 43764 26514
rect 43708 26460 43764 26462
rect 43596 26402 43652 26404
rect 43596 26350 43598 26402
rect 43598 26350 43650 26402
rect 43650 26350 43652 26402
rect 43596 26348 43652 26350
rect 43484 23154 43540 23156
rect 43484 23102 43486 23154
rect 43486 23102 43538 23154
rect 43538 23102 43540 23154
rect 43484 23100 43540 23102
rect 42812 21756 42868 21812
rect 42588 21196 42644 21252
rect 42364 20802 42420 20804
rect 42364 20750 42366 20802
rect 42366 20750 42418 20802
rect 42418 20750 42420 20802
rect 42364 20748 42420 20750
rect 43484 21308 43540 21364
rect 43148 21196 43204 21252
rect 43820 26012 43876 26068
rect 44268 25900 44324 25956
rect 44716 28588 44772 28644
rect 44604 28140 44660 28196
rect 44492 27132 44548 27188
rect 43932 25506 43988 25508
rect 43932 25454 43934 25506
rect 43934 25454 43986 25506
rect 43986 25454 43988 25506
rect 43932 25452 43988 25454
rect 44044 25282 44100 25284
rect 44044 25230 44046 25282
rect 44046 25230 44098 25282
rect 44098 25230 44100 25282
rect 44044 25228 44100 25230
rect 43932 23996 43988 24052
rect 43820 23436 43876 23492
rect 44156 21756 44212 21812
rect 43932 21474 43988 21476
rect 43932 21422 43934 21474
rect 43934 21422 43986 21474
rect 43986 21422 43988 21474
rect 43932 21420 43988 21422
rect 43708 21084 43764 21140
rect 43036 20748 43092 20804
rect 41580 18844 41636 18900
rect 41580 18620 41636 18676
rect 42252 18620 42308 18676
rect 42588 19964 42644 20020
rect 42924 19180 42980 19236
rect 42812 19068 42868 19124
rect 44044 19234 44100 19236
rect 44044 19182 44046 19234
rect 44046 19182 44098 19234
rect 44098 19182 44100 19234
rect 44044 19180 44100 19182
rect 44156 19122 44212 19124
rect 44156 19070 44158 19122
rect 44158 19070 44210 19122
rect 44210 19070 44212 19122
rect 44156 19068 44212 19070
rect 44940 25340 44996 25396
rect 44380 25228 44436 25284
rect 44604 25282 44660 25284
rect 44604 25230 44606 25282
rect 44606 25230 44658 25282
rect 44658 25230 44660 25282
rect 44604 25228 44660 25230
rect 45500 35922 45556 35924
rect 45500 35870 45502 35922
rect 45502 35870 45554 35922
rect 45554 35870 45556 35922
rect 45500 35868 45556 35870
rect 45388 35810 45444 35812
rect 45388 35758 45390 35810
rect 45390 35758 45442 35810
rect 45442 35758 45444 35810
rect 45388 35756 45444 35758
rect 46508 39394 46564 39396
rect 46508 39342 46510 39394
rect 46510 39342 46562 39394
rect 46562 39342 46564 39394
rect 46508 39340 46564 39342
rect 45948 35756 46004 35812
rect 46060 38668 46116 38724
rect 45948 35532 46004 35588
rect 45724 35420 45780 35476
rect 45500 33852 45556 33908
rect 45164 32284 45220 32340
rect 45500 32450 45556 32452
rect 45500 32398 45502 32450
rect 45502 32398 45554 32450
rect 45554 32398 45556 32450
rect 45500 32396 45556 32398
rect 45836 34412 45892 34468
rect 46956 40348 47012 40404
rect 46284 38722 46340 38724
rect 46284 38670 46286 38722
rect 46286 38670 46338 38722
rect 46338 38670 46340 38722
rect 46284 38668 46340 38670
rect 46732 38780 46788 38836
rect 46172 38556 46228 38612
rect 46284 37772 46340 37828
rect 46284 36988 46340 37044
rect 46844 37324 46900 37380
rect 46732 36988 46788 37044
rect 46508 35868 46564 35924
rect 46620 36092 46676 36148
rect 46172 35586 46228 35588
rect 46172 35534 46174 35586
rect 46174 35534 46226 35586
rect 46226 35534 46228 35586
rect 46172 35532 46228 35534
rect 45388 30604 45444 30660
rect 45164 29708 45220 29764
rect 45388 28754 45444 28756
rect 45388 28702 45390 28754
rect 45390 28702 45442 28754
rect 45442 28702 45444 28754
rect 45388 28700 45444 28702
rect 46060 33852 46116 33908
rect 46060 33068 46116 33124
rect 45612 30044 45668 30100
rect 46060 31778 46116 31780
rect 46060 31726 46062 31778
rect 46062 31726 46114 31778
rect 46114 31726 46116 31778
rect 46060 31724 46116 31726
rect 45836 31666 45892 31668
rect 45836 31614 45838 31666
rect 45838 31614 45890 31666
rect 45890 31614 45892 31666
rect 45836 31612 45892 31614
rect 45948 31554 46004 31556
rect 45948 31502 45950 31554
rect 45950 31502 46002 31554
rect 46002 31502 46004 31554
rect 45948 31500 46004 31502
rect 46060 29986 46116 29988
rect 46060 29934 46062 29986
rect 46062 29934 46114 29986
rect 46114 29934 46116 29986
rect 46060 29932 46116 29934
rect 45724 29314 45780 29316
rect 45724 29262 45726 29314
rect 45726 29262 45778 29314
rect 45778 29262 45780 29314
rect 45724 29260 45780 29262
rect 45612 27970 45668 27972
rect 45612 27918 45614 27970
rect 45614 27918 45666 27970
rect 45666 27918 45668 27970
rect 45612 27916 45668 27918
rect 45500 27804 45556 27860
rect 45612 27298 45668 27300
rect 45612 27246 45614 27298
rect 45614 27246 45666 27298
rect 45666 27246 45668 27298
rect 45612 27244 45668 27246
rect 46508 33122 46564 33124
rect 46508 33070 46510 33122
rect 46510 33070 46562 33122
rect 46562 33070 46564 33122
rect 46508 33068 46564 33070
rect 46396 30770 46452 30772
rect 46396 30718 46398 30770
rect 46398 30718 46450 30770
rect 46450 30718 46452 30770
rect 46396 30716 46452 30718
rect 47068 39340 47124 39396
rect 47852 40348 47908 40404
rect 47292 39618 47348 39620
rect 47292 39566 47294 39618
rect 47294 39566 47346 39618
rect 47346 39566 47348 39618
rect 47292 39564 47348 39566
rect 47404 36988 47460 37044
rect 47180 35980 47236 36036
rect 46620 30604 46676 30660
rect 46956 34242 47012 34244
rect 46956 34190 46958 34242
rect 46958 34190 47010 34242
rect 47010 34190 47012 34242
rect 46956 34188 47012 34190
rect 47068 33122 47124 33124
rect 47068 33070 47070 33122
rect 47070 33070 47122 33122
rect 47122 33070 47124 33122
rect 47068 33068 47124 33070
rect 47292 35868 47348 35924
rect 47516 35196 47572 35252
rect 47964 39452 48020 39508
rect 48524 40514 48580 40516
rect 48524 40462 48526 40514
rect 48526 40462 48578 40514
rect 48578 40462 48580 40514
rect 48524 40460 48580 40462
rect 48636 39394 48692 39396
rect 48636 39342 48638 39394
rect 48638 39342 48690 39394
rect 48690 39342 48692 39394
rect 48636 39340 48692 39342
rect 48076 38834 48132 38836
rect 48076 38782 48078 38834
rect 48078 38782 48130 38834
rect 48130 38782 48132 38834
rect 48076 38780 48132 38782
rect 48748 38722 48804 38724
rect 48748 38670 48750 38722
rect 48750 38670 48802 38722
rect 48802 38670 48804 38722
rect 48748 38668 48804 38670
rect 47852 36988 47908 37044
rect 47740 35586 47796 35588
rect 47740 35534 47742 35586
rect 47742 35534 47794 35586
rect 47794 35534 47796 35586
rect 47740 35532 47796 35534
rect 47628 34972 47684 35028
rect 47740 35308 47796 35364
rect 47404 34188 47460 34244
rect 47628 34018 47684 34020
rect 47628 33966 47630 34018
rect 47630 33966 47682 34018
rect 47682 33966 47684 34018
rect 47628 33964 47684 33966
rect 47180 31724 47236 31780
rect 47404 31052 47460 31108
rect 46284 29820 46340 29876
rect 46396 29708 46452 29764
rect 46284 29650 46340 29652
rect 46284 29598 46286 29650
rect 46286 29598 46338 29650
rect 46338 29598 46340 29650
rect 46284 29596 46340 29598
rect 46060 29148 46116 29204
rect 46172 29314 46228 29316
rect 46172 29262 46174 29314
rect 46174 29262 46226 29314
rect 46226 29262 46228 29314
rect 46172 29260 46228 29262
rect 45836 28140 45892 28196
rect 45948 28700 46004 28756
rect 46284 28754 46340 28756
rect 46284 28702 46286 28754
rect 46286 28702 46338 28754
rect 46338 28702 46340 28754
rect 46284 28700 46340 28702
rect 45948 27858 46004 27860
rect 45948 27806 45950 27858
rect 45950 27806 46002 27858
rect 46002 27806 46004 27858
rect 45948 27804 46004 27806
rect 46620 28588 46676 28644
rect 45388 26572 45444 26628
rect 44380 24050 44436 24052
rect 44380 23998 44382 24050
rect 44382 23998 44434 24050
rect 44434 23998 44436 24050
rect 44380 23996 44436 23998
rect 45500 26348 45556 26404
rect 45612 26290 45668 26292
rect 45612 26238 45614 26290
rect 45614 26238 45666 26290
rect 45666 26238 45668 26290
rect 45612 26236 45668 26238
rect 46060 27356 46116 27412
rect 46508 28140 46564 28196
rect 46172 27186 46228 27188
rect 46172 27134 46174 27186
rect 46174 27134 46226 27186
rect 46226 27134 46228 27186
rect 46172 27132 46228 27134
rect 46508 26908 46564 26964
rect 45948 26796 46004 26852
rect 46060 26402 46116 26404
rect 46060 26350 46062 26402
rect 46062 26350 46114 26402
rect 46114 26350 46116 26402
rect 46060 26348 46116 26350
rect 45948 26236 46004 26292
rect 45500 25394 45556 25396
rect 45500 25342 45502 25394
rect 45502 25342 45554 25394
rect 45554 25342 45556 25394
rect 45500 25340 45556 25342
rect 45388 24722 45444 24724
rect 45388 24670 45390 24722
rect 45390 24670 45442 24722
rect 45442 24670 45444 24722
rect 45388 24668 45444 24670
rect 44940 23212 44996 23268
rect 45052 23996 45108 24052
rect 45612 25282 45668 25284
rect 45612 25230 45614 25282
rect 45614 25230 45666 25282
rect 45666 25230 45668 25282
rect 45612 25228 45668 25230
rect 45836 23938 45892 23940
rect 45836 23886 45838 23938
rect 45838 23886 45890 23938
rect 45890 23886 45892 23938
rect 45836 23884 45892 23886
rect 46060 24498 46116 24500
rect 46060 24446 46062 24498
rect 46062 24446 46114 24498
rect 46114 24446 46116 24498
rect 46060 24444 46116 24446
rect 45724 23436 45780 23492
rect 45388 22876 45444 22932
rect 45612 22988 45668 23044
rect 44828 22370 44884 22372
rect 44828 22318 44830 22370
rect 44830 22318 44882 22370
rect 44882 22318 44884 22370
rect 44828 22316 44884 22318
rect 45500 22370 45556 22372
rect 45500 22318 45502 22370
rect 45502 22318 45554 22370
rect 45554 22318 45556 22370
rect 45500 22316 45556 22318
rect 45052 21698 45108 21700
rect 45052 21646 45054 21698
rect 45054 21646 45106 21698
rect 45106 21646 45108 21698
rect 45052 21644 45108 21646
rect 44716 21474 44772 21476
rect 44716 21422 44718 21474
rect 44718 21422 44770 21474
rect 44770 21422 44772 21474
rect 44716 21420 44772 21422
rect 44492 21308 44548 21364
rect 45724 22204 45780 22260
rect 46060 22370 46116 22372
rect 46060 22318 46062 22370
rect 46062 22318 46114 22370
rect 46114 22318 46116 22370
rect 46060 22316 46116 22318
rect 46620 26572 46676 26628
rect 46732 27916 46788 27972
rect 46732 26236 46788 26292
rect 47852 34188 47908 34244
rect 47740 31164 47796 31220
rect 47516 30156 47572 30212
rect 47292 29986 47348 29988
rect 47292 29934 47294 29986
rect 47294 29934 47346 29986
rect 47346 29934 47348 29986
rect 47292 29932 47348 29934
rect 46956 29820 47012 29876
rect 47068 28754 47124 28756
rect 47068 28702 47070 28754
rect 47070 28702 47122 28754
rect 47122 28702 47124 28754
rect 47068 28700 47124 28702
rect 47516 29596 47572 29652
rect 47740 29932 47796 29988
rect 47180 28642 47236 28644
rect 47180 28590 47182 28642
rect 47182 28590 47234 28642
rect 47234 28590 47236 28642
rect 47180 28588 47236 28590
rect 47404 27970 47460 27972
rect 47404 27918 47406 27970
rect 47406 27918 47458 27970
rect 47458 27918 47460 27970
rect 47404 27916 47460 27918
rect 48300 35644 48356 35700
rect 49084 35084 49140 35140
rect 48188 34972 48244 35028
rect 48972 34972 49028 35028
rect 48972 34076 49028 34132
rect 48188 31164 48244 31220
rect 48524 31836 48580 31892
rect 48412 31778 48468 31780
rect 48412 31726 48414 31778
rect 48414 31726 48466 31778
rect 48466 31726 48468 31778
rect 48412 31724 48468 31726
rect 48412 31164 48468 31220
rect 48188 30604 48244 30660
rect 48412 30322 48468 30324
rect 48412 30270 48414 30322
rect 48414 30270 48466 30322
rect 48466 30270 48468 30322
rect 48412 30268 48468 30270
rect 48524 30156 48580 30212
rect 48300 29986 48356 29988
rect 48300 29934 48302 29986
rect 48302 29934 48354 29986
rect 48354 29934 48356 29986
rect 48300 29932 48356 29934
rect 48076 29596 48132 29652
rect 49196 32732 49252 32788
rect 49420 41186 49476 41188
rect 49420 41134 49422 41186
rect 49422 41134 49474 41186
rect 49474 41134 49476 41186
rect 49420 41132 49476 41134
rect 49308 39340 49364 39396
rect 49084 31666 49140 31668
rect 49084 31614 49086 31666
rect 49086 31614 49138 31666
rect 49138 31614 49140 31666
rect 49084 31612 49140 31614
rect 49756 41804 49812 41860
rect 49980 41356 50036 41412
rect 50204 40962 50260 40964
rect 50204 40910 50206 40962
rect 50206 40910 50258 40962
rect 50258 40910 50260 40962
rect 50204 40908 50260 40910
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 50764 40962 50820 40964
rect 50764 40910 50766 40962
rect 50766 40910 50818 40962
rect 50818 40910 50820 40962
rect 50764 40908 50820 40910
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 50764 40514 50820 40516
rect 50764 40462 50766 40514
rect 50766 40462 50818 40514
rect 50818 40462 50820 40514
rect 50764 40460 50820 40462
rect 49868 39340 49924 39396
rect 49868 38892 49924 38948
rect 50092 38780 50148 38836
rect 49980 38668 50036 38724
rect 51548 44940 51604 44996
rect 51884 47458 51940 47460
rect 51884 47406 51886 47458
rect 51886 47406 51938 47458
rect 51938 47406 51940 47458
rect 51884 47404 51940 47406
rect 53116 50034 53172 50036
rect 53116 49982 53118 50034
rect 53118 49982 53170 50034
rect 53170 49982 53172 50034
rect 53116 49980 53172 49982
rect 53340 48914 53396 48916
rect 53340 48862 53342 48914
rect 53342 48862 53394 48914
rect 53394 48862 53396 48914
rect 53340 48860 53396 48862
rect 53676 50204 53732 50260
rect 53564 49308 53620 49364
rect 53788 49698 53844 49700
rect 53788 49646 53790 49698
rect 53790 49646 53842 49698
rect 53842 49646 53844 49698
rect 53788 49644 53844 49646
rect 53116 48466 53172 48468
rect 53116 48414 53118 48466
rect 53118 48414 53170 48466
rect 53170 48414 53172 48466
rect 53116 48412 53172 48414
rect 52892 45836 52948 45892
rect 51884 45164 51940 45220
rect 53452 46450 53508 46452
rect 53452 46398 53454 46450
rect 53454 46398 53506 46450
rect 53506 46398 53508 46450
rect 53452 46396 53508 46398
rect 53228 45836 53284 45892
rect 51996 44828 52052 44884
rect 52108 45052 52164 45108
rect 53340 45106 53396 45108
rect 53340 45054 53342 45106
rect 53342 45054 53394 45106
rect 53394 45054 53396 45106
rect 53340 45052 53396 45054
rect 51772 42812 51828 42868
rect 52108 44156 52164 44212
rect 51100 41970 51156 41972
rect 51100 41918 51102 41970
rect 51102 41918 51154 41970
rect 51154 41918 51156 41970
rect 51100 41916 51156 41918
rect 51212 41132 51268 41188
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 50876 38892 50932 38948
rect 50540 38834 50596 38836
rect 50540 38782 50542 38834
rect 50542 38782 50594 38834
rect 50594 38782 50596 38834
rect 50540 38780 50596 38782
rect 50764 38162 50820 38164
rect 50764 38110 50766 38162
rect 50766 38110 50818 38162
rect 50818 38110 50820 38162
rect 50764 38108 50820 38110
rect 50428 38050 50484 38052
rect 50428 37998 50430 38050
rect 50430 37998 50482 38050
rect 50482 37998 50484 38050
rect 50428 37996 50484 37998
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 50204 36540 50260 36596
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 51660 40908 51716 40964
rect 51324 38834 51380 38836
rect 51324 38782 51326 38834
rect 51326 38782 51378 38834
rect 51378 38782 51380 38834
rect 51324 38780 51380 38782
rect 51436 38722 51492 38724
rect 51436 38670 51438 38722
rect 51438 38670 51490 38722
rect 51490 38670 51492 38722
rect 51436 38668 51492 38670
rect 53788 45890 53844 45892
rect 53788 45838 53790 45890
rect 53790 45838 53842 45890
rect 53842 45838 53844 45890
rect 53788 45836 53844 45838
rect 53788 44828 53844 44884
rect 54124 50482 54180 50484
rect 54124 50430 54126 50482
rect 54126 50430 54178 50482
rect 54178 50430 54180 50482
rect 54124 50428 54180 50430
rect 54460 49644 54516 49700
rect 54124 49308 54180 49364
rect 55356 49308 55412 49364
rect 55916 49698 55972 49700
rect 55916 49646 55918 49698
rect 55918 49646 55970 49698
rect 55970 49646 55972 49698
rect 55916 49644 55972 49646
rect 55580 49196 55636 49252
rect 54796 48242 54852 48244
rect 54796 48190 54798 48242
rect 54798 48190 54850 48242
rect 54850 48190 54852 48242
rect 54796 48188 54852 48190
rect 54460 47740 54516 47796
rect 54012 46396 54068 46452
rect 54572 47458 54628 47460
rect 54572 47406 54574 47458
rect 54574 47406 54626 47458
rect 54626 47406 54628 47458
rect 54572 47404 54628 47406
rect 55468 48802 55524 48804
rect 55468 48750 55470 48802
rect 55470 48750 55522 48802
rect 55522 48750 55524 48802
rect 55468 48748 55524 48750
rect 55356 47404 55412 47460
rect 55244 47292 55300 47348
rect 55468 46732 55524 46788
rect 55244 46674 55300 46676
rect 55244 46622 55246 46674
rect 55246 46622 55298 46674
rect 55298 46622 55300 46674
rect 55244 46620 55300 46622
rect 55692 47516 55748 47572
rect 55692 47292 55748 47348
rect 56252 50540 56308 50596
rect 56812 50594 56868 50596
rect 56812 50542 56814 50594
rect 56814 50542 56866 50594
rect 56866 50542 56868 50594
rect 56812 50540 56868 50542
rect 56364 49756 56420 49812
rect 56700 49698 56756 49700
rect 56700 49646 56702 49698
rect 56702 49646 56754 49698
rect 56754 49646 56756 49698
rect 56700 49644 56756 49646
rect 56700 49026 56756 49028
rect 56700 48974 56702 49026
rect 56702 48974 56754 49026
rect 56754 48974 56756 49026
rect 56700 48972 56756 48974
rect 56812 48188 56868 48244
rect 56364 47570 56420 47572
rect 56364 47518 56366 47570
rect 56366 47518 56418 47570
rect 56418 47518 56420 47570
rect 56364 47516 56420 47518
rect 56252 47346 56308 47348
rect 56252 47294 56254 47346
rect 56254 47294 56306 47346
rect 56306 47294 56308 47346
rect 56252 47292 56308 47294
rect 55580 46396 55636 46452
rect 56028 46450 56084 46452
rect 56028 46398 56030 46450
rect 56030 46398 56082 46450
rect 56082 46398 56084 46450
rect 56028 46396 56084 46398
rect 55804 46172 55860 46228
rect 54236 45612 54292 45668
rect 54012 45218 54068 45220
rect 54012 45166 54014 45218
rect 54014 45166 54066 45218
rect 54066 45166 54068 45218
rect 54012 45164 54068 45166
rect 53900 44156 53956 44212
rect 53900 42866 53956 42868
rect 53900 42814 53902 42866
rect 53902 42814 53954 42866
rect 53954 42814 53956 42866
rect 53900 42812 53956 42814
rect 53564 42028 53620 42084
rect 52220 41916 52276 41972
rect 52668 41970 52724 41972
rect 52668 41918 52670 41970
rect 52670 41918 52722 41970
rect 52722 41918 52724 41970
rect 52668 41916 52724 41918
rect 53452 41916 53508 41972
rect 52108 41132 52164 41188
rect 52444 41580 52500 41636
rect 51884 40962 51940 40964
rect 51884 40910 51886 40962
rect 51886 40910 51938 40962
rect 51938 40910 51940 40962
rect 51884 40908 51940 40910
rect 53228 41746 53284 41748
rect 53228 41694 53230 41746
rect 53230 41694 53282 41746
rect 53282 41694 53284 41746
rect 53228 41692 53284 41694
rect 53004 41244 53060 41300
rect 53452 41468 53508 41524
rect 53340 41132 53396 41188
rect 52444 40908 52500 40964
rect 52668 40962 52724 40964
rect 52668 40910 52670 40962
rect 52670 40910 52722 40962
rect 52722 40910 52724 40962
rect 52668 40908 52724 40910
rect 53228 40348 53284 40404
rect 52220 38946 52276 38948
rect 52220 38894 52222 38946
rect 52222 38894 52274 38946
rect 52274 38894 52276 38946
rect 52220 38892 52276 38894
rect 51884 38108 51940 38164
rect 51772 37996 51828 38052
rect 50428 35868 50484 35924
rect 51100 35868 51156 35924
rect 49420 35532 49476 35588
rect 49980 35532 50036 35588
rect 49532 35084 49588 35140
rect 51212 34860 51268 34916
rect 49420 34076 49476 34132
rect 50876 34748 50932 34804
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 49980 34130 50036 34132
rect 49980 34078 49982 34130
rect 49982 34078 50034 34130
rect 50034 34078 50036 34130
rect 49980 34076 50036 34078
rect 49084 30156 49140 30212
rect 47964 27916 48020 27972
rect 47740 27804 47796 27860
rect 47404 27356 47460 27412
rect 46956 27244 47012 27300
rect 46620 25340 46676 25396
rect 46844 24444 46900 24500
rect 47516 26908 47572 26964
rect 48412 27298 48468 27300
rect 48412 27246 48414 27298
rect 48414 27246 48466 27298
rect 48466 27246 48468 27298
rect 48412 27244 48468 27246
rect 48188 26908 48244 26964
rect 47180 25340 47236 25396
rect 46508 23826 46564 23828
rect 46508 23774 46510 23826
rect 46510 23774 46562 23826
rect 46562 23774 46564 23826
rect 46508 23772 46564 23774
rect 46284 23436 46340 23492
rect 46396 23548 46452 23604
rect 46956 23548 47012 23604
rect 46732 22988 46788 23044
rect 47628 26796 47684 26852
rect 48636 27970 48692 27972
rect 48636 27918 48638 27970
rect 48638 27918 48690 27970
rect 48690 27918 48692 27970
rect 48636 27916 48692 27918
rect 48972 27804 49028 27860
rect 48412 26850 48468 26852
rect 48412 26798 48414 26850
rect 48414 26798 48466 26850
rect 48466 26798 48468 26850
rect 48412 26796 48468 26798
rect 48300 26460 48356 26516
rect 48300 26290 48356 26292
rect 48300 26238 48302 26290
rect 48302 26238 48354 26290
rect 48354 26238 48356 26290
rect 48300 26236 48356 26238
rect 47740 25340 47796 25396
rect 47852 24892 47908 24948
rect 48412 25340 48468 25396
rect 48860 26460 48916 26516
rect 49196 30098 49252 30100
rect 49196 30046 49198 30098
rect 49198 30046 49250 30098
rect 49250 30046 49252 30098
rect 49196 30044 49252 30046
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 49868 32786 49924 32788
rect 49868 32734 49870 32786
rect 49870 32734 49922 32786
rect 49922 32734 49924 32786
rect 49868 32732 49924 32734
rect 53340 37884 53396 37940
rect 54908 45666 54964 45668
rect 54908 45614 54910 45666
rect 54910 45614 54962 45666
rect 54962 45614 54964 45666
rect 54908 45612 54964 45614
rect 55020 44492 55076 44548
rect 56588 47180 56644 47236
rect 56476 46732 56532 46788
rect 56476 46562 56532 46564
rect 56476 46510 56478 46562
rect 56478 46510 56530 46562
rect 56530 46510 56532 46562
rect 56476 46508 56532 46510
rect 56812 47458 56868 47460
rect 56812 47406 56814 47458
rect 56814 47406 56866 47458
rect 56866 47406 56868 47458
rect 56812 47404 56868 47406
rect 56700 46172 56756 46228
rect 57596 49868 57652 49924
rect 57260 47740 57316 47796
rect 56924 46508 56980 46564
rect 56588 46002 56644 46004
rect 56588 45950 56590 46002
rect 56590 45950 56642 46002
rect 56642 45950 56644 46002
rect 56588 45948 56644 45950
rect 56252 45164 56308 45220
rect 55804 42924 55860 42980
rect 54908 42642 54964 42644
rect 54908 42590 54910 42642
rect 54910 42590 54962 42642
rect 54962 42590 54964 42642
rect 54908 42588 54964 42590
rect 54684 42028 54740 42084
rect 53788 41804 53844 41860
rect 53900 41580 53956 41636
rect 54236 41468 54292 41524
rect 53676 41298 53732 41300
rect 53676 41246 53678 41298
rect 53678 41246 53730 41298
rect 53730 41246 53732 41298
rect 53676 41244 53732 41246
rect 53564 41132 53620 41188
rect 53564 40962 53620 40964
rect 53564 40910 53566 40962
rect 53566 40910 53618 40962
rect 53618 40910 53620 40962
rect 53564 40908 53620 40910
rect 53228 37436 53284 37492
rect 51996 35922 52052 35924
rect 51996 35870 51998 35922
rect 51998 35870 52050 35922
rect 52050 35870 52052 35922
rect 51996 35868 52052 35870
rect 51660 34914 51716 34916
rect 51660 34862 51662 34914
rect 51662 34862 51714 34914
rect 51714 34862 51716 34914
rect 51660 34860 51716 34862
rect 52108 34860 52164 34916
rect 49980 32508 50036 32564
rect 50428 32562 50484 32564
rect 50428 32510 50430 32562
rect 50430 32510 50482 32562
rect 50482 32510 50484 32562
rect 50428 32508 50484 32510
rect 50764 32562 50820 32564
rect 50764 32510 50766 32562
rect 50766 32510 50818 32562
rect 50818 32510 50820 32562
rect 50764 32508 50820 32510
rect 49756 31612 49812 31668
rect 49756 31106 49812 31108
rect 49756 31054 49758 31106
rect 49758 31054 49810 31106
rect 49810 31054 49812 31106
rect 49756 31052 49812 31054
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 49980 31052 50036 31108
rect 49868 30322 49924 30324
rect 49868 30270 49870 30322
rect 49870 30270 49922 30322
rect 49922 30270 49924 30322
rect 49868 30268 49924 30270
rect 50092 30044 50148 30100
rect 49644 27746 49700 27748
rect 49644 27694 49646 27746
rect 49646 27694 49698 27746
rect 49698 27694 49700 27746
rect 49644 27692 49700 27694
rect 49532 27186 49588 27188
rect 49532 27134 49534 27186
rect 49534 27134 49586 27186
rect 49586 27134 49588 27186
rect 49532 27132 49588 27134
rect 49756 27186 49812 27188
rect 49756 27134 49758 27186
rect 49758 27134 49810 27186
rect 49810 27134 49812 27186
rect 49756 27132 49812 27134
rect 49420 26178 49476 26180
rect 49420 26126 49422 26178
rect 49422 26126 49474 26178
rect 49474 26126 49476 26178
rect 49420 26124 49476 26126
rect 49196 25452 49252 25508
rect 48636 24946 48692 24948
rect 48636 24894 48638 24946
rect 48638 24894 48690 24946
rect 48690 24894 48692 24946
rect 48636 24892 48692 24894
rect 47964 24668 48020 24724
rect 47516 24220 47572 24276
rect 48748 24722 48804 24724
rect 48748 24670 48750 24722
rect 48750 24670 48802 24722
rect 48802 24670 48804 24722
rect 48748 24668 48804 24670
rect 47180 23660 47236 23716
rect 47516 23714 47572 23716
rect 47516 23662 47518 23714
rect 47518 23662 47570 23714
rect 47570 23662 47572 23714
rect 47516 23660 47572 23662
rect 48972 23660 49028 23716
rect 46396 22428 46452 22484
rect 46172 22146 46228 22148
rect 46172 22094 46174 22146
rect 46174 22094 46226 22146
rect 46226 22094 46228 22146
rect 46172 22092 46228 22094
rect 45948 21644 46004 21700
rect 44716 19122 44772 19124
rect 44716 19070 44718 19122
rect 44718 19070 44770 19122
rect 44770 19070 44772 19122
rect 44716 19068 44772 19070
rect 41804 18226 41860 18228
rect 41804 18174 41806 18226
rect 41806 18174 41858 18226
rect 41858 18174 41860 18226
rect 41804 18172 41860 18174
rect 43148 18396 43204 18452
rect 41468 17164 41524 17220
rect 41132 13916 41188 13972
rect 40572 12236 40628 12292
rect 40796 13356 40852 13412
rect 41804 15426 41860 15428
rect 41804 15374 41806 15426
rect 41806 15374 41858 15426
rect 41858 15374 41860 15426
rect 41804 15372 41860 15374
rect 41244 13356 41300 13412
rect 41356 14924 41412 14980
rect 40348 11900 40404 11956
rect 40460 11788 40516 11844
rect 40572 11340 40628 11396
rect 40124 10780 40180 10836
rect 41244 12962 41300 12964
rect 41244 12910 41246 12962
rect 41246 12910 41298 12962
rect 41298 12910 41300 12962
rect 41244 12908 41300 12910
rect 42476 17724 42532 17780
rect 42140 17164 42196 17220
rect 42364 15426 42420 15428
rect 42364 15374 42366 15426
rect 42366 15374 42418 15426
rect 42418 15374 42420 15426
rect 42364 15372 42420 15374
rect 41468 13356 41524 13412
rect 42028 13356 42084 13412
rect 41580 12348 41636 12404
rect 42028 12402 42084 12404
rect 42028 12350 42030 12402
rect 42030 12350 42082 12402
rect 42082 12350 42084 12402
rect 42028 12348 42084 12350
rect 41804 12290 41860 12292
rect 41804 12238 41806 12290
rect 41806 12238 41858 12290
rect 41858 12238 41860 12290
rect 41804 12236 41860 12238
rect 40796 11788 40852 11844
rect 41132 11900 41188 11956
rect 41580 11788 41636 11844
rect 38556 9884 38612 9940
rect 38892 10050 38948 10052
rect 38892 9998 38894 10050
rect 38894 9998 38946 10050
rect 38946 9998 38948 10050
rect 38892 9996 38948 9998
rect 38780 9042 38836 9044
rect 38780 8990 38782 9042
rect 38782 8990 38834 9042
rect 38834 8990 38836 9042
rect 38780 8988 38836 8990
rect 39340 9996 39396 10052
rect 40684 10834 40740 10836
rect 40684 10782 40686 10834
rect 40686 10782 40738 10834
rect 40738 10782 40740 10834
rect 40684 10780 40740 10782
rect 40348 9996 40404 10052
rect 40460 9884 40516 9940
rect 40012 9826 40068 9828
rect 40012 9774 40014 9826
rect 40014 9774 40066 9826
rect 40066 9774 40068 9826
rect 40012 9772 40068 9774
rect 40908 9826 40964 9828
rect 40908 9774 40910 9826
rect 40910 9774 40962 9826
rect 40962 9774 40964 9826
rect 40908 9772 40964 9774
rect 40684 9660 40740 9716
rect 41020 11228 41076 11284
rect 40460 9042 40516 9044
rect 40460 8990 40462 9042
rect 40462 8990 40514 9042
rect 40514 8990 40516 9042
rect 40460 8988 40516 8990
rect 39788 8204 39844 8260
rect 40124 8204 40180 8260
rect 39900 8034 39956 8036
rect 39900 7982 39902 8034
rect 39902 7982 39954 8034
rect 39954 7982 39956 8034
rect 39900 7980 39956 7982
rect 38556 7420 38612 7476
rect 39900 7474 39956 7476
rect 39900 7422 39902 7474
rect 39902 7422 39954 7474
rect 39954 7422 39956 7474
rect 39900 7420 39956 7422
rect 40796 8258 40852 8260
rect 40796 8206 40798 8258
rect 40798 8206 40850 8258
rect 40850 8206 40852 8258
rect 40796 8204 40852 8206
rect 40572 8034 40628 8036
rect 40572 7982 40574 8034
rect 40574 7982 40626 8034
rect 40626 7982 40628 8034
rect 40572 7980 40628 7982
rect 39452 5906 39508 5908
rect 39452 5854 39454 5906
rect 39454 5854 39506 5906
rect 39506 5854 39508 5906
rect 39452 5852 39508 5854
rect 38220 5180 38276 5236
rect 37660 5122 37716 5124
rect 37660 5070 37662 5122
rect 37662 5070 37714 5122
rect 37714 5070 37716 5122
rect 37660 5068 37716 5070
rect 38556 5122 38612 5124
rect 38556 5070 38558 5122
rect 38558 5070 38610 5122
rect 38610 5070 38612 5122
rect 38556 5068 38612 5070
rect 39228 5122 39284 5124
rect 39228 5070 39230 5122
rect 39230 5070 39282 5122
rect 39282 5070 39284 5122
rect 39228 5068 39284 5070
rect 39788 4898 39844 4900
rect 39788 4846 39790 4898
rect 39790 4846 39842 4898
rect 39842 4846 39844 4898
rect 39788 4844 39844 4846
rect 41020 7420 41076 7476
rect 42252 13356 42308 13412
rect 41692 9714 41748 9716
rect 41692 9662 41694 9714
rect 41694 9662 41746 9714
rect 41746 9662 41748 9714
rect 41692 9660 41748 9662
rect 41916 9996 41972 10052
rect 41916 9154 41972 9156
rect 41916 9102 41918 9154
rect 41918 9102 41970 9154
rect 41970 9102 41972 9154
rect 41916 9100 41972 9102
rect 42252 11900 42308 11956
rect 42364 11676 42420 11732
rect 42588 17164 42644 17220
rect 42812 18172 42868 18228
rect 43036 17612 43092 17668
rect 42812 17500 42868 17556
rect 42924 17052 42980 17108
rect 43596 18450 43652 18452
rect 43596 18398 43598 18450
rect 43598 18398 43650 18450
rect 43650 18398 43652 18450
rect 43596 18396 43652 18398
rect 43484 17724 43540 17780
rect 43820 17778 43876 17780
rect 43820 17726 43822 17778
rect 43822 17726 43874 17778
rect 43874 17726 43876 17778
rect 43820 17724 43876 17726
rect 43708 17666 43764 17668
rect 43708 17614 43710 17666
rect 43710 17614 43762 17666
rect 43762 17614 43764 17666
rect 43708 17612 43764 17614
rect 45500 18620 45556 18676
rect 44044 17276 44100 17332
rect 44492 18338 44548 18340
rect 44492 18286 44494 18338
rect 44494 18286 44546 18338
rect 44546 18286 44548 18338
rect 44492 18284 44548 18286
rect 44492 17778 44548 17780
rect 44492 17726 44494 17778
rect 44494 17726 44546 17778
rect 44546 17726 44548 17778
rect 44492 17724 44548 17726
rect 44380 17500 44436 17556
rect 45612 18508 45668 18564
rect 46060 20242 46116 20244
rect 46060 20190 46062 20242
rect 46062 20190 46114 20242
rect 46114 20190 46116 20242
rect 46060 20188 46116 20190
rect 45948 18284 46004 18340
rect 46060 19458 46116 19460
rect 46060 19406 46062 19458
rect 46062 19406 46114 19458
rect 46114 19406 46116 19458
rect 46060 19404 46116 19406
rect 43260 17106 43316 17108
rect 43260 17054 43262 17106
rect 43262 17054 43314 17106
rect 43314 17054 43316 17106
rect 43260 17052 43316 17054
rect 44268 17052 44324 17108
rect 43148 16940 43204 16996
rect 43484 16940 43540 16996
rect 42700 16828 42756 16884
rect 42924 16882 42980 16884
rect 42924 16830 42926 16882
rect 42926 16830 42978 16882
rect 42978 16830 42980 16882
rect 42924 16828 42980 16830
rect 42924 16044 42980 16100
rect 42588 15314 42644 15316
rect 42588 15262 42590 15314
rect 42590 15262 42642 15314
rect 42642 15262 42644 15314
rect 42588 15260 42644 15262
rect 42812 15986 42868 15988
rect 42812 15934 42814 15986
rect 42814 15934 42866 15986
rect 42866 15934 42868 15986
rect 42812 15932 42868 15934
rect 42700 14924 42756 14980
rect 43372 16098 43428 16100
rect 43372 16046 43374 16098
rect 43374 16046 43426 16098
rect 43426 16046 43428 16098
rect 43372 16044 43428 16046
rect 43820 16882 43876 16884
rect 43820 16830 43822 16882
rect 43822 16830 43874 16882
rect 43874 16830 43876 16882
rect 43820 16828 43876 16830
rect 43708 16604 43764 16660
rect 43708 15874 43764 15876
rect 43708 15822 43710 15874
rect 43710 15822 43762 15874
rect 43762 15822 43764 15874
rect 43708 15820 43764 15822
rect 43148 15372 43204 15428
rect 43036 13858 43092 13860
rect 43036 13806 43038 13858
rect 43038 13806 43090 13858
rect 43090 13806 43092 13858
rect 43036 13804 43092 13806
rect 43708 15426 43764 15428
rect 43708 15374 43710 15426
rect 43710 15374 43762 15426
rect 43762 15374 43764 15426
rect 43708 15372 43764 15374
rect 43484 15314 43540 15316
rect 43484 15262 43486 15314
rect 43486 15262 43538 15314
rect 43538 15262 43540 15314
rect 43484 15260 43540 15262
rect 43260 13356 43316 13412
rect 45164 17106 45220 17108
rect 45164 17054 45166 17106
rect 45166 17054 45218 17106
rect 45218 17054 45220 17106
rect 45164 17052 45220 17054
rect 45612 17106 45668 17108
rect 45612 17054 45614 17106
rect 45614 17054 45666 17106
rect 45666 17054 45668 17106
rect 45612 17052 45668 17054
rect 44716 16994 44772 16996
rect 44716 16942 44718 16994
rect 44718 16942 44770 16994
rect 44770 16942 44772 16994
rect 44716 16940 44772 16942
rect 44604 15986 44660 15988
rect 44604 15934 44606 15986
rect 44606 15934 44658 15986
rect 44658 15934 44660 15986
rect 44604 15932 44660 15934
rect 45052 15426 45108 15428
rect 45052 15374 45054 15426
rect 45054 15374 45106 15426
rect 45106 15374 45108 15426
rect 45052 15372 45108 15374
rect 45948 17052 46004 17108
rect 46732 22428 46788 22484
rect 47740 22258 47796 22260
rect 47740 22206 47742 22258
rect 47742 22206 47794 22258
rect 47794 22206 47796 22258
rect 47740 22204 47796 22206
rect 46844 21756 46900 21812
rect 46620 21084 46676 21140
rect 47628 22146 47684 22148
rect 47628 22094 47630 22146
rect 47630 22094 47682 22146
rect 47682 22094 47684 22146
rect 47628 22092 47684 22094
rect 48300 23042 48356 23044
rect 48300 22990 48302 23042
rect 48302 22990 48354 23042
rect 48354 22990 48356 23042
rect 48300 22988 48356 22990
rect 48188 22482 48244 22484
rect 48188 22430 48190 22482
rect 48190 22430 48242 22482
rect 48242 22430 48244 22482
rect 48188 22428 48244 22430
rect 47404 21810 47460 21812
rect 47404 21758 47406 21810
rect 47406 21758 47458 21810
rect 47458 21758 47460 21810
rect 47404 21756 47460 21758
rect 47292 21586 47348 21588
rect 47292 21534 47294 21586
rect 47294 21534 47346 21586
rect 47346 21534 47348 21586
rect 47292 21532 47348 21534
rect 47180 21084 47236 21140
rect 46508 20188 46564 20244
rect 47404 19122 47460 19124
rect 47404 19070 47406 19122
rect 47406 19070 47458 19122
rect 47458 19070 47460 19122
rect 47404 19068 47460 19070
rect 46508 18956 46564 19012
rect 47292 19010 47348 19012
rect 47292 18958 47294 19010
rect 47294 18958 47346 19010
rect 47346 18958 47348 19010
rect 47292 18956 47348 18958
rect 46620 17778 46676 17780
rect 46620 17726 46622 17778
rect 46622 17726 46674 17778
rect 46674 17726 46676 17778
rect 46620 17724 46676 17726
rect 47852 21084 47908 21140
rect 48300 20242 48356 20244
rect 48300 20190 48302 20242
rect 48302 20190 48354 20242
rect 48354 20190 48356 20242
rect 48300 20188 48356 20190
rect 48636 19180 48692 19236
rect 47516 17724 47572 17780
rect 47852 17612 47908 17668
rect 48076 18450 48132 18452
rect 48076 18398 48078 18450
rect 48078 18398 48130 18450
rect 48130 18398 48132 18450
rect 48076 18396 48132 18398
rect 46284 17052 46340 17108
rect 43708 13804 43764 13860
rect 44156 13804 44212 13860
rect 42588 12290 42644 12292
rect 42588 12238 42590 12290
rect 42590 12238 42642 12290
rect 42642 12238 42644 12290
rect 42588 12236 42644 12238
rect 42812 11676 42868 11732
rect 43596 12348 43652 12404
rect 43596 11676 43652 11732
rect 43484 11452 43540 11508
rect 42924 11170 42980 11172
rect 42924 11118 42926 11170
rect 42926 11118 42978 11170
rect 42978 11118 42980 11170
rect 42924 11116 42980 11118
rect 43708 11116 43764 11172
rect 42028 9436 42084 9492
rect 42252 9324 42308 9380
rect 43036 9826 43092 9828
rect 43036 9774 43038 9826
rect 43038 9774 43090 9826
rect 43090 9774 43092 9826
rect 43036 9772 43092 9774
rect 43036 9548 43092 9604
rect 43260 9660 43316 9716
rect 42028 8988 42084 9044
rect 42588 9100 42644 9156
rect 42028 8204 42084 8260
rect 43148 9324 43204 9380
rect 43260 9212 43316 9268
rect 43708 9100 43764 9156
rect 43932 12402 43988 12404
rect 43932 12350 43934 12402
rect 43934 12350 43986 12402
rect 43986 12350 43988 12402
rect 43932 12348 43988 12350
rect 43932 11564 43988 11620
rect 44044 11452 44100 11508
rect 44716 14642 44772 14644
rect 44716 14590 44718 14642
rect 44718 14590 44770 14642
rect 44770 14590 44772 14642
rect 44716 14588 44772 14590
rect 45724 14028 45780 14084
rect 45612 13634 45668 13636
rect 45612 13582 45614 13634
rect 45614 13582 45666 13634
rect 45666 13582 45668 13634
rect 45612 13580 45668 13582
rect 45164 11452 45220 11508
rect 45500 11506 45556 11508
rect 45500 11454 45502 11506
rect 45502 11454 45554 11506
rect 45554 11454 45556 11506
rect 45500 11452 45556 11454
rect 44604 11394 44660 11396
rect 44604 11342 44606 11394
rect 44606 11342 44658 11394
rect 44658 11342 44660 11394
rect 44604 11340 44660 11342
rect 42700 8258 42756 8260
rect 42700 8206 42702 8258
rect 42702 8206 42754 8258
rect 42754 8206 42756 8258
rect 42700 8204 42756 8206
rect 40908 5292 40964 5348
rect 41468 5346 41524 5348
rect 41468 5294 41470 5346
rect 41470 5294 41522 5346
rect 41522 5294 41524 5346
rect 41468 5292 41524 5294
rect 43148 8370 43204 8372
rect 43148 8318 43150 8370
rect 43150 8318 43202 8370
rect 43202 8318 43204 8370
rect 43148 8316 43204 8318
rect 43036 8204 43092 8260
rect 43148 7474 43204 7476
rect 43148 7422 43150 7474
rect 43150 7422 43202 7474
rect 43202 7422 43204 7474
rect 43148 7420 43204 7422
rect 45724 11394 45780 11396
rect 45724 11342 45726 11394
rect 45726 11342 45778 11394
rect 45778 11342 45780 11394
rect 45724 11340 45780 11342
rect 45948 15426 46004 15428
rect 45948 15374 45950 15426
rect 45950 15374 46002 15426
rect 46002 15374 46004 15426
rect 45948 15372 46004 15374
rect 47292 15202 47348 15204
rect 47292 15150 47294 15202
rect 47294 15150 47346 15202
rect 47346 15150 47348 15202
rect 47292 15148 47348 15150
rect 46508 14642 46564 14644
rect 46508 14590 46510 14642
rect 46510 14590 46562 14642
rect 46562 14590 46564 14642
rect 46508 14588 46564 14590
rect 50764 30098 50820 30100
rect 50764 30046 50766 30098
rect 50766 30046 50818 30098
rect 50818 30046 50820 30098
rect 50764 30044 50820 30046
rect 51212 32508 51268 32564
rect 51548 31106 51604 31108
rect 51548 31054 51550 31106
rect 51550 31054 51602 31106
rect 51602 31054 51604 31106
rect 51548 31052 51604 31054
rect 51772 30828 51828 30884
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 50428 28642 50484 28644
rect 50428 28590 50430 28642
rect 50430 28590 50482 28642
rect 50482 28590 50484 28642
rect 50428 28588 50484 28590
rect 50876 28588 50932 28644
rect 50092 27692 50148 27748
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 50652 27804 50708 27860
rect 50428 27186 50484 27188
rect 50428 27134 50430 27186
rect 50430 27134 50482 27186
rect 50482 27134 50484 27186
rect 50428 27132 50484 27134
rect 50652 27298 50708 27300
rect 50652 27246 50654 27298
rect 50654 27246 50706 27298
rect 50706 27246 50708 27298
rect 50652 27244 50708 27246
rect 51100 27858 51156 27860
rect 51100 27806 51102 27858
rect 51102 27806 51154 27858
rect 51154 27806 51156 27858
rect 51100 27804 51156 27806
rect 51100 27580 51156 27636
rect 51324 30604 51380 30660
rect 51212 27468 51268 27524
rect 51212 27186 51268 27188
rect 51212 27134 51214 27186
rect 51214 27134 51266 27186
rect 51266 27134 51268 27186
rect 51212 27132 51268 27134
rect 50540 26908 50596 26964
rect 51324 26962 51380 26964
rect 51324 26910 51326 26962
rect 51326 26910 51378 26962
rect 51378 26910 51380 26962
rect 51324 26908 51380 26910
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 49868 26178 49924 26180
rect 49868 26126 49870 26178
rect 49870 26126 49922 26178
rect 49922 26126 49924 26178
rect 49868 26124 49924 26126
rect 50540 26124 50596 26180
rect 49420 25452 49476 25508
rect 49756 24668 49812 24724
rect 50540 25564 50596 25620
rect 51324 25618 51380 25620
rect 51324 25566 51326 25618
rect 51326 25566 51378 25618
rect 51378 25566 51380 25618
rect 51324 25564 51380 25566
rect 50764 25506 50820 25508
rect 50764 25454 50766 25506
rect 50766 25454 50818 25506
rect 50818 25454 50820 25506
rect 50764 25452 50820 25454
rect 49980 24946 50036 24948
rect 49980 24894 49982 24946
rect 49982 24894 50034 24946
rect 50034 24894 50036 24946
rect 49980 24892 50036 24894
rect 50876 25394 50932 25396
rect 50876 25342 50878 25394
rect 50878 25342 50930 25394
rect 50930 25342 50932 25394
rect 50876 25340 50932 25342
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 49308 23324 49364 23380
rect 49196 22988 49252 23044
rect 49308 21644 49364 21700
rect 49644 21644 49700 21700
rect 49868 21586 49924 21588
rect 49868 21534 49870 21586
rect 49870 21534 49922 21586
rect 49922 21534 49924 21586
rect 49868 21532 49924 21534
rect 49644 21308 49700 21364
rect 49084 19234 49140 19236
rect 49084 19182 49086 19234
rect 49086 19182 49138 19234
rect 49138 19182 49140 19234
rect 49084 19180 49140 19182
rect 49196 19122 49252 19124
rect 49196 19070 49198 19122
rect 49198 19070 49250 19122
rect 49250 19070 49252 19122
rect 49196 19068 49252 19070
rect 48972 17890 49028 17892
rect 48972 17838 48974 17890
rect 48974 17838 49026 17890
rect 49026 17838 49028 17890
rect 48972 17836 49028 17838
rect 48748 17724 48804 17780
rect 48860 17666 48916 17668
rect 48860 17614 48862 17666
rect 48862 17614 48914 17666
rect 48914 17614 48916 17666
rect 48860 17612 48916 17614
rect 48076 17500 48132 17556
rect 48972 17554 49028 17556
rect 48972 17502 48974 17554
rect 48974 17502 49026 17554
rect 49026 17502 49028 17554
rect 48972 17500 49028 17502
rect 48636 15820 48692 15876
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 50540 22370 50596 22372
rect 50540 22318 50542 22370
rect 50542 22318 50594 22370
rect 50594 22318 50596 22370
rect 50540 22316 50596 22318
rect 51324 23266 51380 23268
rect 51324 23214 51326 23266
rect 51326 23214 51378 23266
rect 51378 23214 51380 23266
rect 51324 23212 51380 23214
rect 51100 22316 51156 22372
rect 51212 22258 51268 22260
rect 51212 22206 51214 22258
rect 51214 22206 51266 22258
rect 51266 22206 51268 22258
rect 51212 22204 51268 22206
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 50540 21698 50596 21700
rect 50540 21646 50542 21698
rect 50542 21646 50594 21698
rect 50594 21646 50596 21698
rect 50540 21644 50596 21646
rect 51100 21586 51156 21588
rect 51100 21534 51102 21586
rect 51102 21534 51154 21586
rect 51154 21534 51156 21586
rect 51100 21532 51156 21534
rect 51324 21362 51380 21364
rect 51324 21310 51326 21362
rect 51326 21310 51378 21362
rect 51378 21310 51380 21362
rect 51324 21308 51380 21310
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 50316 20076 50372 20132
rect 50092 19180 50148 19236
rect 49980 19068 50036 19124
rect 51772 27746 51828 27748
rect 51772 27694 51774 27746
rect 51774 27694 51826 27746
rect 51826 27694 51828 27746
rect 51772 27692 51828 27694
rect 51772 27468 51828 27524
rect 52108 34354 52164 34356
rect 52108 34302 52110 34354
rect 52110 34302 52162 34354
rect 52162 34302 52164 34354
rect 52108 34300 52164 34302
rect 53564 39506 53620 39508
rect 53564 39454 53566 39506
rect 53566 39454 53618 39506
rect 53618 39454 53620 39506
rect 53564 39452 53620 39454
rect 53564 38892 53620 38948
rect 53900 38722 53956 38724
rect 53900 38670 53902 38722
rect 53902 38670 53954 38722
rect 53954 38670 53956 38722
rect 53900 38668 53956 38670
rect 54348 41692 54404 41748
rect 54572 41746 54628 41748
rect 54572 41694 54574 41746
rect 54574 41694 54626 41746
rect 54626 41694 54628 41746
rect 54572 41692 54628 41694
rect 54460 41244 54516 41300
rect 55468 42476 55524 42532
rect 54460 40908 54516 40964
rect 55916 42476 55972 42532
rect 55916 42140 55972 42196
rect 56700 45164 56756 45220
rect 56700 44546 56756 44548
rect 56700 44494 56702 44546
rect 56702 44494 56754 44546
rect 56754 44494 56756 44546
rect 56700 44492 56756 44494
rect 56588 43762 56644 43764
rect 56588 43710 56590 43762
rect 56590 43710 56642 43762
rect 56642 43710 56644 43762
rect 56588 43708 56644 43710
rect 56476 43538 56532 43540
rect 56476 43486 56478 43538
rect 56478 43486 56530 43538
rect 56530 43486 56532 43538
rect 56476 43484 56532 43486
rect 56812 43484 56868 43540
rect 57484 48748 57540 48804
rect 58268 49026 58324 49028
rect 58268 48974 58270 49026
rect 58270 48974 58322 49026
rect 58322 48974 58324 49026
rect 58268 48972 58324 48974
rect 57932 48242 57988 48244
rect 57932 48190 57934 48242
rect 57934 48190 57986 48242
rect 57986 48190 57988 48242
rect 57932 48188 57988 48190
rect 58492 49922 58548 49924
rect 58492 49870 58494 49922
rect 58494 49870 58546 49922
rect 58546 49870 58548 49922
rect 58492 49868 58548 49870
rect 58380 48188 58436 48244
rect 57596 47740 57652 47796
rect 57372 47404 57428 47460
rect 57484 47180 57540 47236
rect 56476 42924 56532 42980
rect 56140 42530 56196 42532
rect 56140 42478 56142 42530
rect 56142 42478 56194 42530
rect 56194 42478 56196 42530
rect 56140 42476 56196 42478
rect 56364 42476 56420 42532
rect 56364 42028 56420 42084
rect 55020 40908 55076 40964
rect 55804 40962 55860 40964
rect 55804 40910 55806 40962
rect 55806 40910 55858 40962
rect 55858 40910 55860 40962
rect 55804 40908 55860 40910
rect 54684 39506 54740 39508
rect 54684 39454 54686 39506
rect 54686 39454 54738 39506
rect 54738 39454 54740 39506
rect 54684 39452 54740 39454
rect 54572 38668 54628 38724
rect 55580 38722 55636 38724
rect 55580 38670 55582 38722
rect 55582 38670 55634 38722
rect 55634 38670 55636 38722
rect 55580 38668 55636 38670
rect 54908 37938 54964 37940
rect 54908 37886 54910 37938
rect 54910 37886 54962 37938
rect 54962 37886 54964 37938
rect 54908 37884 54964 37886
rect 54348 37490 54404 37492
rect 54348 37438 54350 37490
rect 54350 37438 54402 37490
rect 54402 37438 54404 37490
rect 54348 37436 54404 37438
rect 57036 45948 57092 46004
rect 56700 42140 56756 42196
rect 57484 43708 57540 43764
rect 57260 43484 57316 43540
rect 56588 41356 56644 41412
rect 57820 45106 57876 45108
rect 57820 45054 57822 45106
rect 57822 45054 57874 45106
rect 57874 45054 57876 45106
rect 57820 45052 57876 45054
rect 57708 44434 57764 44436
rect 57708 44382 57710 44434
rect 57710 44382 57762 44434
rect 57762 44382 57764 44434
rect 57708 44380 57764 44382
rect 58492 45106 58548 45108
rect 58492 45054 58494 45106
rect 58494 45054 58546 45106
rect 58546 45054 58548 45106
rect 58492 45052 58548 45054
rect 57484 42082 57540 42084
rect 57484 42030 57486 42082
rect 57486 42030 57538 42082
rect 57538 42030 57540 42082
rect 57484 42028 57540 42030
rect 57372 41356 57428 41412
rect 57036 40908 57092 40964
rect 56812 39564 56868 39620
rect 56700 38834 56756 38836
rect 56700 38782 56702 38834
rect 56702 38782 56754 38834
rect 56754 38782 56756 38834
rect 56700 38780 56756 38782
rect 56364 38722 56420 38724
rect 56364 38670 56366 38722
rect 56366 38670 56418 38722
rect 56418 38670 56420 38722
rect 56364 38668 56420 38670
rect 55244 37436 55300 37492
rect 53004 35698 53060 35700
rect 53004 35646 53006 35698
rect 53006 35646 53058 35698
rect 53058 35646 53060 35698
rect 53004 35644 53060 35646
rect 52556 34914 52612 34916
rect 52556 34862 52558 34914
rect 52558 34862 52610 34914
rect 52610 34862 52612 34914
rect 52556 34860 52612 34862
rect 52668 34354 52724 34356
rect 52668 34302 52670 34354
rect 52670 34302 52722 34354
rect 52722 34302 52724 34354
rect 52668 34300 52724 34302
rect 53676 35644 53732 35700
rect 53228 35196 53284 35252
rect 53564 34914 53620 34916
rect 53564 34862 53566 34914
rect 53566 34862 53618 34914
rect 53618 34862 53620 34914
rect 53564 34860 53620 34862
rect 53900 35810 53956 35812
rect 53900 35758 53902 35810
rect 53902 35758 53954 35810
rect 53954 35758 53956 35810
rect 53900 35756 53956 35758
rect 54012 34860 54068 34916
rect 53788 34748 53844 34804
rect 54796 35756 54852 35812
rect 55580 35698 55636 35700
rect 55580 35646 55582 35698
rect 55582 35646 55634 35698
rect 55634 35646 55636 35698
rect 55580 35644 55636 35646
rect 54460 33404 54516 33460
rect 52668 31666 52724 31668
rect 52668 31614 52670 31666
rect 52670 31614 52722 31666
rect 52722 31614 52724 31666
rect 52668 31612 52724 31614
rect 52780 31218 52836 31220
rect 52780 31166 52782 31218
rect 52782 31166 52834 31218
rect 52834 31166 52836 31218
rect 52780 31164 52836 31166
rect 52444 31106 52500 31108
rect 52444 31054 52446 31106
rect 52446 31054 52498 31106
rect 52498 31054 52500 31106
rect 52444 31052 52500 31054
rect 52556 30828 52612 30884
rect 52668 30940 52724 30996
rect 53116 30882 53172 30884
rect 53116 30830 53118 30882
rect 53118 30830 53170 30882
rect 53170 30830 53172 30882
rect 53116 30828 53172 30830
rect 52668 30210 52724 30212
rect 52668 30158 52670 30210
rect 52670 30158 52722 30210
rect 52722 30158 52724 30210
rect 52668 30156 52724 30158
rect 52108 30044 52164 30100
rect 53004 29538 53060 29540
rect 53004 29486 53006 29538
rect 53006 29486 53058 29538
rect 53058 29486 53060 29538
rect 53004 29484 53060 29486
rect 52668 28866 52724 28868
rect 52668 28814 52670 28866
rect 52670 28814 52722 28866
rect 52722 28814 52724 28866
rect 52668 28812 52724 28814
rect 52108 28642 52164 28644
rect 52108 28590 52110 28642
rect 52110 28590 52162 28642
rect 52162 28590 52164 28642
rect 52108 28588 52164 28590
rect 52444 27746 52500 27748
rect 52444 27694 52446 27746
rect 52446 27694 52498 27746
rect 52498 27694 52500 27746
rect 52444 27692 52500 27694
rect 52108 27020 52164 27076
rect 51996 26962 52052 26964
rect 51996 26910 51998 26962
rect 51998 26910 52050 26962
rect 52050 26910 52052 26962
rect 51996 26908 52052 26910
rect 52668 26908 52724 26964
rect 52780 27074 52836 27076
rect 52780 27022 52782 27074
rect 52782 27022 52834 27074
rect 52834 27022 52836 27074
rect 52780 27020 52836 27022
rect 51884 24780 51940 24836
rect 52780 25228 52836 25284
rect 53340 31164 53396 31220
rect 54796 32508 54852 32564
rect 55356 32562 55412 32564
rect 55356 32510 55358 32562
rect 55358 32510 55410 32562
rect 55410 32510 55412 32562
rect 55356 32508 55412 32510
rect 53900 31948 53956 32004
rect 54460 31890 54516 31892
rect 54460 31838 54462 31890
rect 54462 31838 54514 31890
rect 54514 31838 54516 31890
rect 54460 31836 54516 31838
rect 54796 31836 54852 31892
rect 54012 31666 54068 31668
rect 54012 31614 54014 31666
rect 54014 31614 54066 31666
rect 54066 31614 54068 31666
rect 54012 31612 54068 31614
rect 53676 30210 53732 30212
rect 53676 30158 53678 30210
rect 53678 30158 53730 30210
rect 53730 30158 53732 30210
rect 53676 30156 53732 30158
rect 55132 31836 55188 31892
rect 55468 31890 55524 31892
rect 55468 31838 55470 31890
rect 55470 31838 55522 31890
rect 55522 31838 55524 31890
rect 55468 31836 55524 31838
rect 55244 31500 55300 31556
rect 54124 29484 54180 29540
rect 53452 28812 53508 28868
rect 54908 30156 54964 30212
rect 55468 30210 55524 30212
rect 55468 30158 55470 30210
rect 55470 30158 55522 30210
rect 55522 30158 55524 30210
rect 55468 30156 55524 30158
rect 54572 29314 54628 29316
rect 54572 29262 54574 29314
rect 54574 29262 54626 29314
rect 54626 29262 54628 29314
rect 54572 29260 54628 29262
rect 53564 28700 53620 28756
rect 54348 29036 54404 29092
rect 55132 29036 55188 29092
rect 55356 29314 55412 29316
rect 55356 29262 55358 29314
rect 55358 29262 55410 29314
rect 55410 29262 55412 29314
rect 55356 29260 55412 29262
rect 55356 28588 55412 28644
rect 55020 28476 55076 28532
rect 55020 27132 55076 27188
rect 53676 27074 53732 27076
rect 53676 27022 53678 27074
rect 53678 27022 53730 27074
rect 53730 27022 53732 27074
rect 53676 27020 53732 27022
rect 53676 26850 53732 26852
rect 53676 26798 53678 26850
rect 53678 26798 53730 26850
rect 53730 26798 53732 26850
rect 53676 26796 53732 26798
rect 53676 26066 53732 26068
rect 53676 26014 53678 26066
rect 53678 26014 53730 26066
rect 53730 26014 53732 26066
rect 53676 26012 53732 26014
rect 54348 26066 54404 26068
rect 54348 26014 54350 26066
rect 54350 26014 54402 26066
rect 54402 26014 54404 26066
rect 54348 26012 54404 26014
rect 53900 25506 53956 25508
rect 53900 25454 53902 25506
rect 53902 25454 53954 25506
rect 53954 25454 53956 25506
rect 53900 25452 53956 25454
rect 56252 35868 56308 35924
rect 56364 35644 56420 35700
rect 56700 35644 56756 35700
rect 56476 33458 56532 33460
rect 56476 33406 56478 33458
rect 56478 33406 56530 33458
rect 56530 33406 56532 33458
rect 56476 33404 56532 33406
rect 56924 32508 56980 32564
rect 55692 29372 55748 29428
rect 55692 29202 55748 29204
rect 55692 29150 55694 29202
rect 55694 29150 55746 29202
rect 55746 29150 55748 29202
rect 55692 29148 55748 29150
rect 54572 25452 54628 25508
rect 52668 23772 52724 23828
rect 53228 24610 53284 24612
rect 53228 24558 53230 24610
rect 53230 24558 53282 24610
rect 53282 24558 53284 24610
rect 53228 24556 53284 24558
rect 53004 23772 53060 23828
rect 51996 22258 52052 22260
rect 51996 22206 51998 22258
rect 51998 22206 52050 22258
rect 52050 22206 52052 22258
rect 51996 22204 52052 22206
rect 52220 22258 52276 22260
rect 52220 22206 52222 22258
rect 52222 22206 52274 22258
rect 52274 22206 52276 22258
rect 52220 22204 52276 22206
rect 52332 21644 52388 21700
rect 52108 21308 52164 21364
rect 51436 19180 51492 19236
rect 50428 19010 50484 19012
rect 50428 18958 50430 19010
rect 50430 18958 50482 19010
rect 50482 18958 50484 19010
rect 50428 18956 50484 18958
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 50316 18226 50372 18228
rect 50316 18174 50318 18226
rect 50318 18174 50370 18226
rect 50370 18174 50372 18226
rect 50316 18172 50372 18174
rect 49980 17778 50036 17780
rect 49980 17726 49982 17778
rect 49982 17726 50034 17778
rect 50034 17726 50036 17778
rect 49980 17724 50036 17726
rect 50876 18172 50932 18228
rect 52892 19906 52948 19908
rect 52892 19854 52894 19906
rect 52894 19854 52946 19906
rect 52946 19854 52948 19906
rect 52892 19852 52948 19854
rect 52220 19068 52276 19124
rect 52668 19122 52724 19124
rect 52668 19070 52670 19122
rect 52670 19070 52722 19122
rect 52722 19070 52724 19122
rect 52668 19068 52724 19070
rect 51436 19010 51492 19012
rect 51436 18958 51438 19010
rect 51438 18958 51490 19010
rect 51490 18958 51492 19010
rect 51436 18956 51492 18958
rect 52780 18562 52836 18564
rect 52780 18510 52782 18562
rect 52782 18510 52834 18562
rect 52834 18510 52836 18562
rect 52780 18508 52836 18510
rect 52108 17836 52164 17892
rect 52332 17836 52388 17892
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 55132 24780 55188 24836
rect 54012 23212 54068 23268
rect 53564 23100 53620 23156
rect 53452 23042 53508 23044
rect 53452 22990 53454 23042
rect 53454 22990 53506 23042
rect 53506 22990 53508 23042
rect 53452 22988 53508 22990
rect 53564 22204 53620 22260
rect 53788 22988 53844 23044
rect 54460 23212 54516 23268
rect 54348 23154 54404 23156
rect 54348 23102 54350 23154
rect 54350 23102 54402 23154
rect 54402 23102 54404 23154
rect 54348 23100 54404 23102
rect 54460 23042 54516 23044
rect 54460 22990 54462 23042
rect 54462 22990 54514 23042
rect 54514 22990 54516 23042
rect 54460 22988 54516 22990
rect 56028 29484 56084 29540
rect 56140 29036 56196 29092
rect 56588 30716 56644 30772
rect 56812 30716 56868 30772
rect 56364 28924 56420 28980
rect 56364 28642 56420 28644
rect 56364 28590 56366 28642
rect 56366 28590 56418 28642
rect 56418 28590 56420 28642
rect 56364 28588 56420 28590
rect 56476 26796 56532 26852
rect 56028 25394 56084 25396
rect 56028 25342 56030 25394
rect 56030 25342 56082 25394
rect 56082 25342 56084 25394
rect 56028 25340 56084 25342
rect 55580 24834 55636 24836
rect 55580 24782 55582 24834
rect 55582 24782 55634 24834
rect 55634 24782 55636 24834
rect 55580 24780 55636 24782
rect 55132 23826 55188 23828
rect 55132 23774 55134 23826
rect 55134 23774 55186 23826
rect 55186 23774 55188 23826
rect 55132 23772 55188 23774
rect 56700 28924 56756 28980
rect 56700 26290 56756 26292
rect 56700 26238 56702 26290
rect 56702 26238 56754 26290
rect 56754 26238 56756 26290
rect 56700 26236 56756 26238
rect 56924 26236 56980 26292
rect 57148 41186 57204 41188
rect 57148 41134 57150 41186
rect 57150 41134 57202 41186
rect 57202 41134 57204 41186
rect 57148 41132 57204 41134
rect 57596 41132 57652 41188
rect 57932 41356 57988 41412
rect 57708 40514 57764 40516
rect 57708 40462 57710 40514
rect 57710 40462 57762 40514
rect 57762 40462 57764 40514
rect 57708 40460 57764 40462
rect 58268 40236 58324 40292
rect 57596 38722 57652 38724
rect 57596 38670 57598 38722
rect 57598 38670 57650 38722
rect 57650 38670 57652 38722
rect 57596 38668 57652 38670
rect 57820 39618 57876 39620
rect 57820 39566 57822 39618
rect 57822 39566 57874 39618
rect 57874 39566 57876 39618
rect 57820 39564 57876 39566
rect 58268 39564 58324 39620
rect 57932 38834 57988 38836
rect 57932 38782 57934 38834
rect 57934 38782 57986 38834
rect 57986 38782 57988 38834
rect 57932 38780 57988 38782
rect 57708 36092 57764 36148
rect 58044 35980 58100 36036
rect 57932 35698 57988 35700
rect 57932 35646 57934 35698
rect 57934 35646 57986 35698
rect 57986 35646 57988 35698
rect 57932 35644 57988 35646
rect 57372 31948 57428 32004
rect 57820 32562 57876 32564
rect 57820 32510 57822 32562
rect 57822 32510 57874 32562
rect 57874 32510 57876 32562
rect 57820 32508 57876 32510
rect 57372 30716 57428 30772
rect 57484 29538 57540 29540
rect 57484 29486 57486 29538
rect 57486 29486 57538 29538
rect 57538 29486 57540 29538
rect 57484 29484 57540 29486
rect 57260 28924 57316 28980
rect 57708 30770 57764 30772
rect 57708 30718 57710 30770
rect 57710 30718 57762 30770
rect 57762 30718 57764 30770
rect 57708 30716 57764 30718
rect 58044 29148 58100 29204
rect 57708 28924 57764 28980
rect 56252 24892 56308 24948
rect 57932 26796 57988 26852
rect 57596 26290 57652 26292
rect 57596 26238 57598 26290
rect 57598 26238 57650 26290
rect 57650 26238 57652 26290
rect 57596 26236 57652 26238
rect 56364 23772 56420 23828
rect 54348 21308 54404 21364
rect 54796 21308 54852 21364
rect 54684 20690 54740 20692
rect 54684 20638 54686 20690
rect 54686 20638 54738 20690
rect 54738 20638 54740 20690
rect 54684 20636 54740 20638
rect 53676 20412 53732 20468
rect 53788 20076 53844 20132
rect 54460 19852 54516 19908
rect 56364 22092 56420 22148
rect 55356 21308 55412 21364
rect 55020 20412 55076 20468
rect 56028 20690 56084 20692
rect 56028 20638 56030 20690
rect 56030 20638 56082 20690
rect 56082 20638 56084 20690
rect 56028 20636 56084 20638
rect 53788 19740 53844 19796
rect 54012 19740 54068 19796
rect 53788 19180 53844 19236
rect 53452 19068 53508 19124
rect 53564 18620 53620 18676
rect 53452 18508 53508 18564
rect 53900 19122 53956 19124
rect 53900 19070 53902 19122
rect 53902 19070 53954 19122
rect 53954 19070 53956 19122
rect 53900 19068 53956 19070
rect 54348 19234 54404 19236
rect 54348 19182 54350 19234
rect 54350 19182 54402 19234
rect 54402 19182 54404 19234
rect 54348 19180 54404 19182
rect 54012 18620 54068 18676
rect 54124 18396 54180 18452
rect 55692 19964 55748 20020
rect 55020 19906 55076 19908
rect 55020 19854 55022 19906
rect 55022 19854 55074 19906
rect 55074 19854 55076 19906
rect 55020 19852 55076 19854
rect 55468 19234 55524 19236
rect 55468 19182 55470 19234
rect 55470 19182 55522 19234
rect 55522 19182 55524 19234
rect 55468 19180 55524 19182
rect 55356 19122 55412 19124
rect 55356 19070 55358 19122
rect 55358 19070 55410 19122
rect 55410 19070 55412 19122
rect 55356 19068 55412 19070
rect 56028 19852 56084 19908
rect 56588 21420 56644 21476
rect 56476 21362 56532 21364
rect 56476 21310 56478 21362
rect 56478 21310 56530 21362
rect 56530 21310 56532 21362
rect 56476 21308 56532 21310
rect 56140 19180 56196 19236
rect 55580 19068 55636 19124
rect 56028 18508 56084 18564
rect 55916 18396 55972 18452
rect 53788 17276 53844 17332
rect 49756 15820 49812 15876
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 49196 15372 49252 15428
rect 48412 15202 48468 15204
rect 48412 15150 48414 15202
rect 48414 15150 48466 15202
rect 48466 15150 48468 15202
rect 48412 15148 48468 15150
rect 46956 14588 47012 14644
rect 46060 14028 46116 14084
rect 46620 14028 46676 14084
rect 45948 13580 46004 13636
rect 46396 13580 46452 13636
rect 46060 13020 46116 13076
rect 46844 13580 46900 13636
rect 49980 15426 50036 15428
rect 49980 15374 49982 15426
rect 49982 15374 50034 15426
rect 50034 15374 50036 15426
rect 49980 15372 50036 15374
rect 49644 15314 49700 15316
rect 49644 15262 49646 15314
rect 49646 15262 49698 15314
rect 49698 15262 49700 15314
rect 49644 15260 49700 15262
rect 49532 15148 49588 15204
rect 48748 14588 48804 14644
rect 49644 14642 49700 14644
rect 49644 14590 49646 14642
rect 49646 14590 49698 14642
rect 49698 14590 49700 14642
rect 49644 14588 49700 14590
rect 52444 15986 52500 15988
rect 52444 15934 52446 15986
rect 52446 15934 52498 15986
rect 52498 15934 52500 15986
rect 52444 15932 52500 15934
rect 52668 15932 52724 15988
rect 53452 15986 53508 15988
rect 53452 15934 53454 15986
rect 53454 15934 53506 15986
rect 53506 15934 53508 15986
rect 53452 15932 53508 15934
rect 52556 15874 52612 15876
rect 52556 15822 52558 15874
rect 52558 15822 52610 15874
rect 52610 15822 52612 15874
rect 52556 15820 52612 15822
rect 50876 14700 50932 14756
rect 51884 14754 51940 14756
rect 51884 14702 51886 14754
rect 51886 14702 51938 14754
rect 51938 14702 51940 14754
rect 51884 14700 51940 14702
rect 52668 15314 52724 15316
rect 52668 15262 52670 15314
rect 52670 15262 52722 15314
rect 52722 15262 52724 15314
rect 52668 15260 52724 15262
rect 52332 14700 52388 14756
rect 47292 13020 47348 13076
rect 47740 14028 47796 14084
rect 48188 14028 48244 14084
rect 47628 13580 47684 13636
rect 47628 12402 47684 12404
rect 47628 12350 47630 12402
rect 47630 12350 47682 12402
rect 47682 12350 47684 12402
rect 47628 12348 47684 12350
rect 44268 10050 44324 10052
rect 44268 9998 44270 10050
rect 44270 9998 44322 10050
rect 44322 9998 44324 10050
rect 44268 9996 44324 9998
rect 44604 9826 44660 9828
rect 44604 9774 44606 9826
rect 44606 9774 44658 9826
rect 44658 9774 44660 9826
rect 44604 9772 44660 9774
rect 44268 9660 44324 9716
rect 44156 9548 44212 9604
rect 44156 9100 44212 9156
rect 43932 8316 43988 8372
rect 44716 9154 44772 9156
rect 44716 9102 44718 9154
rect 44718 9102 44770 9154
rect 44770 9102 44772 9154
rect 44716 9100 44772 9102
rect 44940 9154 44996 9156
rect 44940 9102 44942 9154
rect 44942 9102 44994 9154
rect 44994 9102 44996 9154
rect 44940 9100 44996 9102
rect 45836 11228 45892 11284
rect 45612 9996 45668 10052
rect 45164 9772 45220 9828
rect 45388 9602 45444 9604
rect 45388 9550 45390 9602
rect 45390 9550 45442 9602
rect 45442 9550 45444 9602
rect 45388 9548 45444 9550
rect 47068 11282 47124 11284
rect 47068 11230 47070 11282
rect 47070 11230 47122 11282
rect 47122 11230 47124 11282
rect 47068 11228 47124 11230
rect 46732 11170 46788 11172
rect 46732 11118 46734 11170
rect 46734 11118 46786 11170
rect 46786 11118 46788 11170
rect 46732 11116 46788 11118
rect 46844 11004 46900 11060
rect 47068 9826 47124 9828
rect 47068 9774 47070 9826
rect 47070 9774 47122 9826
rect 47122 9774 47124 9826
rect 47068 9772 47124 9774
rect 43932 7644 43988 7700
rect 44492 7698 44548 7700
rect 44492 7646 44494 7698
rect 44494 7646 44546 7698
rect 44546 7646 44548 7698
rect 44492 7644 44548 7646
rect 43820 7420 43876 7476
rect 42476 5964 42532 6020
rect 40124 4508 40180 4564
rect 40572 4844 40628 4900
rect 41804 5122 41860 5124
rect 41804 5070 41806 5122
rect 41806 5070 41858 5122
rect 41858 5070 41860 5122
rect 41804 5068 41860 5070
rect 41916 5010 41972 5012
rect 41916 4958 41918 5010
rect 41918 4958 41970 5010
rect 41970 4958 41972 5010
rect 41916 4956 41972 4958
rect 41692 4844 41748 4900
rect 40684 4562 40740 4564
rect 40684 4510 40686 4562
rect 40686 4510 40738 4562
rect 40738 4510 40740 4562
rect 40684 4508 40740 4510
rect 42924 5234 42980 5236
rect 42924 5182 42926 5234
rect 42926 5182 42978 5234
rect 42978 5182 42980 5234
rect 42924 5180 42980 5182
rect 42476 5010 42532 5012
rect 42476 4958 42478 5010
rect 42478 4958 42530 5010
rect 42530 4958 42532 5010
rect 42476 4956 42532 4958
rect 42028 4508 42084 4564
rect 37324 4172 37380 4228
rect 37436 3836 37492 3892
rect 34972 3442 35028 3444
rect 34972 3390 34974 3442
rect 34974 3390 35026 3442
rect 35026 3390 35028 3442
rect 34972 3388 35028 3390
rect 33628 3276 33684 3332
rect 37884 4114 37940 4116
rect 37884 4062 37886 4114
rect 37886 4062 37938 4114
rect 37938 4062 37940 4114
rect 37884 4060 37940 4062
rect 39004 4114 39060 4116
rect 39004 4062 39006 4114
rect 39006 4062 39058 4114
rect 39058 4062 39060 4114
rect 39004 4060 39060 4062
rect 39340 4114 39396 4116
rect 39340 4062 39342 4114
rect 39342 4062 39394 4114
rect 39394 4062 39396 4114
rect 39340 4060 39396 4062
rect 41020 4060 41076 4116
rect 38780 3836 38836 3892
rect 39452 3666 39508 3668
rect 39452 3614 39454 3666
rect 39454 3614 39506 3666
rect 39506 3614 39508 3666
rect 39452 3612 39508 3614
rect 41916 4060 41972 4116
rect 41916 3836 41972 3892
rect 40348 3442 40404 3444
rect 40348 3390 40350 3442
rect 40350 3390 40402 3442
rect 40402 3390 40404 3442
rect 40348 3388 40404 3390
rect 41132 3442 41188 3444
rect 41132 3390 41134 3442
rect 41134 3390 41186 3442
rect 41186 3390 41188 3442
rect 41132 3388 41188 3390
rect 42140 4732 42196 4788
rect 44492 6188 44548 6244
rect 44044 6076 44100 6132
rect 43260 5794 43316 5796
rect 43260 5742 43262 5794
rect 43262 5742 43314 5794
rect 43314 5742 43316 5794
rect 43260 5740 43316 5742
rect 43820 5180 43876 5236
rect 43932 5852 43988 5908
rect 43148 4956 43204 5012
rect 42700 4844 42756 4900
rect 43148 4562 43204 4564
rect 43148 4510 43150 4562
rect 43150 4510 43202 4562
rect 43202 4510 43204 4562
rect 43148 4508 43204 4510
rect 44044 5740 44100 5796
rect 44156 5068 44212 5124
rect 44604 5906 44660 5908
rect 44604 5854 44606 5906
rect 44606 5854 44658 5906
rect 44658 5854 44660 5906
rect 44604 5852 44660 5854
rect 46508 9154 46564 9156
rect 46508 9102 46510 9154
rect 46510 9102 46562 9154
rect 46562 9102 46564 9154
rect 46508 9100 46564 9102
rect 46956 9100 47012 9156
rect 46620 8988 46676 9044
rect 49308 13074 49364 13076
rect 49308 13022 49310 13074
rect 49310 13022 49362 13074
rect 49362 13022 49364 13074
rect 49308 13020 49364 13022
rect 49644 12796 49700 12852
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 52332 13804 52388 13860
rect 51212 13074 51268 13076
rect 51212 13022 51214 13074
rect 51214 13022 51266 13074
rect 51266 13022 51268 13074
rect 51212 13020 51268 13022
rect 53900 16994 53956 16996
rect 53900 16942 53902 16994
rect 53902 16942 53954 16994
rect 53954 16942 53956 16994
rect 53900 16940 53956 16942
rect 53676 16828 53732 16884
rect 54012 16882 54068 16884
rect 54012 16830 54014 16882
rect 54014 16830 54066 16882
rect 54066 16830 54068 16882
rect 54012 16828 54068 16830
rect 55020 16828 55076 16884
rect 54460 15932 54516 15988
rect 53676 15874 53732 15876
rect 53676 15822 53678 15874
rect 53678 15822 53730 15874
rect 53730 15822 53732 15874
rect 53676 15820 53732 15822
rect 54236 15820 54292 15876
rect 53564 14812 53620 14868
rect 55244 15986 55300 15988
rect 55244 15934 55246 15986
rect 55246 15934 55298 15986
rect 55298 15934 55300 15986
rect 55244 15932 55300 15934
rect 54796 15314 54852 15316
rect 54796 15262 54798 15314
rect 54798 15262 54850 15314
rect 54850 15262 54852 15314
rect 54796 15260 54852 15262
rect 54684 14642 54740 14644
rect 54684 14590 54686 14642
rect 54686 14590 54738 14642
rect 54738 14590 54740 14642
rect 54684 14588 54740 14590
rect 55580 16882 55636 16884
rect 55580 16830 55582 16882
rect 55582 16830 55634 16882
rect 55634 16830 55636 16882
rect 55580 16828 55636 16830
rect 56028 16828 56084 16884
rect 56252 18396 56308 18452
rect 56476 20242 56532 20244
rect 56476 20190 56478 20242
rect 56478 20190 56530 20242
rect 56530 20190 56532 20242
rect 56476 20188 56532 20190
rect 56812 19964 56868 20020
rect 56700 18732 56756 18788
rect 56588 18620 56644 18676
rect 56476 18396 56532 18452
rect 57148 24668 57204 24724
rect 57260 25340 57316 25396
rect 57484 24946 57540 24948
rect 57484 24894 57486 24946
rect 57486 24894 57538 24946
rect 57538 24894 57540 24946
rect 57484 24892 57540 24894
rect 57820 24722 57876 24724
rect 57820 24670 57822 24722
rect 57822 24670 57874 24722
rect 57874 24670 57876 24722
rect 57820 24668 57876 24670
rect 58044 24610 58100 24612
rect 58044 24558 58046 24610
rect 58046 24558 58098 24610
rect 58098 24558 58100 24610
rect 58044 24556 58100 24558
rect 57260 21532 57316 21588
rect 57708 21586 57764 21588
rect 57708 21534 57710 21586
rect 57710 21534 57762 21586
rect 57762 21534 57764 21586
rect 57708 21532 57764 21534
rect 57596 21474 57652 21476
rect 57596 21422 57598 21474
rect 57598 21422 57650 21474
rect 57650 21422 57652 21474
rect 57596 21420 57652 21422
rect 57596 21196 57652 21252
rect 58156 22146 58212 22148
rect 58156 22094 58158 22146
rect 58158 22094 58210 22146
rect 58210 22094 58212 22146
rect 58156 22092 58212 22094
rect 58492 21586 58548 21588
rect 58492 21534 58494 21586
rect 58494 21534 58546 21586
rect 58546 21534 58548 21586
rect 58492 21532 58548 21534
rect 58044 20636 58100 20692
rect 57932 20076 57988 20132
rect 57820 20018 57876 20020
rect 57820 19966 57822 20018
rect 57822 19966 57874 20018
rect 57874 19966 57876 20018
rect 57820 19964 57876 19966
rect 57260 19740 57316 19796
rect 58380 20412 58436 20468
rect 58156 19852 58212 19908
rect 57372 18732 57428 18788
rect 56476 17052 56532 17108
rect 56364 16994 56420 16996
rect 56364 16942 56366 16994
rect 56366 16942 56418 16994
rect 56418 16942 56420 16994
rect 56364 16940 56420 16942
rect 57708 18732 57764 18788
rect 57596 18674 57652 18676
rect 57596 18622 57598 18674
rect 57598 18622 57650 18674
rect 57650 18622 57652 18674
rect 57596 18620 57652 18622
rect 57820 18562 57876 18564
rect 57820 18510 57822 18562
rect 57822 18510 57874 18562
rect 57874 18510 57876 18562
rect 57820 18508 57876 18510
rect 57036 16940 57092 16996
rect 57260 17276 57316 17332
rect 56812 16604 56868 16660
rect 55692 15932 55748 15988
rect 56364 15484 56420 15540
rect 55580 15314 55636 15316
rect 55580 15262 55582 15314
rect 55582 15262 55634 15314
rect 55634 15262 55636 15314
rect 55580 15260 55636 15262
rect 56700 15314 56756 15316
rect 56700 15262 56702 15314
rect 56702 15262 56754 15314
rect 56754 15262 56756 15314
rect 56700 15260 56756 15262
rect 56476 14642 56532 14644
rect 56476 14590 56478 14642
rect 56478 14590 56530 14642
rect 56530 14590 56532 14642
rect 56476 14588 56532 14590
rect 56588 13916 56644 13972
rect 53788 13858 53844 13860
rect 53788 13806 53790 13858
rect 53790 13806 53842 13858
rect 53842 13806 53844 13858
rect 53788 13804 53844 13806
rect 54796 13522 54852 13524
rect 54796 13470 54798 13522
rect 54798 13470 54850 13522
rect 54850 13470 54852 13522
rect 54796 13468 54852 13470
rect 55468 13468 55524 13524
rect 52108 13074 52164 13076
rect 52108 13022 52110 13074
rect 52110 13022 52162 13074
rect 52162 13022 52164 13074
rect 52108 13020 52164 13022
rect 50316 12908 50372 12964
rect 50988 12962 51044 12964
rect 50988 12910 50990 12962
rect 50990 12910 51042 12962
rect 51042 12910 51044 12962
rect 50988 12908 51044 12910
rect 50764 12850 50820 12852
rect 50764 12798 50766 12850
rect 50766 12798 50818 12850
rect 50818 12798 50820 12850
rect 50764 12796 50820 12798
rect 50204 12684 50260 12740
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 49756 12402 49812 12404
rect 49756 12350 49758 12402
rect 49758 12350 49810 12402
rect 49810 12350 49812 12402
rect 49756 12348 49812 12350
rect 49532 11116 49588 11172
rect 48748 10834 48804 10836
rect 48748 10782 48750 10834
rect 48750 10782 48802 10834
rect 48802 10782 48804 10834
rect 48748 10780 48804 10782
rect 49196 10780 49252 10836
rect 48524 10108 48580 10164
rect 48300 9938 48356 9940
rect 48300 9886 48302 9938
rect 48302 9886 48354 9938
rect 48354 9886 48356 9938
rect 48300 9884 48356 9886
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 49756 10834 49812 10836
rect 49756 10782 49758 10834
rect 49758 10782 49810 10834
rect 49810 10782 49812 10834
rect 49756 10780 49812 10782
rect 49196 9884 49252 9940
rect 51324 12684 51380 12740
rect 51660 11282 51716 11284
rect 51660 11230 51662 11282
rect 51662 11230 51714 11282
rect 51714 11230 51716 11282
rect 51660 11228 51716 11230
rect 53116 11228 53172 11284
rect 53676 11228 53732 11284
rect 49868 10386 49924 10388
rect 49868 10334 49870 10386
rect 49870 10334 49922 10386
rect 49922 10334 49924 10386
rect 49868 10332 49924 10334
rect 49532 10108 49588 10164
rect 47404 9154 47460 9156
rect 47404 9102 47406 9154
rect 47406 9102 47458 9154
rect 47458 9102 47460 9154
rect 47404 9100 47460 9102
rect 47180 9042 47236 9044
rect 47180 8990 47182 9042
rect 47182 8990 47234 9042
rect 47234 8990 47236 9042
rect 47628 9154 47684 9156
rect 47628 9102 47630 9154
rect 47630 9102 47682 9154
rect 47682 9102 47684 9154
rect 47628 9100 47684 9102
rect 49084 9100 49140 9156
rect 47180 8988 47236 8990
rect 47068 8370 47124 8372
rect 47068 8318 47070 8370
rect 47070 8318 47122 8370
rect 47122 8318 47124 8370
rect 47068 8316 47124 8318
rect 47740 8316 47796 8372
rect 53340 10444 53396 10500
rect 51660 10332 51716 10388
rect 51548 9772 51604 9828
rect 52108 9772 52164 9828
rect 49868 9714 49924 9716
rect 49868 9662 49870 9714
rect 49870 9662 49922 9714
rect 49922 9662 49924 9714
rect 49868 9660 49924 9662
rect 50428 9660 50484 9716
rect 49756 9154 49812 9156
rect 49756 9102 49758 9154
rect 49758 9102 49810 9154
rect 49810 9102 49812 9154
rect 49756 9100 49812 9102
rect 50876 9548 50932 9604
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 51548 9602 51604 9604
rect 51548 9550 51550 9602
rect 51550 9550 51602 9602
rect 51602 9550 51604 9602
rect 51548 9548 51604 9550
rect 50428 9154 50484 9156
rect 50428 9102 50430 9154
rect 50430 9102 50482 9154
rect 50482 9102 50484 9154
rect 50428 9100 50484 9102
rect 45276 6130 45332 6132
rect 45276 6078 45278 6130
rect 45278 6078 45330 6130
rect 45330 6078 45332 6130
rect 45276 6076 45332 6078
rect 45500 6018 45556 6020
rect 45500 5966 45502 6018
rect 45502 5966 45554 6018
rect 45554 5966 45556 6018
rect 45500 5964 45556 5966
rect 46284 6018 46340 6020
rect 46284 5966 46286 6018
rect 46286 5966 46338 6018
rect 46338 5966 46340 6018
rect 46284 5964 46340 5966
rect 47068 6018 47124 6020
rect 47068 5966 47070 6018
rect 47070 5966 47122 6018
rect 47122 5966 47124 6018
rect 47068 5964 47124 5966
rect 45388 5852 45444 5908
rect 46172 5906 46228 5908
rect 46172 5854 46174 5906
rect 46174 5854 46226 5906
rect 46226 5854 46228 5906
rect 46172 5852 46228 5854
rect 45836 5234 45892 5236
rect 45836 5182 45838 5234
rect 45838 5182 45890 5234
rect 45890 5182 45892 5234
rect 45836 5180 45892 5182
rect 44380 4732 44436 4788
rect 44492 4956 44548 5012
rect 44492 4508 44548 4564
rect 45724 4732 45780 4788
rect 45724 4562 45780 4564
rect 45724 4510 45726 4562
rect 45726 4510 45778 4562
rect 45778 4510 45780 4562
rect 45724 4508 45780 4510
rect 46956 5906 47012 5908
rect 46956 5854 46958 5906
rect 46958 5854 47010 5906
rect 47010 5854 47012 5906
rect 46956 5852 47012 5854
rect 49756 7980 49812 8036
rect 49644 7644 49700 7700
rect 48636 6412 48692 6468
rect 47964 6130 48020 6132
rect 47964 6078 47966 6130
rect 47966 6078 48018 6130
rect 48018 6078 48020 6130
rect 47964 6076 48020 6078
rect 46284 5682 46340 5684
rect 46284 5630 46286 5682
rect 46286 5630 46338 5682
rect 46338 5630 46340 5682
rect 46284 5628 46340 5630
rect 47292 5628 47348 5684
rect 48524 5292 48580 5348
rect 48076 5180 48132 5236
rect 44828 4396 44884 4452
rect 45612 4450 45668 4452
rect 45612 4398 45614 4450
rect 45614 4398 45666 4450
rect 45666 4398 45668 4450
rect 45612 4396 45668 4398
rect 48188 5068 48244 5124
rect 48748 6188 48804 6244
rect 48748 5292 48804 5348
rect 50652 9042 50708 9044
rect 50652 8990 50654 9042
rect 50654 8990 50706 9042
rect 50706 8990 50708 9042
rect 50652 8988 50708 8990
rect 51660 9154 51716 9156
rect 51660 9102 51662 9154
rect 51662 9102 51714 9154
rect 51714 9102 51716 9154
rect 51660 9100 51716 9102
rect 51548 9042 51604 9044
rect 51548 8990 51550 9042
rect 51550 8990 51602 9042
rect 51602 8990 51604 9042
rect 51548 8988 51604 8990
rect 51100 8764 51156 8820
rect 51884 8316 51940 8372
rect 50876 8204 50932 8260
rect 50652 7980 50708 8036
rect 50876 7980 50932 8036
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 52780 9772 52836 9828
rect 56028 12290 56084 12292
rect 56028 12238 56030 12290
rect 56030 12238 56082 12290
rect 56082 12238 56084 12290
rect 56028 12236 56084 12238
rect 55580 12178 55636 12180
rect 55580 12126 55582 12178
rect 55582 12126 55634 12178
rect 55634 12126 55636 12178
rect 55580 12124 55636 12126
rect 53900 10444 53956 10500
rect 55356 11676 55412 11732
rect 54684 11282 54740 11284
rect 54684 11230 54686 11282
rect 54686 11230 54738 11282
rect 54738 11230 54740 11282
rect 54684 11228 54740 11230
rect 54796 11116 54852 11172
rect 56028 11116 56084 11172
rect 56140 11788 56196 11844
rect 54572 10498 54628 10500
rect 54572 10446 54574 10498
rect 54574 10446 54626 10498
rect 54626 10446 54628 10498
rect 54572 10444 54628 10446
rect 54124 10332 54180 10388
rect 54460 10332 54516 10388
rect 54012 10220 54068 10276
rect 53676 9154 53732 9156
rect 53676 9102 53678 9154
rect 53678 9102 53730 9154
rect 53730 9102 53732 9154
rect 53676 9100 53732 9102
rect 54348 9100 54404 9156
rect 53564 8988 53620 9044
rect 53004 8764 53060 8820
rect 53228 8316 53284 8372
rect 52668 8258 52724 8260
rect 52668 8206 52670 8258
rect 52670 8206 52722 8258
rect 52722 8206 52724 8258
rect 52668 8204 52724 8206
rect 53116 8092 53172 8148
rect 53452 8316 53508 8372
rect 54236 9042 54292 9044
rect 54236 8990 54238 9042
rect 54238 8990 54290 9042
rect 54290 8990 54292 9042
rect 54236 8988 54292 8990
rect 53676 8146 53732 8148
rect 53676 8094 53678 8146
rect 53678 8094 53730 8146
rect 53730 8094 53732 8146
rect 53676 8092 53732 8094
rect 54796 10220 54852 10276
rect 54572 9548 54628 9604
rect 54684 9266 54740 9268
rect 54684 9214 54686 9266
rect 54686 9214 54738 9266
rect 54738 9214 54740 9266
rect 54684 9212 54740 9214
rect 55132 10108 55188 10164
rect 55468 10050 55524 10052
rect 55468 9998 55470 10050
rect 55470 9998 55522 10050
rect 55522 9998 55524 10050
rect 55468 9996 55524 9998
rect 55692 9212 55748 9268
rect 55356 9100 55412 9156
rect 54684 8258 54740 8260
rect 54684 8206 54686 8258
rect 54686 8206 54738 8258
rect 54738 8206 54740 8258
rect 54684 8204 54740 8206
rect 55804 9996 55860 10052
rect 56028 9772 56084 9828
rect 57260 15372 57316 15428
rect 57596 16658 57652 16660
rect 57596 16606 57598 16658
rect 57598 16606 57650 16658
rect 57650 16606 57652 16658
rect 57596 16604 57652 16606
rect 58604 18732 58660 18788
rect 58716 28700 58772 28756
rect 58380 17052 58436 17108
rect 57596 15314 57652 15316
rect 57596 15262 57598 15314
rect 57598 15262 57650 15314
rect 57650 15262 57652 15314
rect 57596 15260 57652 15262
rect 56924 12236 56980 12292
rect 56252 11228 56308 11284
rect 56588 11282 56644 11284
rect 56588 11230 56590 11282
rect 56590 11230 56642 11282
rect 56642 11230 56644 11282
rect 56588 11228 56644 11230
rect 56364 11170 56420 11172
rect 56364 11118 56366 11170
rect 56366 11118 56418 11170
rect 56418 11118 56420 11170
rect 56364 11116 56420 11118
rect 56364 10220 56420 10276
rect 57932 15372 57988 15428
rect 57820 13916 57876 13972
rect 58716 15484 58772 15540
rect 57596 12290 57652 12292
rect 57596 12238 57598 12290
rect 57598 12238 57650 12290
rect 57650 12238 57652 12290
rect 57596 12236 57652 12238
rect 57708 12178 57764 12180
rect 57708 12126 57710 12178
rect 57710 12126 57762 12178
rect 57762 12126 57764 12178
rect 57708 12124 57764 12126
rect 57148 11900 57204 11956
rect 55916 9100 55972 9156
rect 56924 9996 56980 10052
rect 58492 11900 58548 11956
rect 57708 11116 57764 11172
rect 58044 9772 58100 9828
rect 53788 6524 53844 6580
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 57708 7644 57764 7700
rect 56700 6524 56756 6580
rect 55020 6466 55076 6468
rect 55020 6414 55022 6466
rect 55022 6414 55074 6466
rect 55074 6414 55076 6466
rect 55020 6412 55076 6414
rect 55468 6466 55524 6468
rect 55468 6414 55470 6466
rect 55470 6414 55522 6466
rect 55522 6414 55524 6466
rect 55468 6412 55524 6414
rect 53788 6076 53844 6132
rect 49196 5234 49252 5236
rect 49196 5182 49198 5234
rect 49198 5182 49250 5234
rect 49250 5182 49252 5234
rect 49196 5180 49252 5182
rect 48972 5122 49028 5124
rect 48972 5070 48974 5122
rect 48974 5070 49026 5122
rect 49026 5070 49028 5122
rect 48972 5068 49028 5070
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 47516 3724 47572 3780
rect 42028 3388 42084 3444
rect 48076 3388 48132 3444
rect 48748 3442 48804 3444
rect 48748 3390 48750 3442
rect 48750 3390 48802 3442
rect 48802 3390 48804 3442
rect 48748 3388 48804 3390
rect 56028 3388 56084 3444
rect 55356 3330 55412 3332
rect 55356 3278 55358 3330
rect 55358 3278 55410 3330
rect 55410 3278 55412 3330
rect 55356 3276 55412 3278
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
rect 56588 3442 56644 3444
rect 56588 3390 56590 3442
rect 56590 3390 56642 3442
rect 56642 3390 56644 3442
rect 56588 3388 56644 3390
<< metal3 >>
rect 3714 60844 3724 60900
rect 3780 60844 25340 60900
rect 25396 60844 25406 60900
rect 1362 60732 1372 60788
rect 1428 60732 13692 60788
rect 13748 60732 13758 60788
rect 1698 60620 1708 60676
rect 1764 60620 16492 60676
rect 16548 60620 16558 60676
rect 4466 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4750 60396
rect 35186 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35470 60396
rect 30146 60060 30156 60116
rect 30212 60060 31052 60116
rect 31108 60060 31118 60116
rect 50194 60060 50204 60116
rect 50260 60060 51100 60116
rect 51156 60060 51166 60116
rect 4610 59948 4620 60004
rect 4676 59948 4956 60004
rect 5012 59948 9772 60004
rect 9828 59948 14924 60004
rect 14980 59948 14990 60004
rect 5058 59836 5068 59892
rect 5124 59836 5852 59892
rect 5908 59836 5918 59892
rect 6290 59836 6300 59892
rect 6356 59836 7644 59892
rect 7700 59836 7710 59892
rect 14354 59836 14364 59892
rect 14420 59836 14700 59892
rect 14756 59836 14766 59892
rect 3714 59724 3724 59780
rect 3780 59724 10668 59780
rect 10724 59724 10734 59780
rect 11778 59724 11788 59780
rect 11844 59724 12348 59780
rect 12404 59724 12414 59780
rect 14914 59724 14924 59780
rect 14980 59724 15932 59780
rect 15988 59724 15998 59780
rect 24658 59724 24668 59780
rect 24724 59724 29820 59780
rect 29876 59724 30380 59780
rect 30436 59724 30446 59780
rect 35522 59724 35532 59780
rect 35588 59724 36316 59780
rect 36372 59724 36988 59780
rect 37044 59724 37054 59780
rect 39666 59724 39676 59780
rect 39732 59724 49868 59780
rect 49924 59724 50428 59780
rect 50484 59724 50494 59780
rect 8978 59612 8988 59668
rect 9044 59612 10108 59668
rect 10164 59612 12460 59668
rect 12516 59612 12526 59668
rect 13458 59612 13468 59668
rect 13524 59612 15708 59668
rect 15764 59612 15774 59668
rect 23314 59612 23324 59668
rect 23380 59612 24108 59668
rect 24164 59612 25228 59668
rect 25284 59612 25676 59668
rect 25732 59612 33740 59668
rect 33796 59612 33806 59668
rect 19826 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20110 59612
rect 50546 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50830 59612
rect 9874 59500 9884 59556
rect 9940 59500 11844 59556
rect 12786 59500 12796 59556
rect 12852 59500 17612 59556
rect 17668 59500 18060 59556
rect 18116 59500 18508 59556
rect 18564 59500 18574 59556
rect 23538 59500 23548 59556
rect 23604 59500 24556 59556
rect 24612 59500 24892 59556
rect 24948 59500 40796 59556
rect 40852 59500 40862 59556
rect 11788 59444 11844 59500
rect 4610 59388 4620 59444
rect 4676 59388 5740 59444
rect 5796 59388 6748 59444
rect 6804 59388 6814 59444
rect 8082 59388 8092 59444
rect 8148 59388 11564 59444
rect 11620 59388 11630 59444
rect 11788 59388 14700 59444
rect 14756 59388 14766 59444
rect 14914 59388 14924 59444
rect 14980 59388 17948 59444
rect 18004 59388 18014 59444
rect 5058 59276 5068 59332
rect 5124 59276 6412 59332
rect 6468 59276 8652 59332
rect 8708 59276 9772 59332
rect 9828 59276 9838 59332
rect 10658 59276 10668 59332
rect 10724 59276 18396 59332
rect 18452 59276 18462 59332
rect 19506 59276 19516 59332
rect 19572 59276 20076 59332
rect 20132 59276 26684 59332
rect 26740 59276 26908 59332
rect 26964 59276 26974 59332
rect 30146 59276 30156 59332
rect 30212 59276 30716 59332
rect 30772 59276 30782 59332
rect 38210 59276 38220 59332
rect 38276 59276 39340 59332
rect 39396 59276 40572 59332
rect 40628 59276 40638 59332
rect 42018 59276 42028 59332
rect 42084 59276 45500 59332
rect 45556 59276 45566 59332
rect 5842 59164 5852 59220
rect 5908 59164 7196 59220
rect 7252 59164 11004 59220
rect 11060 59164 11070 59220
rect 13010 59164 13020 59220
rect 13076 59164 14364 59220
rect 14420 59164 14430 59220
rect 22978 59164 22988 59220
rect 23044 59164 23884 59220
rect 23940 59164 28028 59220
rect 28084 59164 28094 59220
rect 28690 59164 28700 59220
rect 28756 59164 30828 59220
rect 30884 59164 30894 59220
rect 32834 59164 32844 59220
rect 32900 59164 33964 59220
rect 34020 59164 34524 59220
rect 34580 59164 34590 59220
rect 34748 59164 41468 59220
rect 41524 59164 42364 59220
rect 42420 59164 42430 59220
rect 44930 59164 44940 59220
rect 44996 59164 45388 59220
rect 45444 59164 45454 59220
rect 34748 59108 34804 59164
rect 4834 59052 4844 59108
rect 4900 59052 5964 59108
rect 6020 59052 6030 59108
rect 7634 59052 7644 59108
rect 7700 59052 9324 59108
rect 9380 59052 9390 59108
rect 10770 59052 10780 59108
rect 10836 59052 12348 59108
rect 12404 59052 12414 59108
rect 13234 59052 13244 59108
rect 13300 59052 13916 59108
rect 13972 59052 13982 59108
rect 16034 59052 16044 59108
rect 16100 59052 18620 59108
rect 18676 59052 20076 59108
rect 20132 59052 20142 59108
rect 33842 59052 33852 59108
rect 33908 59052 34804 59108
rect 36754 59052 36764 59108
rect 36820 59052 38108 59108
rect 38164 59052 39284 59108
rect 39228 58996 39284 59052
rect 2706 58940 2716 58996
rect 2772 58940 3612 58996
rect 3668 58940 4060 58996
rect 4116 58940 5852 58996
rect 5908 58940 5918 58996
rect 12114 58940 12124 58996
rect 12180 58940 13468 58996
rect 13524 58940 13534 58996
rect 14690 58940 14700 58996
rect 14756 58940 16604 58996
rect 16660 58940 16670 58996
rect 29922 58940 29932 58996
rect 29988 58940 30716 58996
rect 30772 58940 30782 58996
rect 32834 58940 32844 58996
rect 32900 58940 34076 58996
rect 34132 58940 34142 58996
rect 34738 58940 34748 58996
rect 34804 58940 35420 58996
rect 35476 58940 38668 58996
rect 39218 58940 39228 58996
rect 39284 58940 40348 58996
rect 40404 58940 41804 58996
rect 41860 58940 41870 58996
rect 38612 58884 38668 58940
rect 12898 58828 12908 58884
rect 12964 58828 12974 58884
rect 14018 58828 14028 58884
rect 14084 58828 15764 58884
rect 15922 58828 15932 58884
rect 15988 58828 16492 58884
rect 16548 58828 16558 58884
rect 21858 58828 21868 58884
rect 21924 58828 27692 58884
rect 27748 58828 27758 58884
rect 38612 58828 40572 58884
rect 40628 58828 42476 58884
rect 42532 58828 42542 58884
rect 4466 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4750 58828
rect 12908 58772 12964 58828
rect 15708 58772 15764 58828
rect 35186 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35470 58828
rect 6290 58716 6300 58772
rect 6356 58716 8092 58772
rect 8148 58716 11788 58772
rect 11844 58716 11854 58772
rect 12908 58716 13468 58772
rect 13524 58716 13534 58772
rect 15708 58716 16940 58772
rect 16996 58716 17006 58772
rect 21746 58716 21756 58772
rect 21812 58716 22316 58772
rect 22372 58716 23548 58772
rect 23604 58716 23614 58772
rect 27234 58716 27244 58772
rect 27300 58716 28364 58772
rect 28420 58716 28430 58772
rect 30034 58716 30044 58772
rect 30100 58716 31276 58772
rect 31332 58716 31342 58772
rect 35634 58716 35644 58772
rect 35700 58716 38668 58772
rect 41570 58716 41580 58772
rect 41636 58716 43708 58772
rect 43764 58716 43774 58772
rect 38612 58660 38668 58716
rect 18162 58604 18172 58660
rect 18228 58604 22092 58660
rect 22148 58604 22764 58660
rect 22820 58604 22830 58660
rect 24556 58604 26908 58660
rect 26964 58604 26974 58660
rect 28578 58604 28588 58660
rect 28644 58604 29820 58660
rect 29876 58604 30156 58660
rect 30212 58604 30604 58660
rect 30660 58604 30670 58660
rect 34962 58604 34972 58660
rect 35028 58604 37660 58660
rect 37716 58604 37726 58660
rect 38612 58604 39116 58660
rect 39172 58604 41244 58660
rect 41300 58604 44492 58660
rect 44548 58604 44558 58660
rect 24556 58548 24612 58604
rect 16594 58492 16604 58548
rect 16660 58492 18116 58548
rect 20290 58492 20300 58548
rect 20356 58492 24556 58548
rect 24612 58492 24622 58548
rect 26786 58492 26796 58548
rect 26852 58492 27356 58548
rect 27412 58492 27422 58548
rect 28130 58492 28140 58548
rect 28196 58492 32732 58548
rect 32788 58492 32956 58548
rect 33012 58492 33022 58548
rect 40786 58492 40796 58548
rect 40852 58492 42812 58548
rect 42868 58492 42878 58548
rect 43138 58492 43148 58548
rect 43204 58492 43596 58548
rect 43652 58492 45052 58548
rect 45108 58492 45118 58548
rect 46386 58492 46396 58548
rect 46452 58492 46732 58548
rect 46788 58492 47180 58548
rect 47236 58492 47246 58548
rect 18060 58436 18116 58492
rect 12674 58380 12684 58436
rect 12740 58380 13804 58436
rect 13860 58380 13870 58436
rect 16258 58380 16268 58436
rect 16324 58380 17500 58436
rect 17556 58380 17566 58436
rect 18050 58380 18060 58436
rect 18116 58380 20188 58436
rect 20244 58380 20254 58436
rect 24770 58380 24780 58436
rect 24836 58380 25900 58436
rect 25956 58380 26460 58436
rect 26516 58380 26526 58436
rect 30482 58380 30492 58436
rect 30548 58380 32508 58436
rect 32564 58380 33180 58436
rect 33236 58380 33246 58436
rect 33506 58380 33516 58436
rect 33572 58380 33740 58436
rect 33796 58380 34412 58436
rect 34468 58380 35084 58436
rect 35140 58380 35150 58436
rect 36642 58380 36652 58436
rect 36708 58380 37548 58436
rect 37604 58380 37614 58436
rect 38612 58380 38892 58436
rect 38948 58380 39452 58436
rect 39508 58380 40348 58436
rect 40404 58380 40414 58436
rect 46610 58380 46620 58436
rect 46676 58380 47516 58436
rect 47572 58380 50092 58436
rect 50148 58380 50158 58436
rect 38612 58324 38668 58380
rect 2482 58268 2492 58324
rect 2548 58268 7308 58324
rect 7364 58268 9100 58324
rect 9156 58268 9166 58324
rect 9426 58268 9436 58324
rect 9492 58268 9884 58324
rect 9940 58268 9950 58324
rect 14690 58268 14700 58324
rect 14756 58268 15484 58324
rect 15540 58268 18956 58324
rect 19012 58268 19180 58324
rect 19236 58268 19246 58324
rect 19842 58268 19852 58324
rect 19908 58268 24444 58324
rect 24500 58268 25452 58324
rect 25508 58268 25518 58324
rect 26338 58268 26348 58324
rect 26404 58268 27468 58324
rect 27524 58268 27804 58324
rect 27860 58268 28812 58324
rect 28868 58268 29148 58324
rect 29204 58268 29214 58324
rect 32274 58268 32284 58324
rect 32340 58268 33628 58324
rect 33684 58268 33694 58324
rect 37650 58268 37660 58324
rect 37716 58268 38668 58324
rect 40226 58268 40236 58324
rect 40292 58268 44492 58324
rect 44548 58268 44558 58324
rect 3378 58156 3388 58212
rect 3444 58156 3482 58212
rect 5954 58156 5964 58212
rect 6020 58156 6748 58212
rect 6804 58156 11676 58212
rect 11732 58156 11742 58212
rect 12786 58156 12796 58212
rect 12852 58156 14028 58212
rect 14084 58156 14094 58212
rect 20962 58156 20972 58212
rect 21028 58156 21868 58212
rect 21924 58156 21934 58212
rect 29474 58156 29484 58212
rect 29540 58156 30716 58212
rect 30772 58156 31948 58212
rect 32050 58156 32060 58212
rect 32116 58156 32396 58212
rect 32452 58156 34860 58212
rect 34916 58156 34926 58212
rect 38098 58156 38108 58212
rect 38164 58156 38780 58212
rect 38836 58156 38846 58212
rect 43026 58156 43036 58212
rect 43092 58156 43484 58212
rect 43540 58156 47292 58212
rect 47348 58156 47358 58212
rect 31892 58100 31948 58156
rect 8978 58044 8988 58100
rect 9044 58044 10780 58100
rect 10836 58044 10846 58100
rect 31892 58044 36092 58100
rect 36148 58044 36158 58100
rect 19826 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20110 58044
rect 50546 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50830 58044
rect 4498 57932 4508 57988
rect 4564 57932 11900 57988
rect 11956 57932 11966 57988
rect 27122 57932 27132 57988
rect 27188 57932 27916 57988
rect 27972 57932 28588 57988
rect 28644 57932 28654 57988
rect 44370 57932 44380 57988
rect 44436 57932 44604 57988
rect 44660 57932 46060 57988
rect 46116 57932 46126 57988
rect 4050 57820 4060 57876
rect 4116 57820 4172 57876
rect 4228 57820 4956 57876
rect 5012 57820 5022 57876
rect 8754 57820 8764 57876
rect 8820 57820 14924 57876
rect 14980 57820 14990 57876
rect 38882 57820 38892 57876
rect 38948 57820 43260 57876
rect 43316 57820 43326 57876
rect 43474 57820 43484 57876
rect 43540 57820 44268 57876
rect 44324 57820 44334 57876
rect 45378 57820 45388 57876
rect 45444 57820 53788 57876
rect 53844 57820 53854 57876
rect 2930 57708 2940 57764
rect 2996 57708 4956 57764
rect 5012 57708 8652 57764
rect 8708 57708 11340 57764
rect 11396 57708 15260 57764
rect 15316 57708 15326 57764
rect 22502 57708 22540 57764
rect 22596 57708 22606 57764
rect 30034 57708 30044 57764
rect 30100 57708 35756 57764
rect 35812 57708 36316 57764
rect 36372 57708 36988 57764
rect 37044 57708 37054 57764
rect 3154 57596 3164 57652
rect 3220 57596 9996 57652
rect 10052 57596 10062 57652
rect 10434 57596 10444 57652
rect 10500 57596 13468 57652
rect 13524 57596 13534 57652
rect 19282 57596 19292 57652
rect 19348 57596 19852 57652
rect 19908 57596 19918 57652
rect 28690 57596 28700 57652
rect 28756 57596 31164 57652
rect 31220 57596 32172 57652
rect 32228 57596 32238 57652
rect 34290 57596 34300 57652
rect 34356 57596 34748 57652
rect 34804 57596 35644 57652
rect 35700 57596 35710 57652
rect 38770 57596 38780 57652
rect 38836 57596 39452 57652
rect 39508 57596 39518 57652
rect 46946 57596 46956 57652
rect 47012 57596 47740 57652
rect 47796 57596 48412 57652
rect 48468 57596 48478 57652
rect 51874 57596 51884 57652
rect 51940 57596 52220 57652
rect 52276 57596 52286 57652
rect 3714 57484 3724 57540
rect 3780 57484 4620 57540
rect 4676 57484 4686 57540
rect 5030 57484 5068 57540
rect 5124 57484 5134 57540
rect 6850 57484 6860 57540
rect 6916 57484 8428 57540
rect 8484 57484 8494 57540
rect 12786 57484 12796 57540
rect 12852 57484 13692 57540
rect 13748 57484 14364 57540
rect 14420 57484 14430 57540
rect 14914 57484 14924 57540
rect 14980 57484 15372 57540
rect 15428 57484 17052 57540
rect 17108 57484 17612 57540
rect 17668 57484 18172 57540
rect 18228 57484 18238 57540
rect 23426 57484 23436 57540
rect 23492 57484 23772 57540
rect 23828 57484 24108 57540
rect 24164 57484 24780 57540
rect 24836 57484 25564 57540
rect 25620 57484 25630 57540
rect 31714 57484 31724 57540
rect 31780 57484 32508 57540
rect 32564 57484 32574 57540
rect 40674 57484 40684 57540
rect 40740 57484 43372 57540
rect 43428 57484 43438 57540
rect 49970 57484 49980 57540
rect 50036 57484 50540 57540
rect 50596 57484 51996 57540
rect 52052 57484 52062 57540
rect 2380 57372 4508 57428
rect 4564 57372 4574 57428
rect 8530 57372 8540 57428
rect 8596 57372 9436 57428
rect 9492 57372 9502 57428
rect 11554 57372 11564 57428
rect 11620 57372 13132 57428
rect 13188 57372 13198 57428
rect 36530 57372 36540 57428
rect 36596 57372 37548 57428
rect 37604 57372 37614 57428
rect 47058 57372 47068 57428
rect 47124 57372 47516 57428
rect 47572 57372 48300 57428
rect 48356 57372 51548 57428
rect 51604 57372 51614 57428
rect 2380 57316 2436 57372
rect 2370 57260 2380 57316
rect 2436 57260 2446 57316
rect 8194 57260 8204 57316
rect 8260 57260 10332 57316
rect 10388 57260 10398 57316
rect 11666 57260 11676 57316
rect 11732 57260 13692 57316
rect 13748 57260 13758 57316
rect 19366 57260 19404 57316
rect 19460 57260 19470 57316
rect 19618 57260 19628 57316
rect 19684 57260 27916 57316
rect 27972 57260 27982 57316
rect 38658 57260 38668 57316
rect 38724 57260 42588 57316
rect 42644 57260 42654 57316
rect 4466 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4750 57260
rect 35186 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35470 57260
rect 10546 57148 10556 57204
rect 10612 57148 12124 57204
rect 12180 57148 12348 57204
rect 12404 57148 12414 57204
rect 20514 57148 20524 57204
rect 20580 57148 26348 57204
rect 26404 57148 26414 57204
rect 36530 57148 36540 57204
rect 36596 57148 38108 57204
rect 38164 57148 38174 57204
rect 8194 57036 8204 57092
rect 8260 57036 12012 57092
rect 12068 57036 13580 57092
rect 13636 57036 13646 57092
rect 16482 57036 16492 57092
rect 16548 57036 17724 57092
rect 17780 57036 17790 57092
rect 18610 57036 18620 57092
rect 18676 57036 19404 57092
rect 19460 57036 20188 57092
rect 20244 57036 20254 57092
rect 22754 57036 22764 57092
rect 22820 57036 23660 57092
rect 23716 57036 23996 57092
rect 24052 57036 24062 57092
rect 24780 57036 26124 57092
rect 26180 57036 26572 57092
rect 26628 57036 26638 57092
rect 34962 57036 34972 57092
rect 35028 57036 35868 57092
rect 35924 57036 35934 57092
rect 36306 57036 36316 57092
rect 36372 57036 37436 57092
rect 37492 57036 38220 57092
rect 38276 57036 38286 57092
rect 38434 57036 38444 57092
rect 38500 57036 43820 57092
rect 43876 57036 44156 57092
rect 44212 57036 44222 57092
rect 45490 57036 45500 57092
rect 45556 57036 45948 57092
rect 46004 57036 51996 57092
rect 52052 57036 52062 57092
rect 24780 56980 24836 57036
rect 1138 56924 1148 56980
rect 1204 56924 9156 56980
rect 5180 56812 8092 56868
rect 8148 56812 8158 56868
rect 5180 56644 5236 56812
rect 9100 56756 9156 56924
rect 14140 56924 14812 56980
rect 14868 56924 14878 56980
rect 15474 56924 15484 56980
rect 15540 56924 19180 56980
rect 19236 56924 19246 56980
rect 22082 56924 22092 56980
rect 22148 56924 22540 56980
rect 22596 56924 24108 56980
rect 24164 56924 24836 56980
rect 24994 56924 25004 56980
rect 25060 56924 25788 56980
rect 25844 56924 31500 56980
rect 31556 56924 31566 56980
rect 37762 56924 37772 56980
rect 37828 56924 38556 56980
rect 38612 56924 38622 56980
rect 51650 56924 51660 56980
rect 51716 56924 52332 56980
rect 52388 56924 52398 56980
rect 14140 56868 14196 56924
rect 11106 56812 11116 56868
rect 11172 56812 14140 56868
rect 14196 56812 14206 56868
rect 14354 56812 14364 56868
rect 14420 56812 16044 56868
rect 16100 56812 17500 56868
rect 17556 56812 17566 56868
rect 18386 56812 18396 56868
rect 18452 56812 22596 56868
rect 23762 56812 23772 56868
rect 23828 56812 25116 56868
rect 25172 56812 25182 56868
rect 28802 56812 28812 56868
rect 28868 56812 30492 56868
rect 30548 56812 32284 56868
rect 32340 56812 32350 56868
rect 38322 56812 38332 56868
rect 38388 56812 38780 56868
rect 38836 56812 38846 56868
rect 39330 56812 39340 56868
rect 39396 56812 40348 56868
rect 40404 56812 40414 56868
rect 48178 56812 48188 56868
rect 48244 56812 50092 56868
rect 50148 56812 50158 56868
rect 52098 56812 52108 56868
rect 52164 56812 52174 56868
rect 22540 56756 22596 56812
rect 52108 56756 52164 56812
rect 5842 56700 5852 56756
rect 5908 56700 6748 56756
rect 6804 56700 7644 56756
rect 7700 56700 8764 56756
rect 8820 56700 8830 56756
rect 9100 56700 15148 56756
rect 16482 56700 16492 56756
rect 16548 56700 16828 56756
rect 16884 56700 17276 56756
rect 17332 56700 17342 56756
rect 18050 56700 18060 56756
rect 18116 56700 22316 56756
rect 22372 56700 22382 56756
rect 22540 56700 25676 56756
rect 25732 56700 25742 56756
rect 28018 56700 28028 56756
rect 28084 56700 28588 56756
rect 28644 56700 30044 56756
rect 30100 56700 30110 56756
rect 31490 56700 31500 56756
rect 31556 56700 32172 56756
rect 32228 56700 32238 56756
rect 36418 56700 36428 56756
rect 36484 56700 38556 56756
rect 38612 56700 39116 56756
rect 39172 56700 39182 56756
rect 52108 56700 52332 56756
rect 52388 56700 53900 56756
rect 53956 56700 53966 56756
rect 2594 56588 2604 56644
rect 2660 56588 3500 56644
rect 3556 56588 3566 56644
rect 4274 56588 4284 56644
rect 4340 56588 5180 56644
rect 5236 56588 5246 56644
rect 6402 56588 6412 56644
rect 6468 56588 6524 56644
rect 6580 56588 6590 56644
rect 6850 56588 6860 56644
rect 6916 56588 7420 56644
rect 7476 56588 7486 56644
rect 8082 56588 8092 56644
rect 8148 56588 11564 56644
rect 11620 56588 11630 56644
rect 13570 56588 13580 56644
rect 13636 56588 14588 56644
rect 14644 56588 14654 56644
rect 7858 56476 7868 56532
rect 7924 56476 11228 56532
rect 11284 56476 11294 56532
rect 13010 56476 13020 56532
rect 13076 56476 13468 56532
rect 13524 56476 13534 56532
rect 8530 56364 8540 56420
rect 8596 56364 8876 56420
rect 8932 56364 13244 56420
rect 13300 56364 13310 56420
rect 2146 56252 2156 56308
rect 2212 56252 2716 56308
rect 2772 56252 2782 56308
rect 2930 56252 2940 56308
rect 2996 56252 5404 56308
rect 5460 56252 5470 56308
rect 6850 56252 6860 56308
rect 6916 56252 8988 56308
rect 9044 56252 9054 56308
rect 11106 56252 11116 56308
rect 11172 56252 12908 56308
rect 12964 56252 12974 56308
rect 2716 56196 2772 56252
rect 15092 56196 15148 56700
rect 19842 56588 19852 56644
rect 19908 56588 20972 56644
rect 21028 56588 21038 56644
rect 25218 56588 25228 56644
rect 25284 56588 31052 56644
rect 31108 56588 31118 56644
rect 37202 56588 37212 56644
rect 37268 56588 40236 56644
rect 40292 56588 41020 56644
rect 41076 56588 41086 56644
rect 46498 56588 46508 56644
rect 46564 56588 47740 56644
rect 47796 56588 47806 56644
rect 52210 56588 52220 56644
rect 52276 56588 52892 56644
rect 52948 56588 53564 56644
rect 53620 56588 53630 56644
rect 27010 56476 27020 56532
rect 27076 56476 29260 56532
rect 29316 56476 29326 56532
rect 31378 56476 31388 56532
rect 31444 56476 39004 56532
rect 39060 56476 39070 56532
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 22530 56364 22540 56420
rect 22596 56364 23324 56420
rect 23380 56364 23390 56420
rect 24098 56364 24108 56420
rect 24164 56364 38220 56420
rect 38276 56364 39788 56420
rect 39844 56364 39854 56420
rect 15922 56252 15932 56308
rect 15988 56252 17836 56308
rect 17892 56252 17902 56308
rect 23202 56252 23212 56308
rect 23268 56252 23660 56308
rect 23716 56252 23726 56308
rect 35522 56252 35532 56308
rect 35588 56252 35868 56308
rect 35924 56252 36316 56308
rect 36372 56252 36382 56308
rect 42802 56252 42812 56308
rect 42868 56252 43932 56308
rect 43988 56252 43998 56308
rect 50194 56252 50204 56308
rect 50260 56252 51436 56308
rect 51492 56252 51502 56308
rect 2716 56140 9212 56196
rect 9268 56140 9996 56196
rect 10052 56140 10780 56196
rect 10836 56140 10846 56196
rect 11862 56140 11900 56196
rect 11956 56140 11966 56196
rect 12786 56140 12796 56196
rect 12852 56140 14252 56196
rect 14308 56140 14318 56196
rect 15092 56140 21980 56196
rect 22036 56140 22046 56196
rect 8540 56084 8596 56140
rect 4050 56028 4060 56084
rect 4116 56028 8092 56084
rect 8148 56028 8158 56084
rect 8530 56028 8540 56084
rect 8596 56028 8606 56084
rect 11330 56028 11340 56084
rect 11396 56028 12124 56084
rect 12180 56028 12190 56084
rect 21410 56028 21420 56084
rect 21476 56028 22092 56084
rect 22148 56028 22428 56084
rect 22484 56028 22494 56084
rect 44594 56028 44604 56084
rect 44660 56028 46508 56084
rect 46564 56028 46574 56084
rect 46722 56028 46732 56084
rect 46788 56028 47852 56084
rect 47908 56028 47918 56084
rect 50194 56028 50204 56084
rect 50260 56028 51324 56084
rect 51380 56028 52220 56084
rect 52276 56028 52286 56084
rect 46732 55972 46788 56028
rect 1474 55916 1484 55972
rect 1540 55916 3164 55972
rect 3220 55916 3230 55972
rect 4610 55916 4620 55972
rect 4676 55916 6636 55972
rect 6692 55916 6702 55972
rect 7270 55916 7308 55972
rect 7364 55916 7374 55972
rect 11778 55916 11788 55972
rect 11844 55916 14028 55972
rect 14084 55916 14094 55972
rect 17574 55916 17612 55972
rect 17668 55916 17678 55972
rect 21970 55916 21980 55972
rect 22036 55916 27356 55972
rect 27412 55916 27422 55972
rect 31266 55916 31276 55972
rect 31332 55916 31836 55972
rect 31892 55916 35084 55972
rect 35140 55916 36092 55972
rect 36148 55916 36158 55972
rect 38658 55916 38668 55972
rect 38724 55916 39228 55972
rect 39284 55916 39294 55972
rect 43362 55916 43372 55972
rect 43428 55916 44380 55972
rect 44436 55916 44446 55972
rect 44818 55916 44828 55972
rect 44884 55916 46788 55972
rect 48514 55916 48524 55972
rect 48580 55916 49532 55972
rect 49588 55916 49598 55972
rect 53890 55916 53900 55972
rect 53956 55916 54460 55972
rect 54516 55916 55132 55972
rect 55188 55916 55198 55972
rect 44380 55860 44436 55916
rect 2370 55804 2380 55860
rect 2436 55804 3388 55860
rect 3444 55804 4732 55860
rect 4788 55804 4798 55860
rect 5058 55804 5068 55860
rect 5124 55804 11452 55860
rect 11508 55804 11518 55860
rect 19506 55804 19516 55860
rect 19572 55804 20076 55860
rect 20132 55804 20142 55860
rect 23986 55804 23996 55860
rect 24052 55804 25004 55860
rect 25060 55804 25070 55860
rect 31378 55804 31388 55860
rect 31444 55804 32060 55860
rect 32116 55804 32620 55860
rect 32676 55804 32686 55860
rect 39554 55804 39564 55860
rect 39620 55804 44044 55860
rect 44100 55804 44110 55860
rect 44380 55804 46508 55860
rect 46564 55804 46574 55860
rect 52882 55804 52892 55860
rect 52948 55804 57148 55860
rect 57204 55804 57214 55860
rect 20178 55692 20188 55748
rect 20244 55692 21308 55748
rect 21364 55692 27020 55748
rect 27076 55692 27086 55748
rect 40338 55692 40348 55748
rect 40404 55692 47852 55748
rect 47908 55692 47918 55748
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 2370 55580 2380 55636
rect 2436 55580 3052 55636
rect 3108 55580 3118 55636
rect 3602 55580 3612 55636
rect 3668 55580 4060 55636
rect 4116 55580 4126 55636
rect 12674 55580 12684 55636
rect 12740 55580 12750 55636
rect 18386 55580 18396 55636
rect 18452 55580 18508 55636
rect 18564 55580 18574 55636
rect 23314 55580 23324 55636
rect 23380 55580 23884 55636
rect 23940 55580 23950 55636
rect 25442 55580 25452 55636
rect 25508 55580 28476 55636
rect 28532 55580 28542 55636
rect 2258 55468 2268 55524
rect 2324 55468 4844 55524
rect 4900 55468 5068 55524
rect 5124 55468 5134 55524
rect 7074 55468 7084 55524
rect 7140 55468 7980 55524
rect 8036 55468 8046 55524
rect 12684 55412 12740 55580
rect 17052 55468 18172 55524
rect 18228 55468 18238 55524
rect 23762 55468 23772 55524
rect 23828 55468 38556 55524
rect 38612 55468 38622 55524
rect 43250 55468 43260 55524
rect 43316 55468 46284 55524
rect 46340 55468 46350 55524
rect 1698 55356 1708 55412
rect 1764 55356 10668 55412
rect 10724 55356 10734 55412
rect 10994 55356 11004 55412
rect 11060 55356 12124 55412
rect 12180 55356 13356 55412
rect 13412 55356 13422 55412
rect 15138 55356 15148 55412
rect 15204 55356 16828 55412
rect 16884 55356 16894 55412
rect 17052 55300 17108 55468
rect 20626 55356 20636 55412
rect 20692 55356 25564 55412
rect 25620 55356 26236 55412
rect 26292 55356 26302 55412
rect 2594 55244 2604 55300
rect 2660 55244 2670 55300
rect 3154 55244 3164 55300
rect 3220 55244 4844 55300
rect 4900 55244 4910 55300
rect 7158 55244 7196 55300
rect 7252 55244 7262 55300
rect 8082 55244 8092 55300
rect 8148 55244 8764 55300
rect 8820 55244 8830 55300
rect 10098 55244 10108 55300
rect 10164 55244 10444 55300
rect 10500 55244 11508 55300
rect 12002 55244 12012 55300
rect 12068 55244 17108 55300
rect 18722 55244 18732 55300
rect 18788 55244 19180 55300
rect 19236 55244 19964 55300
rect 20020 55244 20030 55300
rect 21858 55244 21868 55300
rect 21924 55244 22540 55300
rect 22596 55244 24668 55300
rect 24724 55244 24734 55300
rect 26450 55244 26460 55300
rect 26516 55244 27132 55300
rect 27188 55244 27198 55300
rect 32162 55244 32172 55300
rect 32228 55244 32844 55300
rect 32900 55244 33404 55300
rect 33460 55244 33470 55300
rect 34290 55244 34300 55300
rect 34356 55244 35420 55300
rect 35476 55244 35644 55300
rect 35700 55244 35710 55300
rect 38098 55244 38108 55300
rect 38164 55244 39452 55300
rect 39508 55244 39518 55300
rect 39666 55244 39676 55300
rect 39732 55244 40460 55300
rect 40516 55244 40526 55300
rect 41570 55244 41580 55300
rect 41636 55244 42476 55300
rect 42532 55244 42542 55300
rect 47730 55244 47740 55300
rect 47796 55244 48300 55300
rect 48356 55244 51996 55300
rect 52052 55244 52062 55300
rect 2604 55188 2660 55244
rect 11452 55188 11508 55244
rect 2604 55132 2828 55188
rect 2884 55132 7532 55188
rect 7588 55132 7598 55188
rect 9090 55132 9100 55188
rect 9156 55132 9772 55188
rect 9828 55132 9996 55188
rect 10052 55132 11228 55188
rect 11284 55132 11294 55188
rect 11452 55132 12124 55188
rect 12180 55132 12190 55188
rect 13794 55132 13804 55188
rect 13860 55132 15820 55188
rect 15876 55132 16716 55188
rect 16772 55132 16782 55188
rect 19058 55132 19068 55188
rect 19124 55132 19740 55188
rect 19796 55132 27692 55188
rect 27748 55132 27758 55188
rect 36306 55132 36316 55188
rect 36372 55132 37884 55188
rect 37940 55132 38668 55188
rect 38724 55132 40684 55188
rect 40740 55132 40750 55188
rect 48066 55132 48076 55188
rect 48132 55132 48412 55188
rect 48468 55132 48478 55188
rect 2604 55020 3724 55076
rect 3780 55020 3948 55076
rect 4004 55020 4844 55076
rect 4900 55020 7196 55076
rect 7252 55020 7262 55076
rect 7858 55020 7868 55076
rect 7924 55020 8092 55076
rect 8148 55020 8158 55076
rect 8978 55020 8988 55076
rect 9044 55020 9660 55076
rect 9716 55020 10220 55076
rect 10276 55020 10286 55076
rect 15698 55020 15708 55076
rect 15764 55020 16604 55076
rect 16660 55020 16670 55076
rect 20962 55020 20972 55076
rect 21028 55020 21644 55076
rect 21700 55020 24220 55076
rect 24276 55020 24286 55076
rect 26002 55020 26012 55076
rect 26068 55020 26572 55076
rect 26628 55020 26638 55076
rect 28466 55020 28476 55076
rect 28532 55020 33180 55076
rect 33236 55020 33246 55076
rect 40450 55020 40460 55076
rect 40516 55020 43372 55076
rect 43428 55020 43438 55076
rect 54002 55020 54012 55076
rect 54068 55020 54460 55076
rect 54516 55020 55244 55076
rect 55300 55020 57036 55076
rect 57092 55020 57102 55076
rect 2604 54852 2660 55020
rect 3602 54908 3612 54964
rect 3668 54908 4172 54964
rect 4228 54908 4396 54964
rect 4452 54908 10108 54964
rect 10164 54908 10174 54964
rect 14578 54908 14588 54964
rect 14644 54908 17836 54964
rect 17892 54908 17948 54964
rect 18004 54908 18014 54964
rect 22194 54908 22204 54964
rect 22260 54908 22652 54964
rect 22708 54908 25452 54964
rect 25508 54908 25518 54964
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 2594 54796 2604 54852
rect 2660 54796 2670 54852
rect 7410 54796 7420 54852
rect 7476 54796 8092 54852
rect 8148 54796 8158 54852
rect 2706 54684 2716 54740
rect 2772 54684 6188 54740
rect 6244 54684 6254 54740
rect 9090 54684 9100 54740
rect 9156 54684 10332 54740
rect 10388 54684 10398 54740
rect 14130 54684 14140 54740
rect 14196 54684 19628 54740
rect 19684 54684 19694 54740
rect 20178 54684 20188 54740
rect 20244 54684 20748 54740
rect 20804 54684 22764 54740
rect 22820 54684 22830 54740
rect 24434 54684 24444 54740
rect 24500 54684 30940 54740
rect 30996 54684 31276 54740
rect 31332 54684 31342 54740
rect 38770 54684 38780 54740
rect 38836 54684 39788 54740
rect 39844 54684 41804 54740
rect 41860 54684 41870 54740
rect 47954 54684 47964 54740
rect 48020 54684 48412 54740
rect 48468 54684 48478 54740
rect 1810 54572 1820 54628
rect 1876 54572 6076 54628
rect 6132 54572 6142 54628
rect 6402 54572 6412 54628
rect 6468 54572 10108 54628
rect 10164 54572 10174 54628
rect 14018 54572 14028 54628
rect 14084 54572 14252 54628
rect 14308 54572 14318 54628
rect 19282 54572 19292 54628
rect 19348 54572 19516 54628
rect 19572 54572 19582 54628
rect 19954 54572 19964 54628
rect 20020 54572 20300 54628
rect 20356 54572 20366 54628
rect 41906 54572 41916 54628
rect 41972 54572 42588 54628
rect 42644 54572 42654 54628
rect 48514 54572 48524 54628
rect 48580 54572 48692 54628
rect 52434 54572 52444 54628
rect 52500 54572 53228 54628
rect 53284 54572 54348 54628
rect 54404 54572 54414 54628
rect 3332 54460 4396 54516
rect 4452 54460 4462 54516
rect 4946 54460 4956 54516
rect 5012 54460 11788 54516
rect 11844 54460 11854 54516
rect 13346 54460 13356 54516
rect 13412 54460 20188 54516
rect 20244 54460 20254 54516
rect 27234 54460 27244 54516
rect 27300 54460 28140 54516
rect 28196 54460 28206 54516
rect 29026 54460 29036 54516
rect 29092 54460 30156 54516
rect 30212 54460 30222 54516
rect 3266 54348 3276 54404
rect 3332 54348 3388 54460
rect 48636 54404 48692 54572
rect 51762 54460 51772 54516
rect 51828 54460 53004 54516
rect 53060 54460 53070 54516
rect 53666 54460 53676 54516
rect 53732 54460 54236 54516
rect 54292 54460 54302 54516
rect 3938 54348 3948 54404
rect 4004 54348 4172 54404
rect 4228 54348 5740 54404
rect 5796 54348 6300 54404
rect 6356 54348 6366 54404
rect 7298 54348 7308 54404
rect 7364 54348 9996 54404
rect 10052 54348 10062 54404
rect 10210 54348 10220 54404
rect 10276 54348 11340 54404
rect 11396 54348 11406 54404
rect 12012 54348 15148 54404
rect 22082 54348 22092 54404
rect 22148 54348 25004 54404
rect 25060 54348 25070 54404
rect 30818 54348 30828 54404
rect 30884 54348 32508 54404
rect 32564 54348 32574 54404
rect 48626 54348 48636 54404
rect 48692 54348 48702 54404
rect 12012 54292 12068 54348
rect 15092 54292 15148 54348
rect 9734 54236 9772 54292
rect 9828 54236 9838 54292
rect 10546 54236 10556 54292
rect 10612 54236 12068 54292
rect 12226 54236 12236 54292
rect 12292 54236 14588 54292
rect 14644 54236 14654 54292
rect 15092 54236 17724 54292
rect 17780 54236 17790 54292
rect 32610 54236 32620 54292
rect 32676 54236 33628 54292
rect 33684 54236 34076 54292
rect 34132 54236 34142 54292
rect 41682 54236 41692 54292
rect 41748 54236 43148 54292
rect 43204 54236 44044 54292
rect 44100 54236 44110 54292
rect 47506 54236 47516 54292
rect 47572 54236 48300 54292
rect 48356 54236 48366 54292
rect 5068 54124 6748 54180
rect 6804 54124 8540 54180
rect 8596 54124 9660 54180
rect 9716 54124 9726 54180
rect 14018 54124 14028 54180
rect 14084 54124 16380 54180
rect 16436 54124 16940 54180
rect 16996 54124 19404 54180
rect 19460 54124 21196 54180
rect 21252 54124 25564 54180
rect 25620 54124 25630 54180
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 5068 53956 5124 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 5282 54012 5292 54068
rect 5348 54012 6524 54068
rect 6580 54012 10444 54068
rect 10500 54012 10510 54068
rect 11106 54012 11116 54068
rect 11172 54012 12460 54068
rect 12516 54012 12526 54068
rect 13458 54012 13468 54068
rect 13524 54012 15596 54068
rect 15652 54012 32284 54068
rect 32340 54012 32350 54068
rect 16604 53956 16660 54012
rect 1922 53900 1932 53956
rect 1988 53900 3500 53956
rect 3556 53900 4508 53956
rect 4564 53900 5124 53956
rect 6402 53900 6412 53956
rect 6468 53900 12404 53956
rect 13234 53900 13244 53956
rect 13300 53900 14028 53956
rect 14084 53900 14094 53956
rect 15026 53900 15036 53956
rect 15092 53900 15820 53956
rect 15876 53900 15886 53956
rect 16594 53900 16604 53956
rect 16660 53900 16670 53956
rect 19506 53900 19516 53956
rect 19572 53900 20524 53956
rect 20580 53900 20590 53956
rect 23314 53900 23324 53956
rect 23380 53900 23660 53956
rect 23716 53900 23726 53956
rect 40338 53900 40348 53956
rect 40404 53900 41580 53956
rect 41636 53900 41646 53956
rect 48738 53900 48748 53956
rect 48804 53900 52108 53956
rect 52164 53900 53452 53956
rect 53508 53900 53518 53956
rect 2930 53788 2940 53844
rect 2996 53788 3276 53844
rect 3332 53788 3342 53844
rect 4274 53788 4284 53844
rect 4340 53788 9548 53844
rect 9604 53788 9614 53844
rect 3154 53676 3164 53732
rect 3220 53676 3836 53732
rect 3892 53676 4172 53732
rect 4228 53676 4238 53732
rect 4918 53676 4956 53732
rect 5012 53676 5022 53732
rect 5394 53676 5404 53732
rect 5460 53676 5628 53732
rect 5684 53676 6188 53732
rect 6244 53676 6524 53732
rect 6580 53676 6590 53732
rect 6962 53676 6972 53732
rect 7028 53676 7084 53732
rect 7140 53676 7150 53732
rect 7522 53676 7532 53732
rect 7588 53676 8652 53732
rect 8708 53676 8876 53732
rect 8932 53676 9212 53732
rect 9268 53676 10332 53732
rect 10388 53676 10398 53732
rect 2034 53564 2044 53620
rect 2100 53564 6860 53620
rect 6916 53564 6926 53620
rect 7186 53564 7196 53620
rect 7252 53564 8988 53620
rect 9044 53564 9054 53620
rect 12348 53508 12404 53900
rect 17378 53788 17388 53844
rect 17444 53788 17724 53844
rect 17780 53788 18508 53844
rect 18564 53788 18574 53844
rect 19618 53788 19628 53844
rect 19684 53788 20412 53844
rect 20468 53788 20478 53844
rect 22278 53788 22316 53844
rect 22372 53788 22382 53844
rect 26002 53788 26012 53844
rect 26068 53788 29708 53844
rect 29764 53788 29774 53844
rect 40562 53788 40572 53844
rect 40628 53788 41692 53844
rect 41748 53788 41758 53844
rect 44706 53788 44716 53844
rect 44772 53788 45948 53844
rect 46004 53788 46014 53844
rect 12562 53676 12572 53732
rect 12628 53676 13692 53732
rect 13748 53676 14700 53732
rect 14756 53676 14766 53732
rect 17266 53676 17276 53732
rect 17332 53676 18732 53732
rect 18788 53676 18798 53732
rect 22390 53676 22428 53732
rect 22484 53676 23212 53732
rect 23268 53676 23278 53732
rect 24182 53676 24220 53732
rect 24276 53676 24286 53732
rect 27458 53676 27468 53732
rect 27524 53676 28700 53732
rect 28756 53676 28766 53732
rect 29586 53676 29596 53732
rect 29652 53676 29932 53732
rect 29988 53676 30604 53732
rect 30660 53676 30670 53732
rect 38322 53676 38332 53732
rect 38388 53676 39564 53732
rect 39620 53676 39630 53732
rect 46834 53676 46844 53732
rect 46900 53676 48524 53732
rect 48580 53676 50092 53732
rect 50148 53676 50158 53732
rect 52210 53676 52220 53732
rect 52276 53676 52556 53732
rect 52612 53676 53900 53732
rect 53956 53676 53966 53732
rect 19058 53564 19068 53620
rect 19124 53564 22988 53620
rect 23044 53564 23436 53620
rect 23492 53564 23502 53620
rect 25900 53564 28252 53620
rect 28308 53564 28318 53620
rect 32722 53564 32732 53620
rect 32788 53564 33404 53620
rect 33460 53564 33470 53620
rect 35074 53564 35084 53620
rect 35140 53564 36092 53620
rect 36148 53564 37548 53620
rect 37604 53564 37614 53620
rect 48178 53564 48188 53620
rect 48244 53564 49084 53620
rect 49140 53564 49150 53620
rect 3042 53452 3052 53508
rect 3108 53452 5404 53508
rect 5460 53452 5470 53508
rect 6066 53452 6076 53508
rect 6132 53452 6636 53508
rect 6692 53452 6702 53508
rect 7970 53452 7980 53508
rect 8036 53452 11676 53508
rect 11732 53452 11742 53508
rect 12348 53452 14924 53508
rect 14980 53452 14990 53508
rect 15334 53452 15372 53508
rect 15428 53452 15438 53508
rect 19516 53452 22652 53508
rect 22708 53452 22718 53508
rect 22866 53452 22876 53508
rect 22932 53452 23772 53508
rect 23828 53452 24668 53508
rect 24724 53452 24734 53508
rect 7980 53396 8036 53452
rect 19516 53396 19572 53452
rect 25900 53396 25956 53564
rect 35186 53452 35196 53508
rect 35252 53452 36652 53508
rect 36708 53452 36718 53508
rect 47954 53452 47964 53508
rect 48020 53452 49196 53508
rect 49252 53452 49868 53508
rect 49924 53452 49934 53508
rect 2930 53340 2940 53396
rect 2996 53340 3164 53396
rect 3220 53340 3230 53396
rect 5058 53340 5068 53396
rect 5124 53340 8036 53396
rect 12898 53340 12908 53396
rect 12964 53340 19516 53396
rect 19572 53340 19582 53396
rect 22306 53340 22316 53396
rect 22372 53340 25676 53396
rect 25732 53340 25900 53396
rect 25956 53340 25966 53396
rect 28018 53340 28028 53396
rect 28084 53340 45276 53396
rect 45332 53340 45342 53396
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 2940 53228 3724 53284
rect 3780 53228 6748 53284
rect 6804 53228 6814 53284
rect 6962 53228 6972 53284
rect 7028 53228 13804 53284
rect 13860 53228 13870 53284
rect 16118 53228 16156 53284
rect 16212 53228 16222 53284
rect 17154 53228 17164 53284
rect 17220 53228 19068 53284
rect 19124 53228 19134 53284
rect 22754 53228 22764 53284
rect 22820 53228 24220 53284
rect 24276 53228 24286 53284
rect 42130 53228 42140 53284
rect 42196 53228 42700 53284
rect 42756 53228 42924 53284
rect 42980 53228 42990 53284
rect 2940 53172 2996 53228
rect 2156 53116 2716 53172
rect 2772 53116 2782 53172
rect 2930 53116 2940 53172
rect 2996 53116 3006 53172
rect 4946 53116 4956 53172
rect 5012 53116 6300 53172
rect 6356 53116 6366 53172
rect 9090 53116 9100 53172
rect 9156 53116 9884 53172
rect 9940 53116 9950 53172
rect 10098 53116 10108 53172
rect 10164 53116 11900 53172
rect 11956 53116 12684 53172
rect 12740 53116 12750 53172
rect 14578 53116 14588 53172
rect 14644 53116 21420 53172
rect 21476 53116 21486 53172
rect 22530 53116 22540 53172
rect 22596 53116 22876 53172
rect 22932 53116 24892 53172
rect 24948 53116 24958 53172
rect 26002 53116 26012 53172
rect 26068 53116 31948 53172
rect 2156 52724 2212 53116
rect 31892 53060 31948 53116
rect 2370 53004 2380 53060
rect 2436 53004 2446 53060
rect 5394 53004 5404 53060
rect 5460 53004 11116 53060
rect 11172 53004 13580 53060
rect 13636 53004 13646 53060
rect 17042 53004 17052 53060
rect 17108 53004 19852 53060
rect 19908 53004 19918 53060
rect 21186 53004 21196 53060
rect 21252 53004 21644 53060
rect 21700 53004 21980 53060
rect 22036 53004 22988 53060
rect 23044 53004 24668 53060
rect 24724 53004 24734 53060
rect 25666 53004 25676 53060
rect 25732 53004 29036 53060
rect 29092 53004 29102 53060
rect 31892 53004 47292 53060
rect 47348 53004 47358 53060
rect 2380 52836 2436 53004
rect 2818 52892 2828 52948
rect 2884 52892 3276 52948
rect 3332 52892 5516 52948
rect 5572 52892 5582 52948
rect 7158 52892 7196 52948
rect 7252 52892 7262 52948
rect 12338 52892 12348 52948
rect 12404 52892 13524 52948
rect 14802 52892 14812 52948
rect 14868 52892 17276 52948
rect 17332 52892 17342 52948
rect 18050 52892 18060 52948
rect 18116 52892 18126 52948
rect 20626 52892 20636 52948
rect 20692 52892 20860 52948
rect 20916 52892 22316 52948
rect 22372 52892 22540 52948
rect 22596 52892 22606 52948
rect 23622 52892 23660 52948
rect 23716 52892 23726 52948
rect 24182 52892 24220 52948
rect 24276 52892 24286 52948
rect 26338 52892 26348 52948
rect 26404 52892 27020 52948
rect 27076 52892 28588 52948
rect 28644 52892 28654 52948
rect 33058 52892 33068 52948
rect 33124 52892 33628 52948
rect 33684 52892 33694 52948
rect 13468 52836 13524 52892
rect 18060 52836 18116 52892
rect 2380 52780 3052 52836
rect 3108 52780 3118 52836
rect 3378 52780 3388 52836
rect 3444 52780 3500 52836
rect 3556 52780 3566 52836
rect 7298 52780 7308 52836
rect 7364 52780 7756 52836
rect 7812 52780 7822 52836
rect 8082 52780 8092 52836
rect 8148 52780 8316 52836
rect 8372 52780 13132 52836
rect 13188 52780 13198 52836
rect 13458 52780 13468 52836
rect 13524 52780 14364 52836
rect 14420 52780 14430 52836
rect 15250 52780 15260 52836
rect 15316 52780 16044 52836
rect 16100 52780 18116 52836
rect 18274 52780 18284 52836
rect 18340 52780 18396 52836
rect 18452 52780 18462 52836
rect 18918 52780 18956 52836
rect 19012 52780 19022 52836
rect 22418 52780 22428 52836
rect 22484 52780 23324 52836
rect 23380 52780 23390 52836
rect 23874 52780 23884 52836
rect 23940 52780 25004 52836
rect 25060 52780 25070 52836
rect 26852 52780 27244 52836
rect 27300 52780 27310 52836
rect 39554 52780 39564 52836
rect 39620 52780 40348 52836
rect 40404 52780 40414 52836
rect 47730 52780 47740 52836
rect 47796 52780 48636 52836
rect 48692 52780 48702 52836
rect 49074 52780 49084 52836
rect 49140 52780 50092 52836
rect 50148 52780 50158 52836
rect 26852 52724 26908 52780
rect 2146 52668 2156 52724
rect 2212 52668 2222 52724
rect 2818 52668 2828 52724
rect 2884 52668 4956 52724
rect 5012 52668 5022 52724
rect 6850 52668 6860 52724
rect 6916 52668 7644 52724
rect 7700 52668 9436 52724
rect 9492 52668 9502 52724
rect 14914 52668 14924 52724
rect 14980 52668 16268 52724
rect 16324 52668 16492 52724
rect 16548 52668 16558 52724
rect 23426 52668 23436 52724
rect 23492 52668 23996 52724
rect 24052 52668 26908 52724
rect 10322 52556 10332 52612
rect 10388 52556 10892 52612
rect 10948 52556 11228 52612
rect 11284 52556 12236 52612
rect 12292 52556 12302 52612
rect 13794 52556 13804 52612
rect 13860 52556 19292 52612
rect 19348 52556 21756 52612
rect 21812 52556 22204 52612
rect 22260 52556 23100 52612
rect 23156 52556 26124 52612
rect 26180 52556 26796 52612
rect 26852 52556 26862 52612
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 13122 52444 13132 52500
rect 13188 52444 15372 52500
rect 15428 52444 15438 52500
rect 15922 52444 15932 52500
rect 15988 52444 19404 52500
rect 19460 52444 20636 52500
rect 20692 52444 20702 52500
rect 26852 52444 28364 52500
rect 28420 52444 28430 52500
rect 26852 52388 26908 52444
rect 1026 52332 1036 52388
rect 1092 52332 4284 52388
rect 4340 52332 4350 52388
rect 4508 52332 6972 52388
rect 7028 52332 7038 52388
rect 11666 52332 11676 52388
rect 11732 52332 14252 52388
rect 14308 52332 15148 52388
rect 16034 52332 16044 52388
rect 16100 52332 18284 52388
rect 18340 52332 18350 52388
rect 20514 52332 20524 52388
rect 20580 52332 25340 52388
rect 25396 52332 26348 52388
rect 26404 52332 26908 52388
rect 4508 52276 4564 52332
rect 15092 52276 15148 52332
rect 1250 52220 1260 52276
rect 1316 52220 1596 52276
rect 1652 52220 1820 52276
rect 1876 52220 1886 52276
rect 3154 52220 3164 52276
rect 3220 52220 4396 52276
rect 4452 52220 4564 52276
rect 5282 52220 5292 52276
rect 5348 52220 6076 52276
rect 6132 52220 6142 52276
rect 8502 52220 8540 52276
rect 8596 52220 8606 52276
rect 9986 52220 9996 52276
rect 10052 52220 11340 52276
rect 11396 52220 13804 52276
rect 13860 52220 13870 52276
rect 15092 52220 16940 52276
rect 16996 52220 17006 52276
rect 22306 52220 22316 52276
rect 22372 52220 22932 52276
rect 39330 52220 39340 52276
rect 39396 52220 39900 52276
rect 39956 52220 39966 52276
rect 52658 52220 52668 52276
rect 52724 52220 53900 52276
rect 53956 52220 53966 52276
rect 3014 52108 3052 52164
rect 3108 52108 3118 52164
rect 4834 52108 4844 52164
rect 4900 52108 4956 52164
rect 5012 52108 5022 52164
rect 8418 52108 8428 52164
rect 8484 52108 9100 52164
rect 9156 52108 9166 52164
rect 12422 52108 12460 52164
rect 12516 52108 12526 52164
rect 12982 52108 13020 52164
rect 13076 52108 13086 52164
rect 15138 52108 15148 52164
rect 15204 52108 15932 52164
rect 15988 52108 15998 52164
rect 17266 52108 17276 52164
rect 17332 52108 17836 52164
rect 17892 52108 20636 52164
rect 20692 52108 20702 52164
rect 20850 52108 20860 52164
rect 20916 52108 21868 52164
rect 21924 52108 21934 52164
rect 22418 52108 22428 52164
rect 22484 52108 22540 52164
rect 22596 52108 22606 52164
rect 10406 51996 10444 52052
rect 10500 51996 10510 52052
rect 14018 51996 14028 52052
rect 14084 51996 14812 52052
rect 14868 51996 14878 52052
rect 15092 51996 15372 52052
rect 15428 51996 15438 52052
rect 17154 51996 17164 52052
rect 17220 51996 18172 52052
rect 18228 51996 21084 52052
rect 21140 51996 21756 52052
rect 21812 51996 21822 52052
rect 15092 51940 15148 51996
rect 22540 51940 22596 52108
rect 1922 51884 1932 51940
rect 1988 51884 2268 51940
rect 2324 51884 2604 51940
rect 2660 51884 3164 51940
rect 3220 51884 3230 51940
rect 6290 51884 6300 51940
rect 6356 51884 11116 51940
rect 11172 51884 12460 51940
rect 12516 51884 12526 51940
rect 14466 51884 14476 51940
rect 14532 51884 15148 51940
rect 18274 51884 18284 51940
rect 18340 51884 20300 51940
rect 20356 51884 20366 51940
rect 21634 51884 21644 51940
rect 21700 51884 22596 51940
rect 22876 51828 22932 52220
rect 23314 52108 23324 52164
rect 23380 52108 23772 52164
rect 23828 52108 23838 52164
rect 24332 52108 25676 52164
rect 25732 52108 25742 52164
rect 27906 52108 27916 52164
rect 27972 52108 28084 52164
rect 28242 52108 28252 52164
rect 28308 52108 29708 52164
rect 29764 52108 29774 52164
rect 39218 52108 39228 52164
rect 39284 52108 39564 52164
rect 39620 52108 39788 52164
rect 39844 52108 41132 52164
rect 41188 52108 41198 52164
rect 45714 52108 45724 52164
rect 45780 52108 46172 52164
rect 46228 52108 46238 52164
rect 52434 52108 52444 52164
rect 52500 52108 53564 52164
rect 53620 52108 53630 52164
rect 24332 52052 24388 52108
rect 28028 52052 28084 52108
rect 24322 51996 24332 52052
rect 24388 51996 24398 52052
rect 27122 51996 27132 52052
rect 27188 51996 27804 52052
rect 27860 51996 27870 52052
rect 28028 51996 28700 52052
rect 28756 51996 28766 52052
rect 33282 51996 33292 52052
rect 33348 51996 33740 52052
rect 33796 51996 33806 52052
rect 23090 51884 23100 51940
rect 23156 51884 24444 51940
rect 24500 51884 25228 51940
rect 25284 51884 25294 51940
rect 6626 51772 6636 51828
rect 6692 51772 7644 51828
rect 7700 51772 7710 51828
rect 8194 51772 8204 51828
rect 8260 51772 11564 51828
rect 11620 51772 12348 51828
rect 12404 51772 12414 51828
rect 18834 51772 18844 51828
rect 18900 51772 19404 51828
rect 19460 51772 19470 51828
rect 22876 51772 23212 51828
rect 23268 51772 23278 51828
rect 24098 51772 24108 51828
rect 24164 51772 24780 51828
rect 24836 51772 24846 51828
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 9986 51660 9996 51716
rect 10052 51660 11452 51716
rect 11508 51660 11518 51716
rect 21522 51660 21532 51716
rect 21588 51660 21598 51716
rect 30034 51660 30044 51716
rect 30100 51660 30716 51716
rect 30772 51660 31388 51716
rect 31444 51660 31454 51716
rect 21532 51604 21588 51660
rect 4162 51548 4172 51604
rect 4228 51548 4844 51604
rect 4900 51548 4910 51604
rect 5394 51548 5404 51604
rect 5460 51548 5740 51604
rect 5796 51548 6860 51604
rect 6916 51548 6926 51604
rect 15810 51548 15820 51604
rect 15876 51548 17164 51604
rect 17220 51548 17230 51604
rect 21532 51548 25004 51604
rect 25060 51548 25070 51604
rect 30146 51548 30156 51604
rect 30212 51548 31276 51604
rect 31332 51548 31342 51604
rect 36530 51548 36540 51604
rect 36596 51548 37548 51604
rect 37604 51548 37614 51604
rect 6738 51436 6748 51492
rect 6804 51436 7084 51492
rect 7140 51436 7150 51492
rect 8082 51436 8092 51492
rect 8148 51436 13692 51492
rect 13748 51436 14140 51492
rect 14196 51436 14206 51492
rect 17714 51436 17724 51492
rect 17780 51436 21532 51492
rect 21588 51436 21598 51492
rect 24556 51380 24612 51548
rect 45266 51436 45276 51492
rect 45332 51436 47404 51492
rect 47460 51436 47470 51492
rect 3490 51324 3500 51380
rect 3556 51324 3612 51380
rect 3668 51324 3678 51380
rect 6850 51324 6860 51380
rect 6916 51324 8204 51380
rect 8260 51324 8270 51380
rect 8642 51324 8652 51380
rect 8708 51324 11116 51380
rect 11172 51324 11182 51380
rect 14242 51324 14252 51380
rect 14308 51324 16044 51380
rect 16100 51324 16110 51380
rect 24546 51324 24556 51380
rect 24612 51324 24622 51380
rect 26114 51324 26124 51380
rect 26180 51324 28028 51380
rect 28084 51324 28094 51380
rect 31892 51324 32620 51380
rect 32676 51324 33964 51380
rect 34020 51324 34030 51380
rect 36306 51324 36316 51380
rect 36372 51324 37324 51380
rect 37380 51324 37390 51380
rect 42914 51324 42924 51380
rect 42980 51324 43148 51380
rect 43204 51324 43214 51380
rect 44034 51324 44044 51380
rect 44100 51324 44940 51380
rect 44996 51324 47180 51380
rect 47236 51324 47246 51380
rect 31892 51268 31948 51324
rect 1922 51212 1932 51268
rect 1988 51212 2156 51268
rect 2212 51212 2222 51268
rect 3154 51212 3164 51268
rect 3220 51212 5404 51268
rect 5460 51212 5470 51268
rect 7746 51212 7756 51268
rect 7812 51212 8876 51268
rect 8932 51212 9324 51268
rect 9380 51212 10444 51268
rect 10500 51212 17612 51268
rect 17668 51212 17678 51268
rect 18946 51212 18956 51268
rect 19012 51212 19740 51268
rect 19796 51212 19806 51268
rect 31042 51212 31052 51268
rect 31108 51212 31948 51268
rect 32722 51212 32732 51268
rect 32788 51212 34636 51268
rect 34692 51212 34702 51268
rect 3798 51100 3836 51156
rect 3892 51100 3902 51156
rect 4050 51100 4060 51156
rect 4116 51100 4396 51156
rect 4452 51100 4462 51156
rect 6178 51100 6188 51156
rect 6244 51100 9772 51156
rect 9828 51100 9838 51156
rect 11554 51100 11564 51156
rect 11620 51100 18116 51156
rect 4060 50820 4116 51100
rect 18060 51044 18116 51100
rect 31892 51100 44156 51156
rect 44212 51100 44222 51156
rect 45042 51100 45052 51156
rect 45108 51100 46284 51156
rect 46340 51100 47068 51156
rect 47124 51100 47134 51156
rect 12562 50988 12572 51044
rect 12628 50988 16492 51044
rect 16548 50988 16558 51044
rect 18060 50988 20972 51044
rect 21028 50988 21038 51044
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 31892 50932 31948 51100
rect 32050 50988 32060 51044
rect 32116 50988 32396 51044
rect 32452 50988 33740 51044
rect 33796 50988 33806 51044
rect 36418 50988 36428 51044
rect 36484 50988 37660 51044
rect 37716 50988 39788 51044
rect 39844 50988 39854 51044
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 6962 50876 6972 50932
rect 7028 50876 7644 50932
rect 7700 50876 7710 50932
rect 7858 50876 7868 50932
rect 7924 50876 15932 50932
rect 15988 50876 15998 50932
rect 20066 50876 20076 50932
rect 20132 50876 23212 50932
rect 23268 50876 23278 50932
rect 26450 50876 26460 50932
rect 26516 50876 31948 50932
rect 33180 50876 35028 50932
rect 33180 50820 33236 50876
rect 34972 50820 35028 50876
rect 3836 50764 4116 50820
rect 5842 50764 5852 50820
rect 5908 50764 12460 50820
rect 12516 50764 13244 50820
rect 13300 50764 13310 50820
rect 14130 50764 14140 50820
rect 14196 50764 15820 50820
rect 15876 50764 15886 50820
rect 16678 50764 16716 50820
rect 16772 50764 16782 50820
rect 17602 50764 17612 50820
rect 17668 50764 18172 50820
rect 18228 50764 18238 50820
rect 27234 50764 27244 50820
rect 27300 50764 28028 50820
rect 28084 50764 33236 50820
rect 33394 50764 33404 50820
rect 33460 50764 34412 50820
rect 34468 50764 34478 50820
rect 34972 50764 39900 50820
rect 39956 50764 40348 50820
rect 40404 50764 40414 50820
rect 41906 50764 41916 50820
rect 41972 50764 42588 50820
rect 42644 50764 43260 50820
rect 43316 50764 43326 50820
rect 3836 50708 3892 50764
rect 2566 50652 2604 50708
rect 2660 50652 3164 50708
rect 3220 50652 3230 50708
rect 3826 50652 3836 50708
rect 3892 50652 3902 50708
rect 4498 50652 4508 50708
rect 4564 50652 5068 50708
rect 5124 50652 5134 50708
rect 5292 50652 5740 50708
rect 5796 50652 6188 50708
rect 6244 50652 6254 50708
rect 6850 50652 6860 50708
rect 6916 50652 7980 50708
rect 8036 50652 8046 50708
rect 8978 50652 8988 50708
rect 9044 50652 10220 50708
rect 10276 50652 10286 50708
rect 11666 50652 11676 50708
rect 11732 50652 12236 50708
rect 12292 50652 14700 50708
rect 14756 50652 14766 50708
rect 22306 50652 22316 50708
rect 22372 50652 22876 50708
rect 22932 50652 22942 50708
rect 34066 50652 34076 50708
rect 34132 50652 35868 50708
rect 35924 50652 35934 50708
rect 36866 50652 36876 50708
rect 36932 50652 37660 50708
rect 37716 50652 37726 50708
rect 38546 50652 38556 50708
rect 38612 50652 39340 50708
rect 39396 50652 39406 50708
rect 5292 50596 5348 50652
rect 2146 50540 2156 50596
rect 2212 50540 2940 50596
rect 2996 50540 3388 50596
rect 3444 50540 3454 50596
rect 3714 50540 3724 50596
rect 3780 50540 3836 50596
rect 3892 50540 3902 50596
rect 4050 50540 4060 50596
rect 4116 50540 4844 50596
rect 4900 50540 5348 50596
rect 6066 50540 6076 50596
rect 6132 50540 7868 50596
rect 7924 50540 8652 50596
rect 8708 50540 8718 50596
rect 9062 50540 9100 50596
rect 9156 50540 9166 50596
rect 10882 50540 10892 50596
rect 10948 50540 11228 50596
rect 11284 50540 11294 50596
rect 12674 50540 12684 50596
rect 12740 50540 14028 50596
rect 14084 50540 14094 50596
rect 17042 50540 17052 50596
rect 17108 50540 18396 50596
rect 18452 50540 18462 50596
rect 19964 50540 23772 50596
rect 23828 50540 23838 50596
rect 26898 50540 26908 50596
rect 26964 50540 27244 50596
rect 27300 50540 27916 50596
rect 27972 50540 27982 50596
rect 36754 50540 36764 50596
rect 36820 50540 37884 50596
rect 37940 50540 37950 50596
rect 41570 50540 41580 50596
rect 41636 50540 42924 50596
rect 42980 50540 42990 50596
rect 47394 50540 47404 50596
rect 47460 50540 53788 50596
rect 53844 50540 54236 50596
rect 54292 50540 54302 50596
rect 56242 50540 56252 50596
rect 56308 50540 56812 50596
rect 56868 50540 56878 50596
rect 19964 50484 20020 50540
rect 1810 50428 1820 50484
rect 1876 50428 3948 50484
rect 4004 50428 4014 50484
rect 5842 50428 5852 50484
rect 5908 50428 7644 50484
rect 7700 50428 7710 50484
rect 9762 50428 9772 50484
rect 9828 50428 9838 50484
rect 11442 50428 11452 50484
rect 11508 50428 13804 50484
rect 13860 50428 13870 50484
rect 15138 50428 15148 50484
rect 15204 50428 15596 50484
rect 15652 50428 15662 50484
rect 15922 50428 15932 50484
rect 15988 50428 20020 50484
rect 20178 50428 20188 50484
rect 20244 50428 22876 50484
rect 22932 50428 22942 50484
rect 25106 50428 25116 50484
rect 25172 50428 26236 50484
rect 26292 50428 26302 50484
rect 28242 50428 28252 50484
rect 28308 50428 28700 50484
rect 28756 50428 29708 50484
rect 29764 50428 29774 50484
rect 30594 50428 30604 50484
rect 30660 50428 31276 50484
rect 31332 50428 31342 50484
rect 33058 50428 33068 50484
rect 33124 50428 34188 50484
rect 34244 50428 34254 50484
rect 38546 50428 38556 50484
rect 38612 50428 39116 50484
rect 39172 50428 39182 50484
rect 40338 50428 40348 50484
rect 40404 50428 40964 50484
rect 48402 50428 48412 50484
rect 48468 50428 53900 50484
rect 53956 50428 54124 50484
rect 54180 50428 54190 50484
rect 9772 50372 9828 50428
rect 40898 50372 40908 50428
rect 40964 50372 40974 50428
rect 3042 50316 3052 50372
rect 3108 50316 3500 50372
rect 3556 50316 3566 50372
rect 4050 50316 4060 50372
rect 4116 50316 5740 50372
rect 5796 50316 5806 50372
rect 6738 50316 6748 50372
rect 6804 50316 7980 50372
rect 8036 50316 8046 50372
rect 8418 50316 8428 50372
rect 8484 50316 8988 50372
rect 9044 50316 9054 50372
rect 9772 50316 10556 50372
rect 10612 50316 18732 50372
rect 18788 50316 20972 50372
rect 21028 50316 21038 50372
rect 23314 50316 23324 50372
rect 23380 50316 24108 50372
rect 24164 50316 24174 50372
rect 26002 50316 26012 50372
rect 26068 50316 28924 50372
rect 28980 50316 30492 50372
rect 30548 50316 32172 50372
rect 32228 50316 32620 50372
rect 32676 50316 32686 50372
rect 44594 50316 44604 50372
rect 44660 50316 45836 50372
rect 45892 50316 46060 50372
rect 46116 50316 46956 50372
rect 47012 50316 47022 50372
rect 51762 50316 51772 50372
rect 51828 50316 53452 50372
rect 53508 50316 53518 50372
rect 8988 50260 9044 50316
rect 3378 50204 3388 50260
rect 3444 50204 4956 50260
rect 5012 50204 6524 50260
rect 6580 50204 7084 50260
rect 7140 50204 7150 50260
rect 8988 50204 11900 50260
rect 11956 50204 14700 50260
rect 14756 50204 14766 50260
rect 15586 50204 15596 50260
rect 15652 50204 16156 50260
rect 16212 50204 17836 50260
rect 17892 50204 18004 50260
rect 18162 50204 18172 50260
rect 18228 50204 18620 50260
rect 18676 50204 18686 50260
rect 22194 50204 22204 50260
rect 22260 50204 23100 50260
rect 23156 50204 23166 50260
rect 26852 50204 35980 50260
rect 36036 50204 36046 50260
rect 52546 50204 52556 50260
rect 52612 50204 53116 50260
rect 53172 50204 53676 50260
rect 53732 50204 53742 50260
rect 17948 50148 18004 50204
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 26852 50148 26908 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 2930 50092 2940 50148
rect 2996 50092 3612 50148
rect 3668 50092 3678 50148
rect 6962 50092 6972 50148
rect 7028 50092 14084 50148
rect 14802 50092 14812 50148
rect 14868 50092 17724 50148
rect 17780 50092 17790 50148
rect 17948 50092 19068 50148
rect 19124 50092 19134 50148
rect 19282 50092 19292 50148
rect 19348 50092 19404 50148
rect 19460 50092 19470 50148
rect 20850 50092 20860 50148
rect 20916 50092 26908 50148
rect 28018 50092 28028 50148
rect 28084 50092 34076 50148
rect 34132 50092 34142 50148
rect 3490 49980 3500 50036
rect 3556 49980 5628 50036
rect 5684 49980 5694 50036
rect 8306 49980 8316 50036
rect 8372 49980 10668 50036
rect 10724 49980 10734 50036
rect 10882 49980 10892 50036
rect 10948 49980 11452 50036
rect 11508 49980 11518 50036
rect 11666 49980 11676 50036
rect 11732 49980 11742 50036
rect 11676 49924 11732 49980
rect 914 49868 924 49924
rect 980 49868 4732 49924
rect 4788 49868 9996 49924
rect 10052 49868 10062 49924
rect 11452 49868 12460 49924
rect 12516 49868 12526 49924
rect 11452 49812 11508 49868
rect 14028 49812 14084 50092
rect 15698 49980 15708 50036
rect 15764 49980 16380 50036
rect 16436 49980 16446 50036
rect 19394 49980 19404 50036
rect 19460 49980 21308 50036
rect 21364 49980 22540 50036
rect 22596 49980 22764 50036
rect 22820 49980 22830 50036
rect 25666 49980 25676 50036
rect 25732 49980 26908 50036
rect 30594 49980 30604 50036
rect 30660 49980 33852 50036
rect 33908 49980 33918 50036
rect 52098 49980 52108 50036
rect 52164 49980 53116 50036
rect 53172 49980 53182 50036
rect 14466 49868 14476 49924
rect 14532 49868 16940 49924
rect 16996 49868 17276 49924
rect 17332 49868 17342 49924
rect 19842 49868 19852 49924
rect 19908 49868 21644 49924
rect 21700 49868 22092 49924
rect 22148 49868 22158 49924
rect 26852 49812 26908 49980
rect 31714 49868 31724 49924
rect 31780 49868 33964 49924
rect 34020 49868 34030 49924
rect 39666 49868 39676 49924
rect 39732 49868 40348 49924
rect 40404 49868 48412 49924
rect 48468 49868 48478 49924
rect 57586 49868 57596 49924
rect 57652 49868 58492 49924
rect 58548 49868 58558 49924
rect 2370 49756 2380 49812
rect 2436 49756 3276 49812
rect 3332 49756 3948 49812
rect 4004 49756 8372 49812
rect 8530 49756 8540 49812
rect 8596 49756 9548 49812
rect 9604 49756 9614 49812
rect 11442 49756 11452 49812
rect 11508 49756 11518 49812
rect 12338 49756 12348 49812
rect 12404 49756 12414 49812
rect 13766 49756 13804 49812
rect 13860 49756 13870 49812
rect 14028 49756 15148 49812
rect 17602 49756 17612 49812
rect 17668 49756 18508 49812
rect 18564 49756 18574 49812
rect 20738 49756 20748 49812
rect 20804 49756 22204 49812
rect 22260 49756 22270 49812
rect 26852 49756 27356 49812
rect 27412 49756 27916 49812
rect 27972 49756 29540 49812
rect 29698 49756 29708 49812
rect 29764 49756 32396 49812
rect 32452 49756 35308 49812
rect 35364 49756 36596 49812
rect 43586 49756 43596 49812
rect 8316 49700 8372 49756
rect 2902 49644 2940 49700
rect 2996 49644 3006 49700
rect 5170 49644 5180 49700
rect 5236 49644 6300 49700
rect 6356 49644 7308 49700
rect 7364 49644 8092 49700
rect 8148 49644 8158 49700
rect 8306 49644 8316 49700
rect 8372 49644 11228 49700
rect 11284 49644 11294 49700
rect 12348 49588 12404 49756
rect 15092 49700 15148 49756
rect 29484 49700 29540 49756
rect 36540 49700 36596 49756
rect 43652 49700 43708 49812
rect 48178 49756 48188 49812
rect 48244 49756 49084 49812
rect 49140 49756 49532 49812
rect 49588 49756 50204 49812
rect 50260 49756 50270 49812
rect 56354 49756 56364 49812
rect 56420 49756 56430 49812
rect 56364 49700 56420 49756
rect 13234 49644 13244 49700
rect 13300 49644 14812 49700
rect 14868 49644 14878 49700
rect 15092 49644 15260 49700
rect 15316 49644 16044 49700
rect 16100 49644 16110 49700
rect 16930 49644 16940 49700
rect 16996 49644 17388 49700
rect 17444 49644 18956 49700
rect 19012 49644 19022 49700
rect 24770 49644 24780 49700
rect 24836 49644 29148 49700
rect 29204 49644 29214 49700
rect 29484 49644 30268 49700
rect 30324 49644 32508 49700
rect 32564 49644 32574 49700
rect 34626 49644 34636 49700
rect 34692 49644 35756 49700
rect 35812 49644 35822 49700
rect 36530 49644 36540 49700
rect 36596 49644 36764 49700
rect 36820 49644 36830 49700
rect 43652 49644 43820 49700
rect 43876 49644 45164 49700
rect 45220 49644 45230 49700
rect 48514 49644 48524 49700
rect 48580 49644 49756 49700
rect 49812 49644 49822 49700
rect 53778 49644 53788 49700
rect 53844 49644 54460 49700
rect 54516 49644 54526 49700
rect 55906 49644 55916 49700
rect 55972 49644 56700 49700
rect 56756 49644 56766 49700
rect 14812 49588 14868 49644
rect 5058 49532 5068 49588
rect 5124 49532 5852 49588
rect 5908 49532 5918 49588
rect 6710 49532 6748 49588
rect 6804 49532 6814 49588
rect 10770 49532 10780 49588
rect 10836 49532 10892 49588
rect 10948 49532 11004 49588
rect 11060 49532 12796 49588
rect 12852 49532 13132 49588
rect 13188 49532 13198 49588
rect 14812 49532 18228 49588
rect 51426 49532 51436 49588
rect 51492 49532 51884 49588
rect 51940 49532 51950 49588
rect 18172 49476 18228 49532
rect 6850 49420 6860 49476
rect 6916 49420 9212 49476
rect 9268 49420 9278 49476
rect 11712 49420 11788 49476
rect 11844 49420 17836 49476
rect 17892 49420 17902 49476
rect 18162 49420 18172 49476
rect 18228 49420 18396 49476
rect 18452 49420 18462 49476
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 5618 49308 5628 49364
rect 5684 49308 10108 49364
rect 10164 49308 11452 49364
rect 11508 49308 11518 49364
rect 15250 49308 15260 49364
rect 15316 49308 15484 49364
rect 15540 49308 18060 49364
rect 18116 49308 18126 49364
rect 26450 49308 26460 49364
rect 26516 49308 28868 49364
rect 1586 49196 1596 49252
rect 1652 49196 8876 49252
rect 8932 49196 8942 49252
rect 9762 49196 9772 49252
rect 9828 49196 11676 49252
rect 11732 49196 11742 49252
rect 12114 49196 12124 49252
rect 12180 49196 14924 49252
rect 14980 49196 14990 49252
rect 16416 49196 16492 49252
rect 16548 49196 17500 49252
rect 17556 49196 17566 49252
rect 24658 49196 24668 49252
rect 24724 49196 25004 49252
rect 25060 49196 27020 49252
rect 27076 49196 28364 49252
rect 28420 49196 28430 49252
rect 28812 49140 28868 49308
rect 43652 49308 50876 49364
rect 50932 49308 52332 49364
rect 52388 49308 53564 49364
rect 53620 49308 54124 49364
rect 54180 49308 54190 49364
rect 55346 49308 55356 49364
rect 43652 49252 43708 49308
rect 55412 49252 55468 49364
rect 29810 49196 29820 49252
rect 29876 49196 43708 49252
rect 47170 49196 47180 49252
rect 47236 49196 48412 49252
rect 48468 49196 48478 49252
rect 55412 49196 55580 49252
rect 55636 49196 55646 49252
rect 3332 49084 3612 49140
rect 3668 49084 3678 49140
rect 5506 49084 5516 49140
rect 5572 49084 6076 49140
rect 6132 49084 6142 49140
rect 6934 49084 6972 49140
rect 7028 49084 7038 49140
rect 7298 49084 7308 49140
rect 7364 49084 8540 49140
rect 8596 49084 8606 49140
rect 11106 49084 11116 49140
rect 11172 49084 12348 49140
rect 12404 49084 12414 49140
rect 14354 49084 14364 49140
rect 14420 49084 16156 49140
rect 16212 49084 16380 49140
rect 16436 49084 16940 49140
rect 16996 49084 17006 49140
rect 18386 49084 18396 49140
rect 18452 49084 20524 49140
rect 20580 49084 20590 49140
rect 20850 49084 20860 49140
rect 20916 49084 23100 49140
rect 23156 49084 23166 49140
rect 26338 49084 26348 49140
rect 26404 49084 27916 49140
rect 27972 49084 27982 49140
rect 28802 49084 28812 49140
rect 28868 49084 30828 49140
rect 30884 49084 30894 49140
rect 32610 49084 32620 49140
rect 32676 49084 37548 49140
rect 37604 49084 38332 49140
rect 38388 49084 38398 49140
rect 3266 48972 3276 49028
rect 3332 48972 3388 49084
rect 6738 48972 6748 49028
rect 6804 48972 10332 49028
rect 10388 48972 10398 49028
rect 10658 48972 10668 49028
rect 10724 48972 11004 49028
rect 11060 48972 11070 49028
rect 12562 48972 12572 49028
rect 12628 48972 13132 49028
rect 13188 48972 13356 49028
rect 13412 48972 13422 49028
rect 14364 48916 14420 49084
rect 14578 48972 14588 49028
rect 14644 48972 15260 49028
rect 15316 48972 15326 49028
rect 15586 48972 15596 49028
rect 15652 48972 17724 49028
rect 17780 48972 17790 49028
rect 20066 48972 20076 49028
rect 20132 48972 21980 49028
rect 22036 48972 22046 49028
rect 25218 48972 25228 49028
rect 25284 48972 26012 49028
rect 26068 48972 26078 49028
rect 35522 48972 35532 49028
rect 35588 48972 36092 49028
rect 36148 48972 36158 49028
rect 44706 48972 44716 49028
rect 44772 48972 45724 49028
rect 45780 48972 45790 49028
rect 56690 48972 56700 49028
rect 56756 48972 58268 49028
rect 58324 48972 58334 49028
rect 2044 48860 3500 48916
rect 3556 48860 4172 48916
rect 4228 48860 4238 48916
rect 8306 48860 8316 48916
rect 8372 48860 14420 48916
rect 14914 48860 14924 48916
rect 14980 48860 16884 48916
rect 18162 48860 18172 48916
rect 18228 48860 21644 48916
rect 21700 48860 21710 48916
rect 22530 48860 22540 48916
rect 22596 48860 24220 48916
rect 24276 48860 24892 48916
rect 24948 48860 24958 48916
rect 25442 48860 25452 48916
rect 25508 48860 26348 48916
rect 26404 48860 26414 48916
rect 26852 48860 30604 48916
rect 30660 48860 30670 48916
rect 40450 48860 40460 48916
rect 40516 48860 41804 48916
rect 41860 48860 41870 48916
rect 43810 48860 43820 48916
rect 43876 48860 46060 48916
rect 46116 48860 46732 48916
rect 46788 48860 46798 48916
rect 51100 48860 51660 48916
rect 51716 48860 51726 48916
rect 52322 48860 52332 48916
rect 52388 48860 53340 48916
rect 53396 48860 53406 48916
rect 2044 48692 2100 48860
rect 3602 48748 3612 48804
rect 3668 48748 4620 48804
rect 4676 48748 4686 48804
rect 6066 48748 6076 48804
rect 6132 48748 7868 48804
rect 7924 48748 7934 48804
rect 8530 48748 8540 48804
rect 8596 48748 8876 48804
rect 8932 48748 8942 48804
rect 9874 48748 9884 48804
rect 9940 48748 10332 48804
rect 10388 48748 11004 48804
rect 11060 48748 11070 48804
rect 12086 48748 12124 48804
rect 12180 48748 12190 48804
rect 12674 48748 12684 48804
rect 12740 48748 14588 48804
rect 14644 48748 15148 48804
rect 15204 48748 15214 48804
rect 16034 48748 16044 48804
rect 16100 48748 16492 48804
rect 16548 48748 16558 48804
rect 16828 48692 16884 48860
rect 23650 48748 23660 48804
rect 23716 48748 24108 48804
rect 24164 48748 26796 48804
rect 26852 48748 26908 48860
rect 51100 48804 51156 48860
rect 27122 48748 27132 48804
rect 27188 48748 27356 48804
rect 27412 48748 27422 48804
rect 33618 48748 33628 48804
rect 33684 48748 33852 48804
rect 33908 48748 33918 48804
rect 40786 48748 40796 48804
rect 40852 48748 42028 48804
rect 42084 48748 42094 48804
rect 43586 48748 43596 48804
rect 43652 48748 44604 48804
rect 44660 48748 44670 48804
rect 48626 48748 48636 48804
rect 48692 48748 51100 48804
rect 51156 48748 51166 48804
rect 51426 48748 51436 48804
rect 51492 48748 51502 48804
rect 55458 48748 55468 48804
rect 55524 48748 57484 48804
rect 57540 48748 57550 48804
rect 2034 48636 2044 48692
rect 2100 48636 2110 48692
rect 4162 48636 4172 48692
rect 4228 48636 5964 48692
rect 6020 48636 6030 48692
rect 7410 48636 7420 48692
rect 7476 48636 7812 48692
rect 7970 48636 7980 48692
rect 8036 48636 8428 48692
rect 8484 48636 8494 48692
rect 10210 48636 10220 48692
rect 10276 48636 12236 48692
rect 12292 48636 12302 48692
rect 14130 48636 14140 48692
rect 14196 48636 14924 48692
rect 14980 48636 15708 48692
rect 15764 48636 15774 48692
rect 16828 48636 19292 48692
rect 19348 48636 19358 48692
rect 23090 48636 23100 48692
rect 23156 48636 23996 48692
rect 24052 48636 25676 48692
rect 25732 48636 25742 48692
rect 31602 48636 31612 48692
rect 31668 48636 34524 48692
rect 34580 48636 34590 48692
rect 35634 48636 35644 48692
rect 35700 48636 37100 48692
rect 37156 48636 37884 48692
rect 37940 48636 37950 48692
rect 7756 48580 7812 48636
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 1250 48524 1260 48580
rect 1316 48524 7532 48580
rect 7588 48524 7598 48580
rect 7756 48524 15596 48580
rect 15652 48524 15662 48580
rect 16146 48524 16156 48580
rect 16212 48524 18396 48580
rect 18452 48524 18462 48580
rect 25778 48524 25788 48580
rect 25844 48524 26684 48580
rect 26740 48524 34804 48580
rect 2258 48412 2268 48468
rect 2324 48412 2492 48468
rect 2548 48412 3052 48468
rect 3108 48412 3118 48468
rect 5954 48412 5964 48468
rect 6020 48412 8988 48468
rect 9044 48412 9054 48468
rect 9986 48412 9996 48468
rect 10052 48412 10220 48468
rect 10276 48412 10286 48468
rect 10406 48412 10444 48468
rect 10500 48412 10510 48468
rect 10994 48412 11004 48468
rect 11060 48412 11676 48468
rect 11732 48412 11788 48468
rect 11844 48412 11854 48468
rect 15092 48412 15484 48468
rect 15540 48412 15550 48468
rect 16930 48412 16940 48468
rect 16996 48412 19180 48468
rect 19236 48412 19246 48468
rect 21046 48412 21084 48468
rect 21140 48412 21150 48468
rect 21410 48412 21420 48468
rect 21476 48412 23436 48468
rect 23492 48412 23502 48468
rect 28354 48412 28364 48468
rect 28420 48412 30044 48468
rect 30100 48412 30492 48468
rect 30548 48412 31052 48468
rect 31108 48412 34300 48468
rect 34356 48412 34366 48468
rect 2370 48300 2380 48356
rect 2436 48300 6748 48356
rect 6804 48300 6814 48356
rect 15092 48244 15148 48412
rect 34748 48356 34804 48524
rect 51436 48468 51492 48748
rect 34962 48412 34972 48468
rect 35028 48412 52668 48468
rect 52724 48412 53116 48468
rect 53172 48412 53182 48468
rect 17910 48300 17948 48356
rect 18004 48300 18014 48356
rect 18274 48300 18284 48356
rect 18340 48300 20860 48356
rect 20916 48300 21308 48356
rect 21364 48300 21374 48356
rect 22642 48300 22652 48356
rect 22708 48300 22988 48356
rect 23044 48300 23324 48356
rect 23380 48300 26572 48356
rect 26628 48300 28252 48356
rect 28308 48300 28318 48356
rect 30818 48300 30828 48356
rect 30884 48300 34412 48356
rect 34468 48300 34478 48356
rect 34748 48300 40684 48356
rect 40740 48300 40750 48356
rect 1474 48188 1484 48244
rect 1540 48188 3052 48244
rect 3108 48188 5572 48244
rect 5842 48188 5852 48244
rect 5908 48188 8428 48244
rect 8484 48188 8494 48244
rect 8642 48188 8652 48244
rect 8708 48188 8746 48244
rect 10210 48188 10220 48244
rect 10276 48188 11340 48244
rect 11396 48188 12572 48244
rect 12628 48188 12638 48244
rect 12898 48188 12908 48244
rect 12964 48188 14140 48244
rect 14196 48188 14206 48244
rect 14354 48188 14364 48244
rect 14420 48188 15148 48244
rect 15922 48188 15932 48244
rect 15988 48188 16492 48244
rect 16548 48188 18508 48244
rect 18564 48188 18574 48244
rect 32722 48188 32732 48244
rect 32788 48188 34076 48244
rect 34132 48188 34142 48244
rect 36418 48188 36428 48244
rect 36484 48188 37884 48244
rect 37940 48188 38444 48244
rect 38500 48188 38510 48244
rect 46162 48188 46172 48244
rect 46228 48188 46844 48244
rect 46900 48188 46910 48244
rect 52434 48188 52444 48244
rect 52500 48188 54796 48244
rect 54852 48188 54862 48244
rect 56802 48188 56812 48244
rect 56868 48188 57932 48244
rect 57988 48188 58380 48244
rect 58436 48188 58446 48244
rect 5516 48132 5572 48188
rect 3490 48076 3500 48132
rect 3556 48076 5292 48132
rect 5348 48076 5358 48132
rect 5516 48076 10892 48132
rect 10948 48076 10958 48132
rect 12002 48076 12012 48132
rect 12068 48076 13356 48132
rect 13412 48076 13422 48132
rect 14914 48076 14924 48132
rect 14980 48076 17612 48132
rect 17668 48076 17836 48132
rect 17892 48076 17902 48132
rect 18946 48076 18956 48132
rect 19012 48076 19628 48132
rect 19684 48076 19694 48132
rect 23548 48076 24444 48132
rect 24500 48076 24780 48132
rect 24836 48076 27356 48132
rect 27412 48076 27422 48132
rect 28802 48076 28812 48132
rect 28868 48076 29932 48132
rect 29988 48076 30156 48132
rect 30212 48076 32956 48132
rect 33012 48076 33022 48132
rect 38770 48076 38780 48132
rect 38836 48076 39676 48132
rect 39732 48076 39742 48132
rect 23548 48020 23604 48076
rect 2818 47964 2828 48020
rect 2884 47964 3724 48020
rect 3780 47964 6188 48020
rect 6244 47964 6254 48020
rect 7858 47964 7868 48020
rect 7924 47964 9772 48020
rect 9828 47964 14924 48020
rect 14980 47964 14990 48020
rect 15474 47964 15484 48020
rect 15540 47964 16716 48020
rect 16772 47964 18172 48020
rect 18228 47964 18238 48020
rect 23538 47964 23548 48020
rect 23604 47964 23614 48020
rect 25666 47964 25676 48020
rect 25732 47964 31164 48020
rect 31220 47964 31230 48020
rect 4022 47852 4060 47908
rect 4116 47852 4126 47908
rect 4834 47852 4844 47908
rect 4900 47852 7980 47908
rect 8036 47852 8046 47908
rect 8754 47852 8764 47908
rect 8820 47852 24668 47908
rect 24724 47852 24734 47908
rect 28466 47852 28476 47908
rect 28532 47852 34972 47908
rect 35028 47852 35038 47908
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 4134 47740 4172 47796
rect 4228 47740 4238 47796
rect 6962 47740 6972 47796
rect 7028 47740 8988 47796
rect 9044 47740 9054 47796
rect 20402 47740 20412 47796
rect 20468 47740 22764 47796
rect 22820 47740 22830 47796
rect 54450 47740 54460 47796
rect 54516 47740 57260 47796
rect 57316 47740 57596 47796
rect 57652 47740 57662 47796
rect 1586 47628 1596 47684
rect 1652 47628 2828 47684
rect 2884 47628 10220 47684
rect 10276 47628 10286 47684
rect 10546 47628 10556 47684
rect 10612 47628 11452 47684
rect 11508 47628 11518 47684
rect 4274 47516 4284 47572
rect 4340 47516 5628 47572
rect 5684 47516 6076 47572
rect 6132 47516 6142 47572
rect 6738 47516 6748 47572
rect 6804 47516 7756 47572
rect 7812 47516 9436 47572
rect 9492 47516 14364 47572
rect 14420 47516 14430 47572
rect 15138 47516 15148 47572
rect 15204 47516 15596 47572
rect 15652 47516 15662 47572
rect 17602 47516 17612 47572
rect 17668 47516 17724 47572
rect 17780 47516 18956 47572
rect 19012 47516 19852 47572
rect 19908 47516 19918 47572
rect 20066 47516 20076 47572
rect 20132 47516 20860 47572
rect 20916 47516 20926 47572
rect 21970 47516 21980 47572
rect 22036 47516 22316 47572
rect 22372 47516 22382 47572
rect 26852 47516 28812 47572
rect 28868 47516 28878 47572
rect 42466 47516 42476 47572
rect 42532 47516 43260 47572
rect 43316 47516 43326 47572
rect 46050 47516 46060 47572
rect 46116 47516 46732 47572
rect 46788 47516 46798 47572
rect 55682 47516 55692 47572
rect 55748 47516 56364 47572
rect 56420 47516 56430 47572
rect 2594 47404 2604 47460
rect 2660 47404 3276 47460
rect 3332 47404 4060 47460
rect 4116 47404 4126 47460
rect 5506 47404 5516 47460
rect 5572 47404 6524 47460
rect 6580 47404 7644 47460
rect 7700 47404 12124 47460
rect 12180 47404 12190 47460
rect 14466 47404 14476 47460
rect 14532 47404 15708 47460
rect 15764 47404 15774 47460
rect 22316 47348 22372 47516
rect 26852 47460 26908 47516
rect 23314 47404 23324 47460
rect 23380 47404 23772 47460
rect 23828 47404 25116 47460
rect 25172 47404 25676 47460
rect 25732 47404 26908 47460
rect 27346 47404 27356 47460
rect 27412 47404 29484 47460
rect 29540 47404 29550 47460
rect 34066 47404 34076 47460
rect 34132 47404 34412 47460
rect 34468 47404 37436 47460
rect 37492 47404 37502 47460
rect 40002 47404 40012 47460
rect 40068 47404 41020 47460
rect 41076 47404 41580 47460
rect 41636 47404 41646 47460
rect 44594 47404 44604 47460
rect 44660 47404 45388 47460
rect 45444 47404 45454 47460
rect 50866 47404 50876 47460
rect 50932 47404 51884 47460
rect 51940 47404 54572 47460
rect 54628 47404 54638 47460
rect 55346 47404 55356 47460
rect 55412 47404 56308 47460
rect 56802 47404 56812 47460
rect 56868 47404 57372 47460
rect 57428 47404 57438 47460
rect 55692 47348 55748 47404
rect 56252 47348 56308 47404
rect 2258 47292 2268 47348
rect 2324 47292 3612 47348
rect 3668 47292 3678 47348
rect 5954 47292 5964 47348
rect 6020 47292 6860 47348
rect 6916 47292 6926 47348
rect 9202 47292 9212 47348
rect 9268 47292 10556 47348
rect 10612 47292 10622 47348
rect 17938 47292 17948 47348
rect 18004 47292 19292 47348
rect 19348 47292 19358 47348
rect 22316 47292 24556 47348
rect 24612 47292 24622 47348
rect 26002 47292 26012 47348
rect 26068 47292 27580 47348
rect 27636 47292 27916 47348
rect 27972 47292 27982 47348
rect 36978 47292 36988 47348
rect 37044 47292 37548 47348
rect 37604 47292 39452 47348
rect 39508 47292 39518 47348
rect 39666 47292 39676 47348
rect 39732 47292 40348 47348
rect 40404 47292 40414 47348
rect 40562 47292 40572 47348
rect 40628 47292 41244 47348
rect 41300 47292 41804 47348
rect 41860 47292 41870 47348
rect 44034 47292 44044 47348
rect 44100 47292 45836 47348
rect 45892 47292 45902 47348
rect 55234 47292 55244 47348
rect 55300 47292 55468 47348
rect 55682 47292 55692 47348
rect 55748 47292 55758 47348
rect 56242 47292 56252 47348
rect 56308 47292 56318 47348
rect 19292 47236 19348 47292
rect 55412 47236 55468 47292
rect 10546 47180 10556 47236
rect 10612 47180 11116 47236
rect 11172 47180 13692 47236
rect 13748 47180 13758 47236
rect 14802 47180 14812 47236
rect 14868 47180 17724 47236
rect 17780 47180 17790 47236
rect 19292 47180 21868 47236
rect 21924 47180 21934 47236
rect 23762 47180 23772 47236
rect 23828 47180 24332 47236
rect 24388 47180 24398 47236
rect 25218 47180 25228 47236
rect 25284 47180 25564 47236
rect 25620 47180 28364 47236
rect 28420 47180 28430 47236
rect 29698 47180 29708 47236
rect 29764 47180 30716 47236
rect 30772 47180 31724 47236
rect 31780 47180 31790 47236
rect 34402 47180 34412 47236
rect 34468 47180 37772 47236
rect 37828 47180 37838 47236
rect 38098 47180 38108 47236
rect 38164 47180 38668 47236
rect 38724 47180 38734 47236
rect 50194 47180 50204 47236
rect 50260 47180 51100 47236
rect 51156 47180 51660 47236
rect 51716 47180 51726 47236
rect 55412 47180 56588 47236
rect 56644 47180 57484 47236
rect 57540 47180 57550 47236
rect 29708 47124 29764 47180
rect 2380 47068 4396 47124
rect 4452 47068 4462 47124
rect 4956 47068 5068 47124
rect 5124 47068 5134 47124
rect 5282 47068 5292 47124
rect 5348 47068 8372 47124
rect 10994 47068 11004 47124
rect 11060 47068 13412 47124
rect 14466 47068 14476 47124
rect 14532 47068 15708 47124
rect 15764 47068 15932 47124
rect 15988 47068 15998 47124
rect 20178 47068 20188 47124
rect 20244 47068 20636 47124
rect 20692 47068 20702 47124
rect 21522 47068 21532 47124
rect 21588 47068 21598 47124
rect 28242 47068 28252 47124
rect 28308 47068 29764 47124
rect 33282 47068 33292 47124
rect 33348 47068 34300 47124
rect 34356 47068 34366 47124
rect 34738 47068 34748 47124
rect 34804 47068 37996 47124
rect 38052 47068 40460 47124
rect 40516 47068 40526 47124
rect 47170 47068 47180 47124
rect 47236 47068 47852 47124
rect 47908 47068 48300 47124
rect 48356 47068 48860 47124
rect 48916 47068 48926 47124
rect 2380 47012 2436 47068
rect 4834 47012 4844 47068
rect 4900 47012 5012 47068
rect 8316 47012 8372 47068
rect 13356 47012 13412 47068
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 21532 47012 21588 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 2370 46956 2380 47012
rect 2436 46956 2446 47012
rect 3938 46956 3948 47012
rect 4004 46956 4620 47012
rect 4676 46956 4686 47012
rect 7522 46956 7532 47012
rect 7588 46956 8092 47012
rect 8148 46956 8158 47012
rect 8316 46956 8764 47012
rect 8820 46956 8830 47012
rect 11554 46956 11564 47012
rect 11620 46956 12236 47012
rect 12292 46956 12302 47012
rect 13356 46956 14364 47012
rect 14420 46956 14430 47012
rect 15026 46956 15036 47012
rect 15092 46956 16828 47012
rect 16884 46956 18060 47012
rect 18116 46956 18126 47012
rect 20402 46956 20412 47012
rect 20468 46956 21588 47012
rect 25900 46956 26236 47012
rect 26292 46956 26302 47012
rect 31266 46956 31276 47012
rect 31332 46956 31612 47012
rect 31668 46956 32620 47012
rect 32676 46956 32686 47012
rect 34962 46956 34972 47012
rect 35028 46956 35644 47012
rect 35700 46956 36540 47012
rect 36596 46956 36606 47012
rect 45266 46956 45276 47012
rect 45332 46956 48636 47012
rect 48692 46956 48702 47012
rect 14364 46900 14420 46956
rect 25900 46900 25956 46956
rect 4834 46844 4844 46900
rect 4900 46844 5404 46900
rect 5460 46844 5470 46900
rect 6066 46844 6076 46900
rect 6132 46844 9884 46900
rect 9940 46844 10612 46900
rect 10966 46844 11004 46900
rect 11060 46844 11070 46900
rect 11218 46844 11228 46900
rect 11284 46844 14140 46900
rect 14196 46844 14206 46900
rect 14364 46844 16156 46900
rect 16212 46844 16222 46900
rect 25554 46844 25564 46900
rect 25620 46844 25676 46900
rect 25732 46844 25742 46900
rect 25890 46844 25900 46900
rect 25956 46844 25966 46900
rect 34290 46844 34300 46900
rect 34356 46844 38444 46900
rect 38500 46844 41804 46900
rect 41860 46844 41870 46900
rect 48514 46844 48524 46900
rect 48580 46844 49980 46900
rect 50036 46844 50046 46900
rect 10556 46788 10612 46844
rect 2146 46732 2156 46788
rect 2212 46732 2940 46788
rect 2996 46732 3500 46788
rect 3556 46732 3566 46788
rect 4722 46732 4732 46788
rect 4788 46732 6412 46788
rect 6468 46732 6478 46788
rect 6626 46732 6636 46788
rect 6692 46732 7644 46788
rect 7700 46732 7710 46788
rect 10546 46732 10556 46788
rect 10612 46732 11340 46788
rect 11396 46732 11788 46788
rect 11844 46732 11854 46788
rect 13122 46732 13132 46788
rect 13188 46732 15316 46788
rect 15810 46732 15820 46788
rect 15876 46732 23100 46788
rect 23156 46732 23166 46788
rect 23314 46732 23324 46788
rect 23380 46732 23772 46788
rect 23828 46732 24892 46788
rect 24948 46732 27860 46788
rect 44706 46732 44716 46788
rect 44772 46732 45500 46788
rect 45556 46732 45566 46788
rect 55458 46732 55468 46788
rect 55524 46732 56476 46788
rect 56532 46732 56542 46788
rect 15260 46676 15316 46732
rect 2818 46620 2828 46676
rect 2884 46620 7028 46676
rect 7186 46620 7196 46676
rect 7252 46620 7868 46676
rect 7924 46620 7934 46676
rect 9090 46620 9100 46676
rect 9156 46620 13916 46676
rect 13972 46620 13982 46676
rect 14242 46620 14252 46676
rect 14308 46620 15036 46676
rect 15092 46620 15102 46676
rect 15250 46620 15260 46676
rect 15316 46620 15354 46676
rect 16566 46620 16604 46676
rect 16660 46620 16670 46676
rect 22082 46620 22092 46676
rect 22148 46620 23548 46676
rect 23604 46620 23614 46676
rect 24434 46620 24444 46676
rect 24500 46620 26236 46676
rect 26292 46620 26302 46676
rect 6972 46564 7028 46620
rect 27804 46564 27860 46732
rect 28130 46620 28140 46676
rect 28196 46620 28924 46676
rect 28980 46620 29932 46676
rect 29988 46620 29998 46676
rect 35746 46620 35756 46676
rect 35812 46620 36876 46676
rect 36932 46620 36942 46676
rect 48738 46620 48748 46676
rect 48804 46620 49532 46676
rect 49588 46620 49598 46676
rect 55234 46620 55244 46676
rect 55300 46620 55468 46676
rect 55412 46564 55468 46620
rect 4162 46508 4172 46564
rect 4228 46508 5068 46564
rect 5124 46508 5852 46564
rect 5908 46508 5918 46564
rect 6972 46508 8204 46564
rect 8260 46508 8764 46564
rect 8820 46508 8830 46564
rect 9762 46508 9772 46564
rect 9828 46508 11676 46564
rect 11732 46508 11742 46564
rect 16370 46508 16380 46564
rect 16436 46508 17836 46564
rect 17892 46508 17902 46564
rect 20402 46508 20412 46564
rect 20468 46508 23436 46564
rect 23492 46508 23502 46564
rect 25666 46508 25676 46564
rect 25732 46508 25788 46564
rect 25844 46508 25854 46564
rect 27794 46508 27804 46564
rect 27860 46508 28700 46564
rect 28756 46508 32172 46564
rect 32228 46508 32238 46564
rect 35858 46508 35868 46564
rect 35924 46508 36988 46564
rect 37044 46508 37054 46564
rect 55412 46508 56476 46564
rect 56532 46508 56924 46564
rect 56980 46508 56990 46564
rect 1810 46396 1820 46452
rect 1876 46396 2604 46452
rect 2660 46396 6972 46452
rect 7028 46396 7038 46452
rect 8866 46396 8876 46452
rect 8932 46396 18620 46452
rect 18676 46396 18686 46452
rect 21634 46396 21644 46452
rect 21700 46396 22540 46452
rect 22596 46396 24220 46452
rect 24276 46396 24892 46452
rect 24948 46396 28140 46452
rect 28196 46396 28206 46452
rect 28466 46396 28476 46452
rect 28532 46396 30828 46452
rect 30884 46396 30894 46452
rect 32246 46396 32284 46452
rect 32340 46396 32350 46452
rect 33964 46396 41132 46452
rect 41188 46396 41198 46452
rect 53442 46396 53452 46452
rect 53508 46396 54012 46452
rect 54068 46396 54078 46452
rect 55570 46396 55580 46452
rect 55636 46396 56028 46452
rect 56084 46396 56094 46452
rect 5618 46284 5628 46340
rect 5684 46284 10780 46340
rect 10836 46284 11452 46340
rect 11508 46284 11732 46340
rect 14130 46284 14140 46340
rect 14196 46284 14588 46340
rect 14644 46284 17948 46340
rect 18004 46284 18014 46340
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 11676 46228 11732 46284
rect 33964 46228 34020 46396
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 3378 46172 3388 46228
rect 3444 46172 3612 46228
rect 3668 46172 3678 46228
rect 6860 46172 8092 46228
rect 8148 46172 8316 46228
rect 8372 46172 8382 46228
rect 8866 46172 8876 46228
rect 8932 46172 9772 46228
rect 9828 46172 9838 46228
rect 11666 46172 11676 46228
rect 11732 46172 11742 46228
rect 12674 46172 12684 46228
rect 12740 46172 14252 46228
rect 14308 46172 14318 46228
rect 15362 46172 15372 46228
rect 15428 46172 18508 46228
rect 18564 46172 18574 46228
rect 25302 46172 25340 46228
rect 25396 46172 25406 46228
rect 26898 46172 26908 46228
rect 26964 46172 27468 46228
rect 27524 46172 28252 46228
rect 28308 46172 28318 46228
rect 28578 46172 28588 46228
rect 28644 46172 33964 46228
rect 34020 46172 34030 46228
rect 55794 46172 55804 46228
rect 55860 46172 56700 46228
rect 56756 46172 56766 46228
rect 6860 46116 6916 46172
rect 1922 46060 1932 46116
rect 1988 46060 6916 46116
rect 7074 46060 7084 46116
rect 7140 46060 12740 46116
rect 17378 46060 17388 46116
rect 17444 46060 17836 46116
rect 17892 46060 17902 46116
rect 24658 46060 24668 46116
rect 24724 46060 26348 46116
rect 26404 46060 26414 46116
rect 29922 46060 29932 46116
rect 29988 46060 32060 46116
rect 32116 46060 32126 46116
rect 32498 46060 32508 46116
rect 32564 46060 33516 46116
rect 33572 46060 36540 46116
rect 36596 46060 36606 46116
rect 37762 46060 37772 46116
rect 37828 46060 37838 46116
rect 38546 46060 38556 46116
rect 38612 46060 39228 46116
rect 39284 46060 39294 46116
rect 12684 46004 12740 46060
rect 32060 46004 32116 46060
rect 37772 46004 37828 46060
rect 2034 45948 2044 46004
rect 2100 45948 3948 46004
rect 4004 45948 7308 46004
rect 7364 45948 7374 46004
rect 7494 45948 7532 46004
rect 7588 45948 7598 46004
rect 8642 45948 8652 46004
rect 8708 45948 8876 46004
rect 8932 45948 12124 46004
rect 12180 45948 12190 46004
rect 12674 45948 12684 46004
rect 12740 45948 19628 46004
rect 19684 45948 19694 46004
rect 24770 45948 24780 46004
rect 24836 45948 25508 46004
rect 26002 45948 26012 46004
rect 26068 45948 26908 46004
rect 26964 45948 26974 46004
rect 28018 45948 28028 46004
rect 28084 45948 29708 46004
rect 29764 45948 29774 46004
rect 30258 45948 30268 46004
rect 30324 45948 31612 46004
rect 31668 45948 31836 46004
rect 31892 45948 31902 46004
rect 32060 45948 33740 46004
rect 33796 45948 34524 46004
rect 34580 45948 34590 46004
rect 36082 45948 36092 46004
rect 36148 45948 37996 46004
rect 38052 45948 38062 46004
rect 38612 45948 39452 46004
rect 39508 45948 39518 46004
rect 56578 45948 56588 46004
rect 56644 45948 57036 46004
rect 57092 45948 57102 46004
rect 12124 45892 12180 45948
rect 25452 45892 25508 45948
rect 4946 45836 4956 45892
rect 5012 45836 5022 45892
rect 6626 45836 6636 45892
rect 6692 45836 7980 45892
rect 8036 45836 9100 45892
rect 9156 45836 9166 45892
rect 12124 45836 12796 45892
rect 12852 45836 14028 45892
rect 14084 45836 14094 45892
rect 16482 45836 16492 45892
rect 16548 45836 17388 45892
rect 17444 45836 20300 45892
rect 20356 45836 20366 45892
rect 25442 45836 25452 45892
rect 25508 45836 25518 45892
rect 4956 45780 5012 45836
rect 28028 45780 28084 45948
rect 38612 45892 38668 45948
rect 31490 45836 31500 45892
rect 31556 45836 36204 45892
rect 36260 45836 36270 45892
rect 36754 45836 36764 45892
rect 36820 45836 37772 45892
rect 37828 45836 37838 45892
rect 37996 45836 38668 45892
rect 42130 45836 42140 45892
rect 42196 45836 42812 45892
rect 42868 45836 42878 45892
rect 45154 45836 45164 45892
rect 45220 45836 45948 45892
rect 46004 45836 46014 45892
rect 52882 45836 52892 45892
rect 52948 45836 53228 45892
rect 53284 45836 53788 45892
rect 53844 45836 53854 45892
rect 4274 45724 4284 45780
rect 4340 45724 4508 45780
rect 4564 45724 4574 45780
rect 4956 45724 6748 45780
rect 6804 45724 8204 45780
rect 8260 45724 8270 45780
rect 11442 45724 11452 45780
rect 11508 45724 13468 45780
rect 13524 45724 13916 45780
rect 13972 45724 14476 45780
rect 14532 45724 14542 45780
rect 16034 45724 16044 45780
rect 16100 45724 21308 45780
rect 21364 45724 21374 45780
rect 24210 45724 24220 45780
rect 24276 45724 25788 45780
rect 25844 45724 25854 45780
rect 26898 45724 26908 45780
rect 26964 45724 28084 45780
rect 28242 45724 28252 45780
rect 28308 45724 29932 45780
rect 29988 45724 29998 45780
rect 33058 45724 33068 45780
rect 33124 45724 37100 45780
rect 37156 45724 37166 45780
rect 37996 45668 38052 45836
rect 3266 45612 3276 45668
rect 3332 45612 6188 45668
rect 6244 45612 6254 45668
rect 6784 45612 6860 45668
rect 6916 45612 7756 45668
rect 7812 45612 7822 45668
rect 8082 45612 8092 45668
rect 8148 45612 11788 45668
rect 11844 45612 13244 45668
rect 13300 45612 13310 45668
rect 16930 45612 16940 45668
rect 16996 45612 21532 45668
rect 21588 45612 22092 45668
rect 22148 45612 22158 45668
rect 23202 45612 23212 45668
rect 23268 45612 25340 45668
rect 25396 45612 25406 45668
rect 25554 45612 25564 45668
rect 25620 45612 25630 45668
rect 28130 45612 28140 45668
rect 28196 45612 28588 45668
rect 28644 45612 30380 45668
rect 30436 45612 30446 45668
rect 32162 45612 32172 45668
rect 32228 45612 32844 45668
rect 32900 45612 32910 45668
rect 33282 45612 33292 45668
rect 33348 45612 35532 45668
rect 35588 45612 35598 45668
rect 35746 45612 35756 45668
rect 35812 45612 36876 45668
rect 36932 45612 38052 45668
rect 38108 45724 38668 45780
rect 38724 45724 40236 45780
rect 40292 45724 40302 45780
rect 41682 45724 41692 45780
rect 41748 45724 42588 45780
rect 42644 45724 43036 45780
rect 43092 45724 43102 45780
rect 44482 45724 44492 45780
rect 44548 45724 45500 45780
rect 45556 45724 45566 45780
rect 8092 45556 8148 45612
rect 24892 45556 24948 45612
rect 3332 45500 4396 45556
rect 4452 45500 6076 45556
rect 6132 45500 6142 45556
rect 6962 45500 6972 45556
rect 7028 45500 7084 45556
rect 7140 45500 8148 45556
rect 13010 45500 13020 45556
rect 13076 45500 13916 45556
rect 13972 45500 13982 45556
rect 20962 45500 20972 45556
rect 21028 45500 22540 45556
rect 22596 45500 22606 45556
rect 23090 45500 23100 45556
rect 23156 45500 23548 45556
rect 23604 45500 24332 45556
rect 24388 45500 24398 45556
rect 24882 45500 24892 45556
rect 24948 45500 24958 45556
rect 3332 45444 3388 45500
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 25564 45444 25620 45612
rect 32844 45556 32900 45612
rect 35532 45556 35588 45612
rect 38108 45556 38164 45724
rect 38434 45612 38444 45668
rect 38500 45612 39564 45668
rect 39620 45612 39630 45668
rect 40562 45612 40572 45668
rect 40628 45612 41132 45668
rect 41188 45612 42476 45668
rect 42532 45612 42542 45668
rect 44146 45612 44156 45668
rect 44212 45612 45108 45668
rect 54226 45612 54236 45668
rect 54292 45612 54908 45668
rect 54964 45612 54974 45668
rect 28802 45500 28812 45556
rect 28868 45500 29596 45556
rect 29652 45500 29662 45556
rect 32844 45500 34860 45556
rect 34916 45500 34926 45556
rect 35532 45500 37100 45556
rect 37156 45500 38164 45556
rect 45052 45444 45108 45612
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 2482 45388 2492 45444
rect 2548 45388 3388 45444
rect 3602 45388 3612 45444
rect 3668 45388 9660 45444
rect 9716 45388 9726 45444
rect 14018 45388 14028 45444
rect 14084 45388 16604 45444
rect 16660 45388 16670 45444
rect 20402 45388 20412 45444
rect 20468 45388 20860 45444
rect 20916 45388 20926 45444
rect 22866 45388 22876 45444
rect 22932 45388 23996 45444
rect 24052 45388 24062 45444
rect 24322 45388 24332 45444
rect 24388 45388 25620 45444
rect 34738 45388 34748 45444
rect 34804 45388 41468 45444
rect 41524 45388 41534 45444
rect 45042 45388 45052 45444
rect 45108 45388 45724 45444
rect 45780 45388 45790 45444
rect 3088 45276 3164 45332
rect 3220 45276 4284 45332
rect 4340 45276 4350 45332
rect 4834 45276 4844 45332
rect 4900 45276 6972 45332
rect 7028 45276 7038 45332
rect 7522 45276 7532 45332
rect 7588 45276 10780 45332
rect 10836 45276 10846 45332
rect 12674 45276 12684 45332
rect 12740 45276 15596 45332
rect 15652 45276 15662 45332
rect 18274 45276 18284 45332
rect 18340 45276 20524 45332
rect 20580 45276 20590 45332
rect 24994 45276 25004 45332
rect 25060 45276 25228 45332
rect 25284 45276 25294 45332
rect 27346 45276 27356 45332
rect 27412 45276 27580 45332
rect 27636 45276 27646 45332
rect 28018 45276 28028 45332
rect 28084 45276 29260 45332
rect 29316 45276 29326 45332
rect 29474 45276 29484 45332
rect 29540 45276 30492 45332
rect 30548 45276 30558 45332
rect 30902 45276 30940 45332
rect 30996 45276 31006 45332
rect 32050 45276 32060 45332
rect 32116 45276 34636 45332
rect 34692 45276 38780 45332
rect 38836 45276 38846 45332
rect 15596 45220 15652 45276
rect 32060 45220 32116 45276
rect 2118 45164 2156 45220
rect 2212 45164 2222 45220
rect 2818 45164 2828 45220
rect 2884 45164 3612 45220
rect 3668 45164 3678 45220
rect 11666 45164 11676 45220
rect 11732 45164 12796 45220
rect 12852 45164 12862 45220
rect 15596 45164 21644 45220
rect 21700 45164 21710 45220
rect 26786 45164 26796 45220
rect 26852 45164 29372 45220
rect 29428 45164 29438 45220
rect 29586 45164 29596 45220
rect 29652 45164 29932 45220
rect 29988 45164 32116 45220
rect 36642 45164 36652 45220
rect 36708 45164 38220 45220
rect 38276 45164 38286 45220
rect 43586 45164 43596 45220
rect 43652 45164 44268 45220
rect 44324 45164 44334 45220
rect 51874 45164 51884 45220
rect 51940 45164 54012 45220
rect 54068 45164 54078 45220
rect 56242 45164 56252 45220
rect 56308 45164 56700 45220
rect 56756 45164 56766 45220
rect 1810 45052 1820 45108
rect 1876 45052 2492 45108
rect 2548 45052 2558 45108
rect 2930 45052 2940 45108
rect 2996 45052 5964 45108
rect 6020 45052 6030 45108
rect 6626 45052 6636 45108
rect 6692 45052 7308 45108
rect 7364 45052 8204 45108
rect 8260 45052 8270 45108
rect 10434 45052 10444 45108
rect 10500 45052 10780 45108
rect 10836 45052 11452 45108
rect 11508 45052 11518 45108
rect 14802 45052 14812 45108
rect 14868 45052 20188 45108
rect 20244 45052 20254 45108
rect 22642 45052 22652 45108
rect 22708 45052 23772 45108
rect 23828 45052 23838 45108
rect 24210 45052 24220 45108
rect 24276 45052 25676 45108
rect 25732 45052 25742 45108
rect 26852 45052 27020 45108
rect 27076 45052 27086 45108
rect 27794 45052 27804 45108
rect 27860 45052 28028 45108
rect 28084 45052 28094 45108
rect 29250 45052 29260 45108
rect 29316 45052 30044 45108
rect 30100 45052 31388 45108
rect 31444 45052 31454 45108
rect 35074 45052 35084 45108
rect 35140 45052 35532 45108
rect 35588 45052 35756 45108
rect 35812 45052 35822 45108
rect 41346 45052 41356 45108
rect 41412 45052 42252 45108
rect 42308 45052 42318 45108
rect 46722 45052 46732 45108
rect 46788 45052 47068 45108
rect 47124 45052 47740 45108
rect 47796 45052 47806 45108
rect 48738 45052 48748 45108
rect 48804 45052 49868 45108
rect 49924 45052 49934 45108
rect 52098 45052 52108 45108
rect 52164 45052 53340 45108
rect 53396 45052 53406 45108
rect 57810 45052 57820 45108
rect 57876 45052 58492 45108
rect 58548 45052 58558 45108
rect 2940 44996 2996 45052
rect 26852 44996 26908 45052
rect 2370 44940 2380 44996
rect 2436 44940 2996 44996
rect 4498 44940 4508 44996
rect 4564 44940 4844 44996
rect 4900 44940 5068 44996
rect 5124 44940 6412 44996
rect 6468 44940 6478 44996
rect 9650 44940 9660 44996
rect 9716 44940 10332 44996
rect 10388 44940 11564 44996
rect 11620 44940 11630 44996
rect 16370 44940 16380 44996
rect 16436 44940 16492 44996
rect 16548 44940 16558 44996
rect 23874 44940 23884 44996
rect 23940 44940 30156 44996
rect 30212 44940 30940 44996
rect 30996 44940 31006 44996
rect 32498 44940 32508 44996
rect 32564 44940 32956 44996
rect 33012 44940 33628 44996
rect 33684 44940 33694 44996
rect 34850 44940 34860 44996
rect 34916 44940 35980 44996
rect 36036 44940 37548 44996
rect 37604 44940 40348 44996
rect 40404 44940 40414 44996
rect 48514 44940 48524 44996
rect 48580 44940 49084 44996
rect 49140 44940 49644 44996
rect 49700 44940 49710 44996
rect 50530 44940 50540 44996
rect 50596 44940 51100 44996
rect 51156 44940 51548 44996
rect 51604 44940 51614 44996
rect 4050 44828 4060 44884
rect 4116 44828 9212 44884
rect 9268 44828 11900 44884
rect 11956 44828 12348 44884
rect 12404 44828 12572 44884
rect 12628 44828 12638 44884
rect 18610 44828 18620 44884
rect 18676 44828 22204 44884
rect 22260 44828 22270 44884
rect 23650 44828 23660 44884
rect 23716 44828 24332 44884
rect 24388 44828 26012 44884
rect 26068 44828 28700 44884
rect 28756 44828 28766 44884
rect 50866 44828 50876 44884
rect 50932 44828 51996 44884
rect 52052 44828 53788 44884
rect 53844 44828 53854 44884
rect 4834 44716 4844 44772
rect 4900 44716 6076 44772
rect 6132 44716 8540 44772
rect 8596 44716 8606 44772
rect 16146 44716 16156 44772
rect 16212 44716 19292 44772
rect 19348 44716 21308 44772
rect 21364 44716 21374 44772
rect 24994 44716 25004 44772
rect 25060 44716 27244 44772
rect 27300 44716 27310 44772
rect 27542 44716 27580 44772
rect 27636 44716 27646 44772
rect 28018 44716 28028 44772
rect 28084 44716 34412 44772
rect 34468 44716 34478 44772
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 7046 44604 7084 44660
rect 7140 44604 7150 44660
rect 10098 44604 10108 44660
rect 10164 44604 14364 44660
rect 14420 44604 14430 44660
rect 17490 44604 17500 44660
rect 17556 44604 22092 44660
rect 22148 44604 24220 44660
rect 24276 44604 24286 44660
rect 25218 44604 25228 44660
rect 25284 44604 25788 44660
rect 25844 44604 26348 44660
rect 26404 44604 26414 44660
rect 40562 44604 40572 44660
rect 40628 44604 47180 44660
rect 47236 44604 47246 44660
rect 10108 44548 10164 44604
rect 3378 44492 3388 44548
rect 3444 44492 4396 44548
rect 4452 44492 10164 44548
rect 13794 44492 13804 44548
rect 13860 44492 16156 44548
rect 16212 44492 16222 44548
rect 20178 44492 20188 44548
rect 20244 44492 21756 44548
rect 21812 44492 21822 44548
rect 24658 44492 24668 44548
rect 24724 44492 25676 44548
rect 25732 44492 25742 44548
rect 45714 44492 45724 44548
rect 45780 44492 46228 44548
rect 55010 44492 55020 44548
rect 55076 44492 56700 44548
rect 56756 44492 56766 44548
rect 46172 44436 46228 44492
rect 3332 44380 4284 44436
rect 4340 44380 8428 44436
rect 8484 44380 8494 44436
rect 8642 44380 8652 44436
rect 8708 44380 8718 44436
rect 10210 44380 10220 44436
rect 10276 44380 17948 44436
rect 18004 44380 18014 44436
rect 19282 44380 19292 44436
rect 19348 44380 19740 44436
rect 19796 44380 20300 44436
rect 20356 44380 20366 44436
rect 23538 44380 23548 44436
rect 23604 44380 27916 44436
rect 27972 44380 27982 44436
rect 30370 44380 30380 44436
rect 30436 44380 30716 44436
rect 30772 44380 30782 44436
rect 38770 44380 38780 44436
rect 38836 44380 39676 44436
rect 39732 44380 39900 44436
rect 39956 44380 39966 44436
rect 40226 44380 40236 44436
rect 40292 44380 41356 44436
rect 41412 44380 41422 44436
rect 44258 44380 44268 44436
rect 44324 44380 45836 44436
rect 45892 44380 45902 44436
rect 46162 44380 46172 44436
rect 46228 44380 57708 44436
rect 57764 44380 57774 44436
rect 3332 44324 3388 44380
rect 2706 44268 2716 44324
rect 2772 44268 3052 44324
rect 3108 44268 3388 44324
rect 5926 44268 5964 44324
rect 6020 44268 6030 44324
rect 8652 44212 8708 44380
rect 10322 44268 10332 44324
rect 10388 44268 11564 44324
rect 11620 44268 12012 44324
rect 12068 44268 12078 44324
rect 12226 44268 12236 44324
rect 12292 44268 15820 44324
rect 15876 44268 15886 44324
rect 18274 44268 18284 44324
rect 18340 44268 19068 44324
rect 19124 44268 20748 44324
rect 20804 44268 22092 44324
rect 22148 44268 22158 44324
rect 22306 44268 22316 44324
rect 22372 44268 22988 44324
rect 23044 44268 23054 44324
rect 26450 44268 26460 44324
rect 26516 44268 27468 44324
rect 27524 44268 27534 44324
rect 40002 44268 40012 44324
rect 40068 44268 41244 44324
rect 41300 44268 41310 44324
rect 41570 44268 41580 44324
rect 41636 44268 42588 44324
rect 42644 44268 42924 44324
rect 42980 44268 42990 44324
rect 48178 44268 48188 44324
rect 48244 44268 50092 44324
rect 50148 44268 50158 44324
rect 2146 44156 2156 44212
rect 2212 44156 4956 44212
rect 5012 44156 9436 44212
rect 9492 44156 9502 44212
rect 9650 44156 9660 44212
rect 9716 44156 10220 44212
rect 10276 44156 10286 44212
rect 10434 44156 10444 44212
rect 10500 44156 11116 44212
rect 11172 44156 11182 44212
rect 13122 44156 13132 44212
rect 13188 44156 14924 44212
rect 14980 44156 19180 44212
rect 19236 44156 19246 44212
rect 21746 44156 21756 44212
rect 21812 44156 22092 44212
rect 22148 44156 22204 44212
rect 22260 44156 22270 44212
rect 23202 44156 23212 44212
rect 23268 44156 26348 44212
rect 26404 44156 28924 44212
rect 28980 44156 29484 44212
rect 29540 44156 34748 44212
rect 34804 44156 35756 44212
rect 35812 44156 35822 44212
rect 38098 44156 38108 44212
rect 38164 44156 39676 44212
rect 39732 44156 39742 44212
rect 43474 44156 43484 44212
rect 43540 44156 48300 44212
rect 48356 44156 49644 44212
rect 49700 44156 49710 44212
rect 52098 44156 52108 44212
rect 52164 44156 53900 44212
rect 53956 44156 53966 44212
rect 2930 44044 2940 44100
rect 2996 44044 3052 44100
rect 3108 44044 3118 44100
rect 3714 44044 3724 44100
rect 3780 44044 5180 44100
rect 5236 44044 7196 44100
rect 7252 44044 7262 44100
rect 8530 44044 8540 44100
rect 8596 44044 9660 44100
rect 9716 44044 12684 44100
rect 12740 44044 12750 44100
rect 13346 44044 13356 44100
rect 13412 44044 13804 44100
rect 13860 44044 13870 44100
rect 14354 44044 14364 44100
rect 14420 44044 15708 44100
rect 15764 44044 15774 44100
rect 15932 43988 15988 44156
rect 16370 44044 16380 44100
rect 16436 44044 17052 44100
rect 17108 44044 17118 44100
rect 17266 44044 17276 44100
rect 17332 44044 17500 44100
rect 17556 44044 19516 44100
rect 19572 44044 19582 44100
rect 23510 44044 23548 44100
rect 23604 44044 23614 44100
rect 23762 44044 23772 44100
rect 23828 44044 23884 44100
rect 23940 44044 23950 44100
rect 31378 44044 31388 44100
rect 31444 44044 34860 44100
rect 34916 44044 34926 44100
rect 36306 44044 36316 44100
rect 36372 44044 39564 44100
rect 39620 44044 39630 44100
rect 44594 44044 44604 44100
rect 44660 44044 48412 44100
rect 48468 44044 49868 44100
rect 49924 44044 49934 44100
rect 1922 43932 1932 43988
rect 1988 43932 3500 43988
rect 3556 43932 5740 43988
rect 5796 43932 5806 43988
rect 6402 43932 6412 43988
rect 6468 43932 12348 43988
rect 12404 43932 12414 43988
rect 15810 43932 15820 43988
rect 15876 43932 15988 43988
rect 23762 43932 23772 43988
rect 23828 43932 24780 43988
rect 24836 43932 24846 43988
rect 25004 43932 28028 43988
rect 28084 43932 28094 43988
rect 28242 43932 28252 43988
rect 28308 43932 30828 43988
rect 30884 43932 33180 43988
rect 33236 43932 33246 43988
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 25004 43876 25060 43932
rect 28252 43876 28308 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 7858 43820 7868 43876
rect 7924 43820 8540 43876
rect 8596 43820 8606 43876
rect 8866 43820 8876 43876
rect 8932 43820 11788 43876
rect 11844 43820 13020 43876
rect 13076 43820 13086 43876
rect 16818 43820 16828 43876
rect 16884 43820 17052 43876
rect 17108 43820 18060 43876
rect 18116 43820 18126 43876
rect 23996 43820 25060 43876
rect 25330 43820 25340 43876
rect 25396 43820 26012 43876
rect 26068 43820 26460 43876
rect 26516 43820 26526 43876
rect 26852 43820 27132 43876
rect 27188 43820 28308 43876
rect 23996 43764 24052 43820
rect 26852 43764 26908 43820
rect 3378 43708 3388 43764
rect 3444 43708 5124 43764
rect 6514 43708 6524 43764
rect 6580 43708 7868 43764
rect 7924 43708 7934 43764
rect 10210 43708 10220 43764
rect 10276 43708 10332 43764
rect 10388 43708 10398 43764
rect 11554 43708 11564 43764
rect 11620 43708 13580 43764
rect 13636 43708 13646 43764
rect 14690 43708 14700 43764
rect 14756 43708 20412 43764
rect 20468 43708 20478 43764
rect 22754 43708 22764 43764
rect 22820 43708 23996 43764
rect 24052 43708 24062 43764
rect 25106 43708 25116 43764
rect 25172 43708 26908 43764
rect 27010 43708 27020 43764
rect 27076 43708 28140 43764
rect 28196 43708 29036 43764
rect 29092 43708 29102 43764
rect 37538 43708 37548 43764
rect 37604 43708 38220 43764
rect 38276 43708 38286 43764
rect 43586 43708 43596 43764
rect 43652 43708 43662 43764
rect 56578 43708 56588 43764
rect 56644 43708 57484 43764
rect 57540 43708 57550 43764
rect 3042 43596 3052 43652
rect 3108 43596 4844 43652
rect 4900 43596 4910 43652
rect 5068 43540 5124 43708
rect 43596 43652 43652 43708
rect 5282 43596 5292 43652
rect 5348 43596 7084 43652
rect 7140 43596 7150 43652
rect 7858 43596 7868 43652
rect 7924 43596 8764 43652
rect 8820 43596 8830 43652
rect 9734 43596 9772 43652
rect 9828 43596 9838 43652
rect 10098 43596 10108 43652
rect 10164 43596 10444 43652
rect 10500 43596 11228 43652
rect 11284 43596 11294 43652
rect 11414 43596 11452 43652
rect 11508 43596 11518 43652
rect 15250 43596 15260 43652
rect 15316 43596 16268 43652
rect 16324 43596 16334 43652
rect 18806 43596 18844 43652
rect 18900 43596 18910 43652
rect 19394 43596 19404 43652
rect 19460 43596 21196 43652
rect 21252 43596 21262 43652
rect 26898 43596 26908 43652
rect 26964 43596 28476 43652
rect 28532 43596 28542 43652
rect 32162 43596 32172 43652
rect 32228 43596 35308 43652
rect 35364 43596 35374 43652
rect 36194 43596 36204 43652
rect 36260 43596 37884 43652
rect 37940 43596 37950 43652
rect 39666 43596 39676 43652
rect 39732 43596 40348 43652
rect 40404 43596 43652 43652
rect 44706 43596 44716 43652
rect 44772 43596 45276 43652
rect 45332 43596 45342 43652
rect 5068 43484 5180 43540
rect 5236 43484 6748 43540
rect 6804 43484 7420 43540
rect 7476 43484 7486 43540
rect 7634 43484 7644 43540
rect 7700 43484 12740 43540
rect 12898 43484 12908 43540
rect 12964 43484 13244 43540
rect 13300 43484 13356 43540
rect 13412 43484 13422 43540
rect 13580 43484 14252 43540
rect 14308 43484 15148 43540
rect 16258 43484 16268 43540
rect 16324 43484 16380 43540
rect 16436 43484 16446 43540
rect 17266 43484 17276 43540
rect 17332 43484 17948 43540
rect 18004 43484 18956 43540
rect 19012 43484 19022 43540
rect 19618 43484 19628 43540
rect 19684 43484 20300 43540
rect 20356 43484 20366 43540
rect 21298 43484 21308 43540
rect 21364 43484 21644 43540
rect 21700 43484 21980 43540
rect 22036 43484 22046 43540
rect 24546 43484 24556 43540
rect 24612 43484 27356 43540
rect 27412 43484 27916 43540
rect 27972 43484 27982 43540
rect 31154 43484 31164 43540
rect 31220 43484 34076 43540
rect 34132 43484 35084 43540
rect 35140 43484 35980 43540
rect 36036 43484 37324 43540
rect 37380 43484 37390 43540
rect 40562 43484 40572 43540
rect 40628 43484 41580 43540
rect 41636 43484 41646 43540
rect 42242 43484 42252 43540
rect 42308 43484 43932 43540
rect 43988 43484 43998 43540
rect 56466 43484 56476 43540
rect 56532 43484 56812 43540
rect 56868 43484 57260 43540
rect 57316 43484 57326 43540
rect 12684 43428 12740 43484
rect 13580 43428 13636 43484
rect 15092 43428 15148 43484
rect 3154 43372 3164 43428
rect 3220 43372 6300 43428
rect 6356 43372 6366 43428
rect 8642 43372 8652 43428
rect 8708 43372 8988 43428
rect 9044 43372 9054 43428
rect 12684 43372 13020 43428
rect 13076 43372 13580 43428
rect 13636 43372 13646 43428
rect 13906 43372 13916 43428
rect 13972 43372 14812 43428
rect 14868 43372 14878 43428
rect 15092 43372 18732 43428
rect 18788 43372 18798 43428
rect 21074 43372 21084 43428
rect 21140 43372 24108 43428
rect 24164 43372 24174 43428
rect 25442 43372 25452 43428
rect 25508 43372 25564 43428
rect 25620 43372 26796 43428
rect 26852 43372 27020 43428
rect 27076 43372 27086 43428
rect 27234 43372 27244 43428
rect 27300 43372 31948 43428
rect 32004 43372 32014 43428
rect 32946 43372 32956 43428
rect 33012 43372 33516 43428
rect 33572 43372 33582 43428
rect 40450 43372 40460 43428
rect 40516 43372 40796 43428
rect 40852 43372 45836 43428
rect 45892 43372 46956 43428
rect 47012 43372 47628 43428
rect 47684 43372 47852 43428
rect 47908 43372 47918 43428
rect 27244 43316 27300 43372
rect 1026 43260 1036 43316
rect 1092 43260 3836 43316
rect 3892 43260 4060 43316
rect 4116 43260 10220 43316
rect 10276 43260 13020 43316
rect 13076 43260 13086 43316
rect 15026 43260 15036 43316
rect 15092 43260 15484 43316
rect 15540 43260 15550 43316
rect 16146 43260 16156 43316
rect 16212 43260 16380 43316
rect 16436 43260 17276 43316
rect 17332 43260 19180 43316
rect 19236 43260 20524 43316
rect 20580 43260 21420 43316
rect 21476 43260 21486 43316
rect 25554 43260 25564 43316
rect 25620 43260 27300 43316
rect 31266 43260 31276 43316
rect 31332 43260 32508 43316
rect 32564 43260 32574 43316
rect 32834 43260 32844 43316
rect 32900 43260 34188 43316
rect 34244 43260 34254 43316
rect 41794 43260 41804 43316
rect 41860 43260 46060 43316
rect 46116 43260 46732 43316
rect 46788 43260 46798 43316
rect 32508 43204 32564 43260
rect 2482 43148 2492 43204
rect 2548 43148 3276 43204
rect 3332 43148 3342 43204
rect 9090 43148 9100 43204
rect 9156 43148 11900 43204
rect 11956 43148 11966 43204
rect 23090 43148 23100 43204
rect 23156 43148 26684 43204
rect 26740 43148 26750 43204
rect 32508 43148 33852 43204
rect 33908 43148 33918 43204
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 8082 43036 8092 43092
rect 8148 43036 8764 43092
rect 8820 43036 8830 43092
rect 15138 43036 15148 43092
rect 15204 43036 15372 43092
rect 15428 43036 15438 43092
rect 15698 43036 15708 43092
rect 15764 43036 16156 43092
rect 16212 43036 16222 43092
rect 25666 43036 25676 43092
rect 25732 43036 26236 43092
rect 26292 43036 30492 43092
rect 30548 43036 30558 43092
rect 12114 42924 12124 42980
rect 12180 42924 13468 42980
rect 13524 42924 13534 42980
rect 13692 42924 17612 42980
rect 17668 42924 17678 42980
rect 18946 42924 18956 42980
rect 19012 42924 19068 42980
rect 19124 42924 19628 42980
rect 19684 42924 19694 42980
rect 26684 42924 33292 42980
rect 33348 42924 33358 42980
rect 55794 42924 55804 42980
rect 55860 42924 56476 42980
rect 56532 42924 56542 42980
rect 13692 42868 13748 42924
rect 26684 42868 26740 42924
rect 1362 42812 1372 42868
rect 1428 42812 2604 42868
rect 2660 42812 2670 42868
rect 2902 42812 2940 42868
rect 2996 42812 3006 42868
rect 6402 42812 6412 42868
rect 6468 42812 6636 42868
rect 6692 42812 6702 42868
rect 6850 42812 6860 42868
rect 6916 42812 6972 42868
rect 7028 42812 7038 42868
rect 7746 42812 7756 42868
rect 7812 42812 8428 42868
rect 8484 42812 9660 42868
rect 9716 42812 11228 42868
rect 11284 42812 11294 42868
rect 12338 42812 12348 42868
rect 12404 42812 13748 42868
rect 13878 42812 13916 42868
rect 13972 42812 13982 42868
rect 14242 42812 14252 42868
rect 14308 42812 18396 42868
rect 18452 42812 18462 42868
rect 19478 42812 19516 42868
rect 19572 42812 19582 42868
rect 22754 42812 22764 42868
rect 22820 42812 25116 42868
rect 25172 42812 25340 42868
rect 25396 42812 26684 42868
rect 26740 42812 26750 42868
rect 27010 42812 27020 42868
rect 27076 42812 27916 42868
rect 27972 42812 27982 42868
rect 51762 42812 51772 42868
rect 51828 42812 53900 42868
rect 53956 42812 53966 42868
rect 4022 42700 4060 42756
rect 4116 42700 4126 42756
rect 6066 42700 6076 42756
rect 6132 42700 8540 42756
rect 8596 42700 8606 42756
rect 8950 42700 8988 42756
rect 9044 42700 9054 42756
rect 9202 42700 9212 42756
rect 9268 42700 10668 42756
rect 10724 42700 14364 42756
rect 14420 42700 14430 42756
rect 18722 42700 18732 42756
rect 18788 42700 22204 42756
rect 22260 42700 22270 42756
rect 22418 42700 22428 42756
rect 22484 42700 23660 42756
rect 23716 42700 23726 42756
rect 26758 42700 26796 42756
rect 26852 42700 26862 42756
rect 28802 42700 28812 42756
rect 28868 42700 30492 42756
rect 30548 42700 31500 42756
rect 31556 42700 31948 42756
rect 32004 42700 32014 42756
rect 36194 42700 36204 42756
rect 36260 42700 36652 42756
rect 36708 42700 36718 42756
rect 47394 42700 47404 42756
rect 47460 42700 48188 42756
rect 48244 42700 48254 42756
rect 4274 42588 4284 42644
rect 4340 42588 9884 42644
rect 9940 42588 9950 42644
rect 11554 42588 11564 42644
rect 11620 42588 11788 42644
rect 11844 42588 12348 42644
rect 12404 42588 12414 42644
rect 13346 42588 13356 42644
rect 13412 42588 14140 42644
rect 14196 42588 14206 42644
rect 16034 42588 16044 42644
rect 16100 42588 16492 42644
rect 16548 42588 17388 42644
rect 17444 42588 17454 42644
rect 19954 42588 19964 42644
rect 20020 42588 22092 42644
rect 22148 42588 22316 42644
rect 22372 42588 22382 42644
rect 23090 42588 23100 42644
rect 23156 42588 24892 42644
rect 24948 42588 26124 42644
rect 26180 42588 37996 42644
rect 38052 42588 38062 42644
rect 39778 42588 39788 42644
rect 39844 42588 40348 42644
rect 40404 42588 40414 42644
rect 54898 42588 54908 42644
rect 54964 42588 55468 42644
rect 3714 42476 3724 42532
rect 3780 42476 6300 42532
rect 6356 42476 6636 42532
rect 6692 42476 6702 42532
rect 10322 42476 10332 42532
rect 10388 42476 15148 42532
rect 15922 42476 15932 42532
rect 15988 42476 16380 42532
rect 16436 42476 16446 42532
rect 16594 42476 16604 42532
rect 16660 42476 17948 42532
rect 18004 42476 18014 42532
rect 18274 42476 18284 42532
rect 18340 42476 18620 42532
rect 18676 42476 18686 42532
rect 19618 42476 19628 42532
rect 19684 42476 25788 42532
rect 25844 42476 25854 42532
rect 26450 42476 26460 42532
rect 26516 42476 28028 42532
rect 28084 42476 28094 42532
rect 36418 42476 36428 42532
rect 36484 42476 38444 42532
rect 38500 42476 38510 42532
rect 40786 42476 40796 42532
rect 40852 42476 41356 42532
rect 41412 42476 41422 42532
rect 41794 42476 41804 42532
rect 41860 42476 42364 42532
rect 42420 42476 42430 42532
rect 44706 42476 44716 42532
rect 44772 42476 45836 42532
rect 45892 42476 45902 42532
rect 48402 42476 48412 42532
rect 48468 42476 49084 42532
rect 49140 42476 49532 42532
rect 49588 42476 49598 42532
rect 55412 42476 55468 42588
rect 55524 42476 55916 42532
rect 55972 42476 55982 42532
rect 56130 42476 56140 42532
rect 56196 42476 56364 42532
rect 56420 42476 56430 42532
rect 15092 42420 15148 42476
rect 3490 42364 3500 42420
rect 3556 42364 3948 42420
rect 4004 42364 5740 42420
rect 5796 42364 5806 42420
rect 10658 42364 10668 42420
rect 10724 42364 11564 42420
rect 11620 42364 11630 42420
rect 15092 42364 16604 42420
rect 16660 42364 16670 42420
rect 18162 42364 18172 42420
rect 18228 42364 18396 42420
rect 18452 42364 18462 42420
rect 19170 42364 19180 42420
rect 19236 42364 19516 42420
rect 19572 42364 19582 42420
rect 20402 42364 20412 42420
rect 20468 42364 23660 42420
rect 23716 42364 23726 42420
rect 35522 42364 35532 42420
rect 35588 42364 37548 42420
rect 37604 42364 37614 42420
rect 42130 42364 42140 42420
rect 42196 42364 42476 42420
rect 42532 42364 42700 42420
rect 42756 42364 42766 42420
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 6514 42252 6524 42308
rect 6580 42252 8428 42308
rect 8484 42252 8494 42308
rect 8754 42252 8764 42308
rect 8820 42252 9324 42308
rect 9380 42252 9390 42308
rect 13458 42252 13468 42308
rect 13524 42252 15596 42308
rect 15652 42252 15662 42308
rect 16258 42252 16268 42308
rect 16324 42252 18844 42308
rect 18900 42252 19404 42308
rect 19460 42252 19470 42308
rect 20822 42252 20860 42308
rect 20916 42252 25676 42308
rect 25732 42252 25900 42308
rect 25956 42252 25966 42308
rect 34178 42252 34188 42308
rect 34244 42252 37660 42308
rect 37716 42252 37726 42308
rect 3686 42140 3724 42196
rect 3780 42140 3790 42196
rect 5170 42140 5180 42196
rect 5236 42140 6300 42196
rect 6356 42140 13244 42196
rect 13300 42140 13310 42196
rect 13458 42140 13468 42196
rect 13524 42140 14140 42196
rect 14196 42140 14206 42196
rect 14914 42140 14924 42196
rect 14980 42140 21644 42196
rect 21700 42140 21710 42196
rect 21970 42140 21980 42196
rect 22036 42140 22316 42196
rect 22372 42140 22382 42196
rect 27458 42140 27468 42196
rect 27524 42140 28532 42196
rect 30258 42140 30268 42196
rect 30324 42140 30828 42196
rect 30884 42140 30894 42196
rect 37426 42140 37436 42196
rect 37492 42140 42252 42196
rect 42308 42140 42318 42196
rect 55906 42140 55916 42196
rect 55972 42140 56700 42196
rect 56756 42140 56766 42196
rect 28476 42084 28532 42140
rect 2454 42028 2492 42084
rect 2548 42028 2558 42084
rect 4610 42028 4620 42084
rect 4676 42028 8204 42084
rect 8260 42028 8270 42084
rect 8866 42028 8876 42084
rect 8932 42028 10892 42084
rect 10948 42028 10958 42084
rect 11218 42028 11228 42084
rect 11284 42028 13692 42084
rect 13748 42028 14868 42084
rect 17826 42028 17836 42084
rect 17892 42028 21868 42084
rect 21924 42028 21934 42084
rect 24098 42028 24108 42084
rect 24164 42028 24668 42084
rect 24724 42028 24734 42084
rect 28466 42028 28476 42084
rect 28532 42028 29260 42084
rect 29316 42028 31164 42084
rect 31220 42028 34412 42084
rect 34468 42028 34478 42084
rect 36530 42028 36540 42084
rect 36596 42028 37884 42084
rect 37940 42028 37950 42084
rect 43148 42028 43652 42084
rect 46386 42028 46396 42084
rect 46452 42028 46732 42084
rect 46788 42028 53564 42084
rect 53620 42028 53630 42084
rect 53788 42028 54684 42084
rect 54740 42028 54750 42084
rect 56354 42028 56364 42084
rect 56420 42028 57484 42084
rect 57540 42028 57550 42084
rect 4162 41916 4172 41972
rect 4228 41916 5628 41972
rect 5684 41916 5694 41972
rect 6178 41916 6188 41972
rect 6244 41916 6636 41972
rect 6692 41916 6702 41972
rect 7382 41916 7420 41972
rect 7476 41916 7486 41972
rect 11442 41916 11452 41972
rect 11508 41916 12124 41972
rect 12180 41916 12190 41972
rect 13010 41916 13020 41972
rect 13076 41916 14588 41972
rect 14644 41916 14654 41972
rect 14812 41860 14868 42028
rect 43148 41972 43204 42028
rect 43596 41972 43652 42028
rect 15586 41916 15596 41972
rect 15652 41916 21084 41972
rect 21140 41916 21150 41972
rect 22418 41916 22428 41972
rect 22484 41916 24220 41972
rect 24276 41916 24286 41972
rect 28018 41916 28028 41972
rect 28084 41916 29036 41972
rect 29092 41916 29102 41972
rect 34514 41916 34524 41972
rect 34580 41916 35868 41972
rect 35924 41916 37324 41972
rect 37380 41916 37390 41972
rect 38658 41916 38668 41972
rect 38724 41916 38892 41972
rect 38948 41916 38958 41972
rect 40898 41916 40908 41972
rect 40964 41916 43204 41972
rect 43362 41916 43372 41972
rect 43428 41916 43438 41972
rect 43596 41916 45724 41972
rect 45780 41916 46172 41972
rect 46228 41916 46238 41972
rect 47842 41916 47852 41972
rect 47908 41916 48636 41972
rect 48692 41916 51100 41972
rect 51156 41916 51166 41972
rect 52210 41916 52220 41972
rect 52276 41916 52668 41972
rect 52724 41916 53452 41972
rect 53508 41916 53518 41972
rect 43372 41860 43428 41916
rect 53788 41860 53844 42028
rect 1922 41804 1932 41860
rect 1988 41804 2940 41860
rect 2996 41804 4956 41860
rect 5012 41804 5022 41860
rect 5506 41804 5516 41860
rect 5572 41804 5740 41860
rect 5796 41804 5806 41860
rect 6514 41804 6524 41860
rect 6580 41804 6972 41860
rect 7028 41804 8876 41860
rect 8932 41804 14364 41860
rect 14420 41804 14430 41860
rect 14812 41804 17276 41860
rect 17332 41804 17612 41860
rect 17668 41804 17678 41860
rect 17798 41804 17836 41860
rect 17892 41804 17902 41860
rect 19618 41804 19628 41860
rect 19684 41804 19740 41860
rect 19796 41804 19806 41860
rect 23762 41804 23772 41860
rect 23828 41804 25228 41860
rect 25284 41804 25294 41860
rect 29474 41804 29484 41860
rect 29540 41804 31724 41860
rect 31780 41804 32508 41860
rect 32564 41804 32574 41860
rect 39106 41804 39116 41860
rect 39172 41804 39676 41860
rect 39732 41804 43148 41860
rect 43204 41804 43214 41860
rect 43372 41804 43820 41860
rect 43876 41804 43886 41860
rect 47618 41804 47628 41860
rect 47684 41804 48300 41860
rect 48356 41804 49756 41860
rect 49812 41804 49822 41860
rect 53778 41804 53788 41860
rect 53844 41804 53854 41860
rect 5954 41692 5964 41748
rect 6020 41692 15036 41748
rect 15092 41692 15148 41748
rect 15204 41692 15484 41748
rect 15540 41692 15550 41748
rect 16044 41692 16380 41748
rect 16436 41692 18732 41748
rect 18788 41692 19292 41748
rect 19348 41692 19358 41748
rect 20514 41692 20524 41748
rect 20580 41692 21980 41748
rect 22036 41692 22046 41748
rect 24546 41692 24556 41748
rect 24612 41692 26684 41748
rect 26740 41692 26750 41748
rect 32274 41692 32284 41748
rect 32340 41692 33516 41748
rect 33572 41692 33582 41748
rect 34300 41692 36876 41748
rect 36932 41692 36942 41748
rect 43652 41692 45276 41748
rect 45332 41692 45612 41748
rect 45668 41692 45678 41748
rect 53218 41692 53228 41748
rect 53284 41692 54348 41748
rect 54404 41692 54572 41748
rect 54628 41692 54638 41748
rect 16044 41636 16100 41692
rect 34300 41636 34356 41692
rect 43652 41636 43708 41692
rect 1698 41580 1708 41636
rect 1764 41580 3612 41636
rect 3668 41580 3678 41636
rect 5058 41580 5068 41636
rect 5124 41580 8932 41636
rect 9090 41580 9100 41636
rect 9156 41580 9996 41636
rect 10052 41580 10062 41636
rect 12450 41580 12460 41636
rect 12516 41580 15260 41636
rect 15316 41580 15326 41636
rect 15586 41580 15596 41636
rect 15652 41580 16044 41636
rect 16100 41580 16110 41636
rect 16930 41580 16940 41636
rect 16996 41580 19628 41636
rect 19684 41580 19694 41636
rect 23426 41580 23436 41636
rect 23492 41580 24444 41636
rect 24500 41580 24510 41636
rect 30930 41580 30940 41636
rect 30996 41580 34300 41636
rect 34356 41580 34366 41636
rect 37986 41580 37996 41636
rect 38052 41580 43708 41636
rect 52434 41580 52444 41636
rect 52500 41580 53900 41636
rect 53956 41580 53966 41636
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 8876 41412 8932 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 10098 41468 10108 41524
rect 10164 41468 12684 41524
rect 12740 41468 12750 41524
rect 12944 41468 13020 41524
rect 13076 41468 19068 41524
rect 19124 41468 19292 41524
rect 19348 41468 19358 41524
rect 22866 41468 22876 41524
rect 22932 41468 22942 41524
rect 27916 41468 28364 41524
rect 28420 41468 28430 41524
rect 39778 41468 39788 41524
rect 39844 41468 42028 41524
rect 42084 41468 43260 41524
rect 43316 41468 43326 41524
rect 53442 41468 53452 41524
rect 53508 41468 54236 41524
rect 54292 41468 54302 41524
rect 3602 41356 3612 41412
rect 3668 41356 4844 41412
rect 4900 41356 5852 41412
rect 5908 41356 5918 41412
rect 8876 41356 11788 41412
rect 15250 41356 15260 41412
rect 15316 41356 17724 41412
rect 17780 41356 17790 41412
rect 19366 41356 19404 41412
rect 19460 41356 19470 41412
rect 3490 41244 3500 41300
rect 3556 41244 3836 41300
rect 3892 41244 9548 41300
rect 9604 41244 9614 41300
rect 11732 41188 11788 41356
rect 12898 41244 12908 41300
rect 12964 41244 13356 41300
rect 13412 41244 18620 41300
rect 18676 41244 19180 41300
rect 19236 41244 20748 41300
rect 20804 41244 20814 41300
rect 3154 41132 3164 41188
rect 3220 41132 4060 41188
rect 4116 41132 4508 41188
rect 4564 41132 4574 41188
rect 5618 41132 5628 41188
rect 5684 41132 7420 41188
rect 7476 41132 7486 41188
rect 9212 41132 10668 41188
rect 10724 41132 11116 41188
rect 11172 41132 11182 41188
rect 11732 41132 13468 41188
rect 13524 41132 14140 41188
rect 14196 41132 15036 41188
rect 15092 41132 18060 41188
rect 18116 41132 18126 41188
rect 19058 41132 19068 41188
rect 19124 41132 21532 41188
rect 21588 41132 21756 41188
rect 21812 41132 21822 41188
rect 5628 41076 5684 41132
rect 9212 41076 9268 41132
rect 22876 41076 22932 41468
rect 27916 41412 27972 41468
rect 25004 41356 27020 41412
rect 27076 41356 27916 41412
rect 27972 41356 27982 41412
rect 28242 41356 28252 41412
rect 28308 41356 28924 41412
rect 28980 41356 28990 41412
rect 34514 41356 34524 41412
rect 34580 41356 35644 41412
rect 35700 41356 37100 41412
rect 37156 41356 37166 41412
rect 49970 41356 49980 41412
rect 50036 41356 56588 41412
rect 56644 41356 57372 41412
rect 57428 41356 57932 41412
rect 57988 41356 57998 41412
rect 25004 41300 25060 41356
rect 28252 41300 28308 41356
rect 23202 41244 23212 41300
rect 23268 41244 25004 41300
rect 25060 41244 25070 41300
rect 25218 41244 25228 41300
rect 25284 41244 28308 41300
rect 28802 41244 28812 41300
rect 28868 41244 30156 41300
rect 30212 41244 30222 41300
rect 35756 41244 36428 41300
rect 36484 41244 36494 41300
rect 43810 41244 43820 41300
rect 43876 41244 46956 41300
rect 47012 41244 49084 41300
rect 49140 41244 49150 41300
rect 52994 41244 53004 41300
rect 53060 41244 53676 41300
rect 53732 41244 54460 41300
rect 54516 41244 54526 41300
rect 35756 41076 35812 41244
rect 35970 41132 35980 41188
rect 36036 41132 37772 41188
rect 37828 41132 37838 41188
rect 38882 41132 38892 41188
rect 38948 41132 39452 41188
rect 39508 41132 39518 41188
rect 49410 41132 49420 41188
rect 49476 41132 51212 41188
rect 51268 41132 52108 41188
rect 52164 41132 52174 41188
rect 53330 41132 53340 41188
rect 53396 41132 53564 41188
rect 53620 41132 53630 41188
rect 57138 41132 57148 41188
rect 57204 41132 57596 41188
rect 57652 41132 57662 41188
rect 2594 41020 2604 41076
rect 2660 41020 5684 41076
rect 6038 41020 6076 41076
rect 6132 41020 6142 41076
rect 7410 41020 7420 41076
rect 7476 41020 8652 41076
rect 8708 41020 9212 41076
rect 9268 41020 9278 41076
rect 9426 41020 9436 41076
rect 9492 41020 12460 41076
rect 12516 41020 12526 41076
rect 12908 41020 13692 41076
rect 13748 41020 13758 41076
rect 14242 41020 14252 41076
rect 14308 41020 15036 41076
rect 15092 41020 15102 41076
rect 15250 41020 15260 41076
rect 15316 41020 15372 41076
rect 15428 41020 15438 41076
rect 16930 41020 16940 41076
rect 16996 41020 17612 41076
rect 17668 41020 17678 41076
rect 18722 41020 18732 41076
rect 18788 41020 20412 41076
rect 20468 41020 21420 41076
rect 21476 41020 21486 41076
rect 22866 41020 22876 41076
rect 22932 41020 22942 41076
rect 25218 41020 25228 41076
rect 25284 41020 26460 41076
rect 26516 41020 26526 41076
rect 28130 41020 28140 41076
rect 28196 41020 35812 41076
rect 38546 41020 38556 41076
rect 38612 41020 43596 41076
rect 43652 41020 44604 41076
rect 44660 41020 44670 41076
rect 46834 41020 46844 41076
rect 46900 41020 47404 41076
rect 47460 41020 47470 41076
rect 12908 40964 12964 41020
rect 4162 40908 4172 40964
rect 4228 40908 5068 40964
rect 5124 40908 5134 40964
rect 7522 40908 7532 40964
rect 7588 40908 8092 40964
rect 8148 40908 9772 40964
rect 9828 40908 12964 40964
rect 13020 40908 16380 40964
rect 16436 40908 16716 40964
rect 16772 40908 17668 40964
rect 17826 40908 17836 40964
rect 17892 40908 20636 40964
rect 20692 40908 20702 40964
rect 27122 40908 27132 40964
rect 27188 40908 33628 40964
rect 33684 40908 35196 40964
rect 35252 40908 36988 40964
rect 37044 40908 37054 40964
rect 39890 40908 39900 40964
rect 39956 40908 41244 40964
rect 41300 40908 41310 40964
rect 41794 40908 41804 40964
rect 41860 40908 43036 40964
rect 43092 40908 43102 40964
rect 49186 40908 49196 40964
rect 49252 40908 50204 40964
rect 50260 40908 50764 40964
rect 50820 40908 50830 40964
rect 51650 40908 51660 40964
rect 51716 40908 51884 40964
rect 51940 40908 52444 40964
rect 52500 40908 52668 40964
rect 52724 40908 52734 40964
rect 53554 40908 53564 40964
rect 53620 40908 54460 40964
rect 54516 40908 55020 40964
rect 55076 40908 55804 40964
rect 55860 40908 57036 40964
rect 57092 40908 57102 40964
rect 13020 40852 13076 40908
rect 17612 40852 17668 40908
rect 6738 40796 6748 40852
rect 6804 40796 7756 40852
rect 7812 40796 11564 40852
rect 11620 40796 11630 40852
rect 13010 40796 13020 40852
rect 13076 40796 13086 40852
rect 13244 40796 16604 40852
rect 16660 40796 16670 40852
rect 17612 40796 18732 40852
rect 18788 40796 18798 40852
rect 19506 40796 19516 40852
rect 19572 40796 19628 40852
rect 19684 40796 19694 40852
rect 22306 40796 22316 40852
rect 22372 40796 24332 40852
rect 24388 40796 25900 40852
rect 25956 40796 25966 40852
rect 29362 40796 29372 40852
rect 29428 40796 29820 40852
rect 29876 40796 29886 40852
rect 32274 40796 32284 40852
rect 32340 40796 33404 40852
rect 33460 40796 33470 40852
rect 39218 40796 39228 40852
rect 39284 40796 42140 40852
rect 42196 40796 42206 40852
rect 13244 40740 13300 40796
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 25900 40740 25956 40796
rect 43652 40740 43708 40852
rect 43764 40796 43774 40852
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 4722 40684 4732 40740
rect 4788 40684 9100 40740
rect 9156 40684 9166 40740
rect 12674 40684 12684 40740
rect 12740 40684 13300 40740
rect 14466 40684 14476 40740
rect 14532 40684 15596 40740
rect 15652 40684 15662 40740
rect 16370 40684 16380 40740
rect 16436 40684 16604 40740
rect 16660 40684 16670 40740
rect 16864 40684 16940 40740
rect 16996 40684 17388 40740
rect 17444 40684 17454 40740
rect 20738 40684 20748 40740
rect 20804 40684 21756 40740
rect 21812 40684 21822 40740
rect 25900 40684 27580 40740
rect 27636 40684 27804 40740
rect 27860 40684 27870 40740
rect 36306 40684 36316 40740
rect 36372 40684 42700 40740
rect 42756 40684 43148 40740
rect 43204 40684 43708 40740
rect 4274 40572 4284 40628
rect 4340 40572 4844 40628
rect 4900 40572 4910 40628
rect 6374 40572 6412 40628
rect 6468 40572 6478 40628
rect 6962 40572 6972 40628
rect 7028 40572 7196 40628
rect 7252 40572 7262 40628
rect 7970 40572 7980 40628
rect 8036 40572 8316 40628
rect 8372 40572 8382 40628
rect 11638 40572 11676 40628
rect 11732 40572 11742 40628
rect 13906 40572 13916 40628
rect 13972 40572 14364 40628
rect 14420 40572 14430 40628
rect 14662 40572 14700 40628
rect 14756 40572 14766 40628
rect 18162 40572 18172 40628
rect 18228 40572 19180 40628
rect 19236 40572 19628 40628
rect 19684 40572 19694 40628
rect 21298 40572 21308 40628
rect 21364 40572 21980 40628
rect 22036 40572 22046 40628
rect 22194 40572 22204 40628
rect 22260 40572 23996 40628
rect 24052 40572 24444 40628
rect 24500 40572 24510 40628
rect 26562 40572 26572 40628
rect 26628 40572 26796 40628
rect 26852 40572 26862 40628
rect 28018 40572 28028 40628
rect 28084 40572 28588 40628
rect 28644 40572 28654 40628
rect 30818 40572 30828 40628
rect 30884 40572 32284 40628
rect 32340 40572 32350 40628
rect 33506 40572 33516 40628
rect 33572 40572 35980 40628
rect 36036 40572 36046 40628
rect 40674 40572 40684 40628
rect 40740 40572 41468 40628
rect 41524 40572 42476 40628
rect 42532 40572 42542 40628
rect 2818 40460 2828 40516
rect 2884 40460 3500 40516
rect 3556 40460 3566 40516
rect 4946 40460 4956 40516
rect 5012 40460 5964 40516
rect 6020 40460 6636 40516
rect 6692 40460 6702 40516
rect 7858 40460 7868 40516
rect 7924 40460 7980 40516
rect 8036 40460 8046 40516
rect 11190 40460 11228 40516
rect 11284 40460 11294 40516
rect 11974 40460 12012 40516
rect 12068 40460 13020 40516
rect 13076 40460 13086 40516
rect 13468 40460 15036 40516
rect 15092 40460 15102 40516
rect 15222 40460 15260 40516
rect 15316 40460 16268 40516
rect 16324 40460 16334 40516
rect 16482 40460 16492 40516
rect 16548 40460 20524 40516
rect 20580 40460 20590 40516
rect 20962 40460 20972 40516
rect 21028 40460 22316 40516
rect 22372 40460 22382 40516
rect 22642 40460 22652 40516
rect 22708 40460 26908 40516
rect 26964 40460 27244 40516
rect 27300 40460 27692 40516
rect 27748 40460 27758 40516
rect 28028 40460 35532 40516
rect 35588 40460 35598 40516
rect 38434 40460 38444 40516
rect 38500 40460 40012 40516
rect 40068 40460 40078 40516
rect 46162 40460 46172 40516
rect 46228 40460 46844 40516
rect 46900 40460 47180 40516
rect 47236 40460 47246 40516
rect 48514 40460 48524 40516
rect 48580 40460 50764 40516
rect 50820 40460 50830 40516
rect 57698 40460 57708 40516
rect 57764 40460 57774 40516
rect 13468 40404 13524 40460
rect 28028 40404 28084 40460
rect 2706 40348 2716 40404
rect 2772 40348 3388 40404
rect 3444 40348 3454 40404
rect 5058 40348 5068 40404
rect 5124 40348 5134 40404
rect 6738 40348 6748 40404
rect 6804 40348 8652 40404
rect 8708 40348 8718 40404
rect 10546 40348 10556 40404
rect 10612 40348 11564 40404
rect 11620 40348 11630 40404
rect 12114 40348 12124 40404
rect 12180 40348 13524 40404
rect 13682 40348 13692 40404
rect 13748 40348 16044 40404
rect 16100 40348 18284 40404
rect 18340 40348 18350 40404
rect 18470 40348 18508 40404
rect 18564 40348 18574 40404
rect 18834 40348 18844 40404
rect 18900 40348 21196 40404
rect 21252 40348 21262 40404
rect 21522 40348 21532 40404
rect 21588 40348 21868 40404
rect 21924 40348 21934 40404
rect 22866 40348 22876 40404
rect 22932 40348 23660 40404
rect 23716 40348 23726 40404
rect 25330 40348 25340 40404
rect 25396 40348 26236 40404
rect 26292 40348 26302 40404
rect 27122 40348 27132 40404
rect 27188 40348 28028 40404
rect 28084 40348 28094 40404
rect 32386 40348 32396 40404
rect 32452 40348 33068 40404
rect 33124 40348 33134 40404
rect 34738 40348 34748 40404
rect 34804 40348 37660 40404
rect 37716 40348 37726 40404
rect 37986 40348 37996 40404
rect 38052 40348 38556 40404
rect 38612 40348 38892 40404
rect 38948 40348 38958 40404
rect 43698 40348 43708 40404
rect 43764 40348 44268 40404
rect 44324 40348 44334 40404
rect 45042 40348 45052 40404
rect 45108 40348 46060 40404
rect 46116 40348 46956 40404
rect 47012 40348 47022 40404
rect 47842 40348 47852 40404
rect 47908 40348 53228 40404
rect 53284 40348 53294 40404
rect 5068 40292 5124 40348
rect 57708 40292 57764 40460
rect 1586 40236 1596 40292
rect 1652 40236 5124 40292
rect 5842 40236 5852 40292
rect 5908 40236 11116 40292
rect 11172 40236 11182 40292
rect 11330 40236 11340 40292
rect 11396 40236 15372 40292
rect 15428 40236 15438 40292
rect 18610 40236 18620 40292
rect 18676 40236 18844 40292
rect 18900 40236 18910 40292
rect 19282 40236 19292 40292
rect 19348 40236 20188 40292
rect 20244 40236 20254 40292
rect 24770 40236 24780 40292
rect 24836 40236 25564 40292
rect 25620 40236 25630 40292
rect 31714 40236 31724 40292
rect 31780 40236 32844 40292
rect 32900 40236 33516 40292
rect 33572 40236 33582 40292
rect 34178 40236 34188 40292
rect 34244 40236 36092 40292
rect 36148 40236 36428 40292
rect 36484 40236 36494 40292
rect 36642 40236 36652 40292
rect 36708 40236 37324 40292
rect 37380 40236 37390 40292
rect 38994 40236 39004 40292
rect 39060 40236 46732 40292
rect 46788 40236 46798 40292
rect 57708 40236 58268 40292
rect 58324 40236 58334 40292
rect 5068 40180 5124 40236
rect 2034 40124 2044 40180
rect 2100 40124 2380 40180
rect 2436 40124 2604 40180
rect 2660 40124 2670 40180
rect 5068 40124 7308 40180
rect 7364 40124 7374 40180
rect 9426 40124 9436 40180
rect 9492 40124 9772 40180
rect 9828 40124 9838 40180
rect 10546 40124 10556 40180
rect 10612 40124 15372 40180
rect 15428 40124 15438 40180
rect 17938 40124 17948 40180
rect 18004 40124 20188 40180
rect 20244 40124 20254 40180
rect 26114 40124 26124 40180
rect 26180 40124 27692 40180
rect 27748 40124 27758 40180
rect 34290 40124 34300 40180
rect 34356 40124 36484 40180
rect 40226 40124 40236 40180
rect 40292 40124 40796 40180
rect 40852 40124 41132 40180
rect 41188 40124 41198 40180
rect 45490 40124 45500 40180
rect 45556 40124 45724 40180
rect 45780 40124 45790 40180
rect 36428 40068 36484 40124
rect 914 40012 924 40068
rect 980 40012 1596 40068
rect 1652 40012 1662 40068
rect 3378 40012 3388 40068
rect 3444 40012 3948 40068
rect 4004 40012 4014 40068
rect 5058 40012 5068 40068
rect 5124 40012 7308 40068
rect 7364 40012 7374 40068
rect 8530 40012 8540 40068
rect 8596 40012 9996 40068
rect 10052 40012 10444 40068
rect 10500 40012 10948 40068
rect 11666 40012 11676 40068
rect 11732 40012 18844 40068
rect 18900 40012 18910 40068
rect 22978 40012 22988 40068
rect 23044 40012 27244 40068
rect 27300 40012 27310 40068
rect 36418 40012 36428 40068
rect 36484 40012 36494 40068
rect 2370 39900 2380 39956
rect 2436 39900 3388 39956
rect 3444 39900 3454 39956
rect 3948 39844 4004 40012
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 10892 39956 10948 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 5618 39900 5628 39956
rect 5684 39900 5740 39956
rect 5796 39900 5806 39956
rect 7634 39900 7644 39956
rect 7700 39900 7980 39956
rect 8036 39900 8046 39956
rect 10892 39900 12012 39956
rect 12068 39900 12078 39956
rect 12674 39900 12684 39956
rect 12740 39900 14812 39956
rect 14868 39900 14878 39956
rect 27346 39900 27356 39956
rect 27412 39900 29820 39956
rect 29876 39900 31836 39956
rect 31892 39900 31902 39956
rect 3042 39788 3052 39844
rect 3108 39788 3500 39844
rect 3556 39788 3612 39844
rect 3668 39788 3678 39844
rect 3948 39788 7084 39844
rect 7140 39788 7150 39844
rect 7746 39788 7756 39844
rect 7812 39788 14364 39844
rect 14420 39788 14430 39844
rect 15362 39788 15372 39844
rect 15428 39788 16828 39844
rect 16884 39788 16894 39844
rect 17602 39788 17612 39844
rect 17668 39788 18060 39844
rect 18116 39788 18126 39844
rect 23538 39788 23548 39844
rect 23604 39788 23614 39844
rect 26338 39788 26348 39844
rect 26404 39788 27132 39844
rect 27188 39788 27198 39844
rect 23548 39732 23604 39788
rect 3378 39676 3388 39732
rect 3444 39676 4060 39732
rect 4116 39676 5180 39732
rect 5236 39676 5246 39732
rect 6290 39676 6300 39732
rect 6356 39676 10108 39732
rect 10164 39676 10174 39732
rect 12898 39676 12908 39732
rect 12964 39676 15036 39732
rect 15092 39676 15102 39732
rect 16258 39676 16268 39732
rect 16324 39676 17164 39732
rect 17220 39676 17724 39732
rect 17780 39676 17790 39732
rect 18610 39676 18620 39732
rect 18676 39676 19404 39732
rect 19460 39676 19470 39732
rect 19954 39676 19964 39732
rect 20020 39676 23324 39732
rect 23380 39676 23390 39732
rect 23548 39676 25116 39732
rect 25172 39676 40460 39732
rect 40516 39676 42140 39732
rect 42196 39676 42588 39732
rect 42644 39676 42654 39732
rect 3332 39564 4956 39620
rect 5012 39564 5022 39620
rect 6290 39564 6300 39620
rect 6356 39564 6636 39620
rect 6692 39564 6702 39620
rect 7830 39564 7868 39620
rect 7924 39564 7934 39620
rect 8082 39564 8092 39620
rect 8148 39564 9884 39620
rect 9940 39564 9950 39620
rect 10210 39564 10220 39620
rect 10276 39564 11564 39620
rect 11620 39564 13692 39620
rect 13748 39564 13758 39620
rect 16678 39564 16716 39620
rect 16772 39564 16782 39620
rect 16940 39564 18284 39620
rect 18340 39564 18350 39620
rect 18694 39564 18732 39620
rect 18788 39564 18798 39620
rect 20962 39564 20972 39620
rect 21028 39564 23884 39620
rect 23940 39564 23950 39620
rect 27122 39564 27132 39620
rect 27188 39564 27692 39620
rect 27748 39564 32172 39620
rect 32228 39564 32238 39620
rect 34514 39564 34524 39620
rect 34580 39564 34972 39620
rect 35028 39564 36092 39620
rect 36148 39564 36158 39620
rect 41570 39564 41580 39620
rect 41636 39564 42924 39620
rect 42980 39564 43148 39620
rect 43204 39564 43214 39620
rect 46722 39564 46732 39620
rect 46788 39564 47292 39620
rect 47348 39564 47358 39620
rect 56802 39564 56812 39620
rect 56868 39564 57820 39620
rect 57876 39564 58268 39620
rect 58324 39564 58334 39620
rect 3332 39508 3388 39564
rect 16940 39508 16996 39564
rect 2146 39452 2156 39508
rect 2212 39452 3388 39508
rect 3500 39452 4452 39508
rect 4610 39452 4620 39508
rect 4676 39452 11452 39508
rect 11508 39452 11676 39508
rect 11732 39452 11742 39508
rect 11890 39452 11900 39508
rect 11956 39452 11994 39508
rect 12450 39452 12460 39508
rect 12516 39452 14140 39508
rect 14196 39452 16996 39508
rect 17154 39452 17164 39508
rect 17220 39452 17948 39508
rect 18004 39452 18014 39508
rect 18610 39452 18620 39508
rect 18676 39452 19628 39508
rect 19684 39452 19852 39508
rect 19908 39452 19918 39508
rect 26114 39452 26124 39508
rect 26180 39452 28476 39508
rect 28532 39452 28542 39508
rect 34626 39452 34636 39508
rect 34692 39452 35868 39508
rect 35924 39452 35934 39508
rect 44706 39452 44716 39508
rect 44772 39452 47964 39508
rect 48020 39452 48030 39508
rect 53554 39452 53564 39508
rect 53620 39452 54684 39508
rect 54740 39452 54750 39508
rect 3500 39396 3556 39452
rect 2034 39340 2044 39396
rect 2100 39340 3276 39396
rect 3332 39340 3556 39396
rect 2594 39228 2604 39284
rect 2660 39228 3612 39284
rect 3668 39228 3678 39284
rect 3826 39228 3836 39284
rect 3892 39228 4116 39284
rect 4060 39172 4116 39228
rect 3612 39116 3724 39172
rect 3780 39116 3790 39172
rect 4050 39116 4060 39172
rect 4116 39116 4126 39172
rect 1810 38892 1820 38948
rect 1876 38892 3388 38948
rect 3444 38892 3454 38948
rect 3612 38836 3668 39116
rect 4396 39060 4452 39452
rect 5142 39340 5180 39396
rect 5236 39340 5246 39396
rect 6178 39340 6188 39396
rect 6244 39340 7644 39396
rect 7700 39340 11564 39396
rect 11620 39340 12236 39396
rect 12292 39340 12302 39396
rect 13542 39340 13580 39396
rect 13636 39340 14700 39396
rect 14756 39340 14766 39396
rect 15138 39340 15148 39396
rect 15204 39340 15372 39396
rect 15428 39340 15438 39396
rect 15698 39340 15708 39396
rect 15764 39340 16156 39396
rect 16212 39340 18396 39396
rect 18452 39340 18462 39396
rect 18806 39340 18844 39396
rect 18900 39340 18910 39396
rect 19058 39340 19068 39396
rect 19124 39340 20076 39396
rect 20132 39340 20142 39396
rect 25442 39340 25452 39396
rect 25508 39340 31724 39396
rect 31780 39340 33292 39396
rect 33348 39340 33358 39396
rect 46498 39340 46508 39396
rect 46564 39340 47068 39396
rect 47124 39340 47134 39396
rect 48626 39340 48636 39396
rect 48692 39340 49308 39396
rect 49364 39340 49868 39396
rect 49924 39340 49934 39396
rect 6178 39228 6188 39284
rect 6244 39228 10220 39284
rect 10276 39228 10286 39284
rect 11936 39228 12012 39284
rect 12068 39228 12572 39284
rect 12628 39228 12638 39284
rect 13234 39228 13244 39284
rect 13300 39228 16380 39284
rect 16436 39228 16446 39284
rect 16902 39228 16940 39284
rect 16996 39228 17006 39284
rect 17238 39228 17276 39284
rect 17332 39228 17342 39284
rect 17686 39228 17724 39284
rect 17780 39228 17790 39284
rect 18274 39228 18284 39284
rect 18340 39228 19292 39284
rect 19348 39228 19358 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 5506 39116 5516 39172
rect 5572 39116 6860 39172
rect 6916 39116 6926 39172
rect 8306 39116 8316 39172
rect 8372 39116 12180 39172
rect 13794 39116 13804 39172
rect 13860 39116 14028 39172
rect 14084 39116 14476 39172
rect 14532 39116 14542 39172
rect 15026 39116 15036 39172
rect 15092 39116 19348 39172
rect 23062 39116 23100 39172
rect 23156 39116 23166 39172
rect 27794 39116 27804 39172
rect 27860 39116 33852 39172
rect 33908 39116 34524 39172
rect 34580 39116 37548 39172
rect 37604 39116 37614 39172
rect 12124 39060 12180 39116
rect 19292 39060 19348 39116
rect 3798 39004 3836 39060
rect 3892 39004 3902 39060
rect 4396 39004 7756 39060
rect 7812 39004 7980 39060
rect 8036 39004 8372 39060
rect 8978 39004 8988 39060
rect 9044 39004 9772 39060
rect 9828 39004 10444 39060
rect 10500 39004 10510 39060
rect 12114 39004 12124 39060
rect 12180 39004 12460 39060
rect 12516 39004 13916 39060
rect 13972 39004 13982 39060
rect 14130 39004 14140 39060
rect 14196 39004 14924 39060
rect 14980 39004 14990 39060
rect 15082 39004 15092 39060
rect 15148 39004 15484 39060
rect 15540 39004 16268 39060
rect 16324 39004 16334 39060
rect 16706 39004 16716 39060
rect 16772 39004 18508 39060
rect 18564 39004 18574 39060
rect 18918 39004 18956 39060
rect 19012 39004 19022 39060
rect 19292 39004 23548 39060
rect 23604 39004 23614 39060
rect 34066 39004 34076 39060
rect 34132 39004 34636 39060
rect 34692 39004 34702 39060
rect 36530 39004 36540 39060
rect 36596 39004 37100 39060
rect 37156 39004 37166 39060
rect 42018 39004 42028 39060
rect 42084 39004 42812 39060
rect 42868 39004 44996 39060
rect 8316 38948 8372 39004
rect 4208 38892 4284 38948
rect 4340 38892 4620 38948
rect 4676 38892 4686 38948
rect 4834 38892 4844 38948
rect 4900 38892 6300 38948
rect 6356 38892 6366 38948
rect 7298 38892 7308 38948
rect 7364 38892 8092 38948
rect 8148 38892 8158 38948
rect 8306 38892 8316 38948
rect 8372 38892 8382 38948
rect 9986 38892 9996 38948
rect 10052 38892 10668 38948
rect 10724 38892 10734 38948
rect 14018 38892 14028 38948
rect 14084 38892 14476 38948
rect 14532 38892 14542 38948
rect 14802 38892 14812 38948
rect 14868 38892 15372 38948
rect 15428 38892 15438 38948
rect 15586 38892 15596 38948
rect 15652 38892 18284 38948
rect 18340 38892 18350 38948
rect 19170 38892 19180 38948
rect 19236 38892 20188 38948
rect 20244 38892 20636 38948
rect 20692 38892 20702 38948
rect 23090 38892 23100 38948
rect 23156 38892 23996 38948
rect 24052 38892 25788 38948
rect 25844 38892 26348 38948
rect 26404 38892 26414 38948
rect 30716 38892 31500 38948
rect 31556 38892 31566 38948
rect 33618 38892 33628 38948
rect 33684 38892 37324 38948
rect 37380 38892 37390 38948
rect 40786 38892 40796 38948
rect 40852 38892 44268 38948
rect 44324 38892 44334 38948
rect 30716 38836 30772 38892
rect 44940 38836 44996 39004
rect 49858 38892 49868 38948
rect 49924 38892 50876 38948
rect 50932 38892 50942 38948
rect 52210 38892 52220 38948
rect 52276 38892 53564 38948
rect 53620 38892 53630 38948
rect 1362 38780 1372 38836
rect 1428 38780 2044 38836
rect 2100 38780 2492 38836
rect 2548 38780 2558 38836
rect 3612 38780 6076 38836
rect 6132 38780 6142 38836
rect 7606 38780 7644 38836
rect 7700 38780 7710 38836
rect 7970 38780 7980 38836
rect 8036 38780 8428 38836
rect 8484 38780 11788 38836
rect 11844 38780 12348 38836
rect 12404 38780 13356 38836
rect 13412 38780 13422 38836
rect 14802 38780 14812 38836
rect 14868 38780 16156 38836
rect 16212 38780 16222 38836
rect 17350 38780 17388 38836
rect 17444 38780 17454 38836
rect 17826 38780 17836 38836
rect 17892 38780 19404 38836
rect 19460 38780 19470 38836
rect 21494 38780 21532 38836
rect 21588 38780 21598 38836
rect 29036 38780 30044 38836
rect 30100 38780 30716 38836
rect 30772 38780 30782 38836
rect 31266 38780 31276 38836
rect 31332 38780 44492 38836
rect 44548 38780 44558 38836
rect 44930 38780 44940 38836
rect 44996 38780 45780 38836
rect 46722 38780 46732 38836
rect 46788 38780 48076 38836
rect 48132 38780 48142 38836
rect 50082 38780 50092 38836
rect 50148 38780 50540 38836
rect 50596 38780 51324 38836
rect 51380 38780 51390 38836
rect 56690 38780 56700 38836
rect 56756 38780 57932 38836
rect 57988 38780 57998 38836
rect 29036 38724 29092 38780
rect 45724 38724 45780 38780
rect 1922 38668 1932 38724
rect 1988 38668 2324 38724
rect 2482 38668 2492 38724
rect 2548 38668 2940 38724
rect 2996 38668 3388 38724
rect 3444 38668 3454 38724
rect 5590 38668 5628 38724
rect 5684 38668 5694 38724
rect 6262 38668 6300 38724
rect 6356 38668 6366 38724
rect 7074 38668 7084 38724
rect 7140 38668 7980 38724
rect 8036 38668 9212 38724
rect 9268 38668 10108 38724
rect 10164 38668 10174 38724
rect 11788 38668 12684 38724
rect 12740 38668 12750 38724
rect 15138 38668 15148 38724
rect 15204 38668 15372 38724
rect 15428 38668 16604 38724
rect 16660 38668 16670 38724
rect 18162 38668 18172 38724
rect 18228 38668 20748 38724
rect 20804 38668 20814 38724
rect 22978 38668 22988 38724
rect 23044 38668 25900 38724
rect 25956 38668 25966 38724
rect 29026 38668 29036 38724
rect 29092 38668 29102 38724
rect 29810 38668 29820 38724
rect 29876 38668 30604 38724
rect 30660 38668 31500 38724
rect 31556 38668 31566 38724
rect 31826 38668 31836 38724
rect 31892 38668 34188 38724
rect 34244 38668 34254 38724
rect 37090 38668 37100 38724
rect 37156 38668 38668 38724
rect 38724 38668 38780 38724
rect 38836 38668 38846 38724
rect 42914 38668 42924 38724
rect 42980 38668 43708 38724
rect 43764 38668 43774 38724
rect 45714 38668 45724 38724
rect 45780 38668 46060 38724
rect 46116 38668 46284 38724
rect 46340 38668 46350 38724
rect 48738 38668 48748 38724
rect 48804 38668 49980 38724
rect 50036 38668 51436 38724
rect 51492 38668 51502 38724
rect 53890 38668 53900 38724
rect 53956 38668 54572 38724
rect 54628 38668 54638 38724
rect 55570 38668 55580 38724
rect 55636 38668 56364 38724
rect 56420 38668 57596 38724
rect 57652 38668 57662 38724
rect 2258 38612 2268 38668
rect 2324 38612 2334 38668
rect 11788 38612 11844 38668
rect 7084 38556 7756 38612
rect 7812 38556 9324 38612
rect 9380 38556 11844 38612
rect 13244 38556 16940 38612
rect 16996 38556 17006 38612
rect 17602 38556 17612 38612
rect 17668 38556 19292 38612
rect 19348 38556 19628 38612
rect 19684 38556 19694 38612
rect 36866 38556 36876 38612
rect 36932 38556 37772 38612
rect 37828 38556 46172 38612
rect 46228 38556 46238 38612
rect 7084 38500 7140 38556
rect 13244 38500 13300 38556
rect 14812 38500 14868 38556
rect 3826 38444 3836 38500
rect 3892 38444 4172 38500
rect 4228 38444 4238 38500
rect 6626 38444 6636 38500
rect 6692 38444 7140 38500
rect 7410 38444 7420 38500
rect 7476 38444 8204 38500
rect 8260 38444 8270 38500
rect 11218 38444 11228 38500
rect 11284 38444 13300 38500
rect 14802 38444 14812 38500
rect 14868 38444 14878 38500
rect 16034 38444 16044 38500
rect 16100 38444 19404 38500
rect 19460 38444 19470 38500
rect 22866 38444 22876 38500
rect 22932 38444 23548 38500
rect 23604 38444 23772 38500
rect 23828 38444 26572 38500
rect 26628 38444 26638 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 5058 38332 5068 38388
rect 5124 38332 5740 38388
rect 5796 38332 5806 38388
rect 6738 38332 6748 38388
rect 6804 38332 8652 38388
rect 8708 38332 8718 38388
rect 14914 38332 14924 38388
rect 14980 38332 24332 38388
rect 24388 38332 25004 38388
rect 25060 38332 25070 38388
rect 4050 38220 4060 38276
rect 4116 38220 4620 38276
rect 4676 38220 4686 38276
rect 8082 38220 8092 38276
rect 8148 38220 8988 38276
rect 9044 38220 9054 38276
rect 10322 38220 10332 38276
rect 10388 38220 12908 38276
rect 12964 38220 12974 38276
rect 14214 38220 14252 38276
rect 14308 38220 14318 38276
rect 15138 38220 15148 38276
rect 15204 38220 15932 38276
rect 15988 38220 15998 38276
rect 27234 38220 27244 38276
rect 27300 38220 33404 38276
rect 33460 38220 33852 38276
rect 33908 38220 34412 38276
rect 34468 38220 34478 38276
rect 1474 38108 1484 38164
rect 1540 38108 2380 38164
rect 2436 38108 2446 38164
rect 2594 38108 2604 38164
rect 2660 38108 3388 38164
rect 5058 38108 5068 38164
rect 5124 38108 7420 38164
rect 7476 38108 7486 38164
rect 8754 38108 8764 38164
rect 8820 38108 11676 38164
rect 11732 38108 11742 38164
rect 12562 38108 12572 38164
rect 12628 38108 15036 38164
rect 15092 38108 15102 38164
rect 17042 38108 17052 38164
rect 17108 38108 18172 38164
rect 18228 38108 22652 38164
rect 22708 38108 22718 38164
rect 25666 38108 25676 38164
rect 25732 38108 29260 38164
rect 29316 38108 29708 38164
rect 29764 38108 29774 38164
rect 33292 38108 36316 38164
rect 36372 38108 36382 38164
rect 40114 38108 40124 38164
rect 40180 38108 40908 38164
rect 40964 38108 40974 38164
rect 50754 38108 50764 38164
rect 50820 38108 51884 38164
rect 51940 38108 51950 38164
rect 3332 38052 3388 38108
rect 3332 37996 4060 38052
rect 4116 37996 4126 38052
rect 4274 37996 4284 38052
rect 4340 37996 6524 38052
rect 6580 37996 6748 38052
rect 6804 37996 6814 38052
rect 7074 37996 7084 38052
rect 7140 37996 9100 38052
rect 9156 37996 10220 38052
rect 10276 37996 10286 38052
rect 10434 37996 10444 38052
rect 10500 37996 10892 38052
rect 10948 37996 10958 38052
rect 12114 37996 12124 38052
rect 12180 37996 18284 38052
rect 18340 37996 18350 38052
rect 19954 37996 19964 38052
rect 20020 37996 21868 38052
rect 21924 37996 21934 38052
rect 33292 37940 33348 38108
rect 34178 37996 34188 38052
rect 34244 37996 38332 38052
rect 38388 37996 38398 38052
rect 38994 37996 39004 38052
rect 39060 37996 40236 38052
rect 40292 37996 40302 38052
rect 44146 37996 44156 38052
rect 44212 37996 50428 38052
rect 50484 37996 51772 38052
rect 51828 37996 51838 38052
rect 4274 37884 4284 37940
rect 4340 37884 5068 37940
rect 5124 37884 6188 37940
rect 6244 37884 6254 37940
rect 6626 37884 6636 37940
rect 6692 37884 7532 37940
rect 7588 37884 7598 37940
rect 9202 37884 9212 37940
rect 9268 37884 9772 37940
rect 9828 37884 14588 37940
rect 14644 37884 14654 37940
rect 15026 37884 15036 37940
rect 15092 37884 23548 37940
rect 23604 37884 23996 37940
rect 24052 37884 24556 37940
rect 24612 37884 26124 37940
rect 26180 37884 26190 37940
rect 27570 37884 27580 37940
rect 27636 37884 27804 37940
rect 27860 37884 27870 37940
rect 32050 37884 32060 37940
rect 32116 37884 33068 37940
rect 33124 37884 33292 37940
rect 33348 37884 33358 37940
rect 33618 37884 33628 37940
rect 33684 37884 34524 37940
rect 34580 37884 34972 37940
rect 35028 37884 35196 37940
rect 35252 37884 35262 37940
rect 53330 37884 53340 37940
rect 53396 37884 54908 37940
rect 54964 37884 54974 37940
rect 3266 37772 3276 37828
rect 3332 37772 4172 37828
rect 4228 37772 4238 37828
rect 6402 37772 6412 37828
rect 6468 37772 10668 37828
rect 10724 37772 11116 37828
rect 11172 37772 11900 37828
rect 11956 37772 11966 37828
rect 18610 37772 18620 37828
rect 18676 37772 19068 37828
rect 19124 37772 24108 37828
rect 24164 37772 24174 37828
rect 31602 37772 31612 37828
rect 31668 37772 32620 37828
rect 32676 37772 32686 37828
rect 34290 37772 34300 37828
rect 34356 37772 36204 37828
rect 36260 37772 36540 37828
rect 36596 37772 36606 37828
rect 38098 37772 38108 37828
rect 38164 37772 45724 37828
rect 45780 37772 46284 37828
rect 46340 37772 46350 37828
rect 3602 37660 3612 37716
rect 3668 37660 4060 37716
rect 4116 37660 4126 37716
rect 4498 37660 4508 37716
rect 4564 37660 4956 37716
rect 5012 37660 9212 37716
rect 9268 37660 9278 37716
rect 12562 37660 12572 37716
rect 12628 37660 15148 37716
rect 17602 37660 17612 37716
rect 17668 37660 17836 37716
rect 17892 37660 17902 37716
rect 39666 37660 39676 37716
rect 39732 37660 40236 37716
rect 40292 37660 40302 37716
rect 15092 37604 15148 37660
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 3490 37548 3500 37604
rect 3556 37548 10780 37604
rect 10836 37548 11116 37604
rect 11172 37548 11182 37604
rect 11442 37548 11452 37604
rect 11508 37548 12124 37604
rect 12180 37548 12190 37604
rect 12786 37548 12796 37604
rect 12852 37548 13580 37604
rect 13636 37548 13646 37604
rect 13794 37548 13804 37604
rect 13860 37548 13898 37604
rect 14242 37548 14252 37604
rect 14308 37548 14364 37604
rect 14420 37548 14430 37604
rect 15092 37548 15372 37604
rect 15428 37548 18172 37604
rect 18228 37548 18238 37604
rect 27346 37548 27356 37604
rect 27412 37548 27916 37604
rect 27972 37548 27982 37604
rect 31378 37548 31388 37604
rect 31444 37548 34188 37604
rect 34244 37548 35308 37604
rect 35364 37548 35374 37604
rect 38434 37548 38444 37604
rect 38500 37548 38668 37604
rect 38724 37548 38734 37604
rect 38994 37548 39004 37604
rect 39060 37548 39564 37604
rect 39620 37548 39630 37604
rect 1586 37436 1596 37492
rect 1652 37436 5628 37492
rect 5684 37436 5694 37492
rect 6738 37436 6748 37492
rect 6804 37436 10388 37492
rect 10546 37436 10556 37492
rect 10612 37436 19964 37492
rect 20020 37436 21868 37492
rect 21924 37436 21934 37492
rect 22082 37436 22092 37492
rect 22148 37436 22764 37492
rect 22820 37436 22830 37492
rect 22978 37436 22988 37492
rect 23044 37436 28700 37492
rect 28756 37436 28766 37492
rect 29698 37436 29708 37492
rect 29764 37436 30716 37492
rect 30772 37436 31724 37492
rect 31780 37436 31790 37492
rect 32386 37436 32396 37492
rect 32452 37436 33292 37492
rect 33348 37436 33358 37492
rect 38322 37436 38332 37492
rect 38388 37436 38780 37492
rect 38836 37436 38846 37492
rect 39330 37436 39340 37492
rect 39396 37436 39900 37492
rect 39956 37436 41468 37492
rect 41524 37436 41534 37492
rect 53218 37436 53228 37492
rect 53284 37436 54348 37492
rect 54404 37436 55244 37492
rect 55300 37436 55310 37492
rect 10332 37380 10388 37436
rect 39340 37380 39396 37436
rect 3826 37324 3836 37380
rect 3892 37324 7084 37380
rect 7140 37324 7150 37380
rect 9090 37324 9100 37380
rect 9156 37324 9884 37380
rect 9940 37324 9996 37380
rect 10052 37324 10062 37380
rect 10332 37324 10668 37380
rect 10724 37324 10734 37380
rect 12002 37324 12012 37380
rect 12068 37324 15148 37380
rect 16594 37324 16604 37380
rect 16660 37324 20748 37380
rect 20804 37324 20814 37380
rect 20962 37324 20972 37380
rect 21028 37324 21644 37380
rect 21700 37324 21710 37380
rect 26348 37324 29148 37380
rect 29204 37324 29214 37380
rect 30034 37324 30044 37380
rect 30100 37324 39396 37380
rect 45042 37324 45052 37380
rect 45108 37324 46844 37380
rect 46900 37324 46910 37380
rect 15092 37268 15148 37324
rect 26348 37268 26404 37324
rect 3938 37212 3948 37268
rect 4004 37212 5964 37268
rect 6020 37212 6030 37268
rect 6850 37212 6860 37268
rect 6916 37212 8764 37268
rect 8820 37212 8830 37268
rect 10210 37212 10220 37268
rect 10276 37212 12124 37268
rect 12180 37212 12190 37268
rect 12646 37212 12684 37268
rect 12740 37212 12750 37268
rect 13570 37212 13580 37268
rect 13636 37212 14924 37268
rect 14980 37212 14990 37268
rect 15092 37212 15260 37268
rect 15316 37212 15326 37268
rect 15586 37212 15596 37268
rect 15652 37212 16492 37268
rect 16548 37212 16558 37268
rect 17154 37212 17164 37268
rect 17220 37212 18508 37268
rect 18564 37212 18844 37268
rect 18900 37212 19292 37268
rect 19348 37212 19358 37268
rect 20626 37212 20636 37268
rect 20692 37212 21084 37268
rect 21140 37212 21150 37268
rect 21970 37212 21980 37268
rect 22036 37212 26348 37268
rect 26404 37212 26414 37268
rect 27010 37212 27020 37268
rect 27076 37212 27804 37268
rect 27860 37212 27870 37268
rect 33730 37212 33740 37268
rect 33796 37212 35084 37268
rect 35140 37212 37436 37268
rect 37492 37212 37502 37268
rect 2258 37100 2268 37156
rect 2324 37100 3052 37156
rect 3108 37100 3388 37156
rect 3444 37100 3454 37156
rect 4610 37100 4620 37156
rect 4676 37100 5404 37156
rect 5460 37100 5470 37156
rect 5590 37100 5628 37156
rect 5684 37100 5694 37156
rect 6066 37100 6076 37156
rect 6132 37100 6636 37156
rect 6692 37100 6702 37156
rect 7942 37100 7980 37156
rect 8036 37100 8046 37156
rect 9650 37100 9660 37156
rect 9716 37100 11228 37156
rect 11284 37100 12572 37156
rect 12628 37100 12638 37156
rect 13682 37100 13692 37156
rect 13748 37100 17724 37156
rect 17780 37100 17790 37156
rect 26114 37100 26124 37156
rect 26180 37100 27468 37156
rect 27524 37100 27534 37156
rect 29250 37100 29260 37156
rect 29316 37100 29484 37156
rect 29540 37100 30156 37156
rect 30212 37100 30222 37156
rect 31266 37100 31276 37156
rect 31332 37100 36876 37156
rect 36932 37100 36942 37156
rect 40562 37100 40572 37156
rect 40628 37100 42700 37156
rect 42756 37100 42766 37156
rect 43362 37100 43372 37156
rect 43428 37100 44156 37156
rect 44212 37100 44222 37156
rect 30156 37044 30212 37100
rect 2482 36988 2492 37044
rect 2548 36988 3724 37044
rect 3780 36988 4900 37044
rect 5506 36988 5516 37044
rect 5572 36988 7084 37044
rect 7140 36988 7150 37044
rect 7746 36988 7756 37044
rect 7812 36988 9548 37044
rect 9604 36988 10220 37044
rect 10276 36988 10286 37044
rect 10546 36988 10556 37044
rect 10612 36988 10892 37044
rect 10948 36988 10958 37044
rect 12114 36988 12124 37044
rect 12180 36988 13916 37044
rect 13972 36988 13982 37044
rect 15250 36988 15260 37044
rect 15316 36988 16660 37044
rect 16818 36988 16828 37044
rect 16884 36988 17388 37044
rect 17444 36988 17454 37044
rect 19170 36988 19180 37044
rect 19236 36988 19516 37044
rect 19572 36988 20524 37044
rect 20580 36988 20590 37044
rect 24322 36988 24332 37044
rect 24388 36988 27356 37044
rect 27412 36988 27422 37044
rect 30156 36988 31836 37044
rect 31892 36988 31902 37044
rect 32162 36988 32172 37044
rect 32228 36988 32732 37044
rect 32788 36988 32798 37044
rect 36194 36988 36204 37044
rect 36260 36988 38780 37044
rect 38836 36988 38846 37044
rect 39666 36988 39676 37044
rect 39732 36988 39900 37044
rect 39956 36988 39966 37044
rect 46274 36988 46284 37044
rect 46340 36988 46732 37044
rect 46788 36988 47404 37044
rect 47460 36988 47852 37044
rect 47908 36988 47918 37044
rect 4844 36932 4900 36988
rect 16604 36932 16660 36988
rect 4844 36876 7196 36932
rect 7252 36876 7868 36932
rect 7924 36876 7934 36932
rect 8642 36876 8652 36932
rect 8708 36876 9996 36932
rect 10052 36876 10062 36932
rect 10658 36876 10668 36932
rect 10724 36876 13076 36932
rect 13346 36876 13356 36932
rect 13412 36876 15484 36932
rect 15540 36876 15550 36932
rect 16604 36876 16716 36932
rect 16772 36876 16828 36932
rect 16884 36876 16894 36932
rect 18050 36876 18060 36932
rect 18116 36876 19180 36932
rect 19236 36876 19246 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 5730 36764 5740 36820
rect 5796 36764 6524 36820
rect 6580 36764 11564 36820
rect 11620 36764 11630 36820
rect 13020 36708 13076 36876
rect 13346 36764 13356 36820
rect 13412 36764 13580 36820
rect 13636 36764 16380 36820
rect 16436 36764 16446 36820
rect 18610 36764 18620 36820
rect 18676 36764 18956 36820
rect 19012 36764 19022 36820
rect 6178 36652 6188 36708
rect 6244 36652 8652 36708
rect 8708 36652 8718 36708
rect 9100 36652 10556 36708
rect 10612 36652 10622 36708
rect 10882 36652 10892 36708
rect 10948 36652 12796 36708
rect 12852 36652 12862 36708
rect 13020 36652 13580 36708
rect 13636 36652 13646 36708
rect 13794 36652 13804 36708
rect 13860 36652 14252 36708
rect 14308 36652 14318 36708
rect 14550 36652 14588 36708
rect 14644 36652 14654 36708
rect 16482 36652 16492 36708
rect 16548 36652 16716 36708
rect 16772 36652 20748 36708
rect 20804 36652 20814 36708
rect 2930 36540 2940 36596
rect 2996 36540 7308 36596
rect 7364 36540 7374 36596
rect 7858 36540 7868 36596
rect 7924 36540 8428 36596
rect 8484 36540 8494 36596
rect 9100 36484 9156 36652
rect 9426 36540 9436 36596
rect 9492 36540 9996 36596
rect 10052 36540 10062 36596
rect 10882 36540 10892 36596
rect 10948 36540 14476 36596
rect 14532 36540 14542 36596
rect 15138 36540 15148 36596
rect 15204 36540 17836 36596
rect 17892 36540 17902 36596
rect 18246 36540 18284 36596
rect 18340 36540 18350 36596
rect 1698 36428 1708 36484
rect 1764 36428 2828 36484
rect 2884 36428 3276 36484
rect 3332 36428 3342 36484
rect 4172 36428 9156 36484
rect 9314 36428 9324 36484
rect 9380 36428 10108 36484
rect 10164 36428 10174 36484
rect 10770 36428 10780 36484
rect 10836 36428 11452 36484
rect 11508 36428 11518 36484
rect 12898 36428 12908 36484
rect 12964 36428 15260 36484
rect 15316 36428 16716 36484
rect 16772 36428 16782 36484
rect 18162 36428 18172 36484
rect 18228 36428 22092 36484
rect 22148 36428 22158 36484
rect 1474 36316 1484 36372
rect 1540 36316 3948 36372
rect 4004 36316 4014 36372
rect 4172 36260 4228 36428
rect 26012 36372 26068 36988
rect 38658 36876 38668 36932
rect 38724 36876 38762 36932
rect 42130 36876 42140 36932
rect 42196 36876 42588 36932
rect 42644 36876 42654 36932
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 28354 36652 28364 36708
rect 28420 36652 30380 36708
rect 30436 36652 30446 36708
rect 32162 36652 32172 36708
rect 32228 36652 32956 36708
rect 33012 36652 33404 36708
rect 33460 36652 34300 36708
rect 34356 36652 36428 36708
rect 36484 36652 36494 36708
rect 28578 36540 28588 36596
rect 28644 36540 29484 36596
rect 29540 36540 29550 36596
rect 31938 36540 31948 36596
rect 32004 36540 38668 36596
rect 41682 36540 41692 36596
rect 41748 36540 43820 36596
rect 43876 36540 44380 36596
rect 44436 36540 44446 36596
rect 45042 36540 45052 36596
rect 45108 36540 50204 36596
rect 50260 36540 50270 36596
rect 38612 36484 38668 36540
rect 26562 36428 26572 36484
rect 26628 36428 28028 36484
rect 28084 36428 28476 36484
rect 28532 36428 30268 36484
rect 30324 36428 30334 36484
rect 34850 36428 34860 36484
rect 34916 36428 35308 36484
rect 35364 36428 37884 36484
rect 37940 36428 37950 36484
rect 38612 36428 41356 36484
rect 41412 36428 41804 36484
rect 41860 36428 41870 36484
rect 37884 36372 37940 36428
rect 7410 36316 7420 36372
rect 7476 36316 7644 36372
rect 7700 36316 7710 36372
rect 10434 36316 10444 36372
rect 10500 36316 10556 36372
rect 10612 36316 10622 36372
rect 13794 36316 13804 36372
rect 13860 36316 14140 36372
rect 14196 36316 14206 36372
rect 14438 36316 14476 36372
rect 14532 36316 14542 36372
rect 16818 36316 16828 36372
rect 16884 36316 17052 36372
rect 17108 36316 17118 36372
rect 19954 36316 19964 36372
rect 20020 36316 21868 36372
rect 21924 36316 22428 36372
rect 22484 36316 22494 36372
rect 26002 36316 26012 36372
rect 26068 36316 26078 36372
rect 29586 36316 29596 36372
rect 29652 36316 30156 36372
rect 30212 36316 32060 36372
rect 32116 36316 32844 36372
rect 32900 36316 33012 36372
rect 37884 36316 39564 36372
rect 39620 36316 39630 36372
rect 32956 36260 33012 36316
rect 2258 36204 2268 36260
rect 2324 36204 4228 36260
rect 5058 36204 5068 36260
rect 5124 36204 6412 36260
rect 6468 36204 6478 36260
rect 8988 36204 10892 36260
rect 10948 36204 14364 36260
rect 14420 36204 14924 36260
rect 14980 36204 14990 36260
rect 20850 36204 20860 36260
rect 20916 36204 22876 36260
rect 22932 36204 22942 36260
rect 24434 36204 24444 36260
rect 24500 36204 25900 36260
rect 25956 36204 25966 36260
rect 32386 36204 32396 36260
rect 32452 36204 32620 36260
rect 32676 36204 32686 36260
rect 32956 36204 35980 36260
rect 36036 36204 36652 36260
rect 36708 36204 37436 36260
rect 37492 36204 37502 36260
rect 39890 36204 39900 36260
rect 39956 36204 42252 36260
rect 42308 36204 44156 36260
rect 44212 36204 44222 36260
rect 8988 36148 9044 36204
rect 3378 36092 3388 36148
rect 3444 36092 3836 36148
rect 3892 36092 3902 36148
rect 5842 36092 5852 36148
rect 5908 36092 7644 36148
rect 7700 36092 7710 36148
rect 8530 36092 8540 36148
rect 8596 36092 8988 36148
rect 9044 36092 9054 36148
rect 9314 36092 9324 36148
rect 9380 36092 12012 36148
rect 12068 36092 12684 36148
rect 12740 36092 12750 36148
rect 12898 36092 12908 36148
rect 12964 36092 18060 36148
rect 18116 36092 18126 36148
rect 22194 36092 22204 36148
rect 22260 36092 22270 36148
rect 23986 36092 23996 36148
rect 24052 36092 25228 36148
rect 25284 36092 26124 36148
rect 26180 36092 26190 36148
rect 38332 36092 46620 36148
rect 46676 36092 46686 36148
rect 57698 36092 57708 36148
rect 57764 36092 57774 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 22204 36036 22260 36092
rect 38332 36036 38388 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 57708 36036 57764 36092
rect 3332 35980 9884 36036
rect 9940 35980 9950 36036
rect 16940 35980 17836 36036
rect 17892 35980 18956 36036
rect 19012 35980 19022 36036
rect 20402 35980 20412 36036
rect 20468 35980 20860 36036
rect 20916 35980 22260 36036
rect 25778 35980 25788 36036
rect 25844 35980 35756 36036
rect 35812 35980 36876 36036
rect 36932 35980 38332 36036
rect 38388 35980 38398 36036
rect 42466 35980 42476 36036
rect 42532 35980 47180 36036
rect 47236 35980 47246 36036
rect 57708 35980 58044 36036
rect 58100 35980 58110 36036
rect 3266 35868 3276 35924
rect 3332 35868 3388 35980
rect 16940 35924 16996 35980
rect 7298 35868 7308 35924
rect 7364 35868 8540 35924
rect 8596 35868 8606 35924
rect 13430 35868 13468 35924
rect 13524 35868 13534 35924
rect 15026 35868 15036 35924
rect 15092 35868 15148 35924
rect 15204 35868 15214 35924
rect 16930 35868 16940 35924
rect 16996 35868 17006 35924
rect 17154 35868 17164 35924
rect 17220 35868 18284 35924
rect 18340 35868 18350 35924
rect 19366 35868 19404 35924
rect 19460 35868 20300 35924
rect 20356 35868 20412 35924
rect 20468 35868 20478 35924
rect 20626 35868 20636 35924
rect 20692 35868 20730 35924
rect 22166 35868 22204 35924
rect 22260 35868 23324 35924
rect 23380 35868 23390 35924
rect 24994 35868 25004 35924
rect 25060 35868 26012 35924
rect 26068 35868 26078 35924
rect 32274 35868 32284 35924
rect 32340 35868 32620 35924
rect 32676 35868 32686 35924
rect 33842 35868 33852 35924
rect 33908 35868 34524 35924
rect 34580 35868 34590 35924
rect 34962 35868 34972 35924
rect 35028 35868 42700 35924
rect 42756 35868 44380 35924
rect 44436 35868 44446 35924
rect 45490 35868 45500 35924
rect 45556 35868 46508 35924
rect 46564 35868 47292 35924
rect 47348 35868 47358 35924
rect 50418 35868 50428 35924
rect 50484 35868 51100 35924
rect 51156 35868 51996 35924
rect 52052 35868 56252 35924
rect 56308 35868 56318 35924
rect 2034 35756 2044 35812
rect 2100 35756 10108 35812
rect 10164 35756 10174 35812
rect 13682 35756 13692 35812
rect 13748 35756 15260 35812
rect 15316 35756 16044 35812
rect 16100 35756 16110 35812
rect 16258 35756 16268 35812
rect 16324 35756 16492 35812
rect 16548 35756 16558 35812
rect 17826 35756 17836 35812
rect 17892 35756 20580 35812
rect 30818 35756 30828 35812
rect 30884 35756 32396 35812
rect 32452 35756 32462 35812
rect 41794 35756 41804 35812
rect 41860 35756 43484 35812
rect 43540 35756 43550 35812
rect 44482 35756 44492 35812
rect 44548 35756 44940 35812
rect 44996 35756 45388 35812
rect 45444 35756 45454 35812
rect 45724 35756 45948 35812
rect 46004 35756 46014 35812
rect 53890 35756 53900 35812
rect 53956 35756 54796 35812
rect 54852 35756 54862 35812
rect 20524 35700 20580 35756
rect 4722 35644 4732 35700
rect 4788 35644 5740 35700
rect 5796 35644 5806 35700
rect 9538 35644 9548 35700
rect 9604 35644 10780 35700
rect 10836 35644 11788 35700
rect 11844 35644 11854 35700
rect 12338 35644 12348 35700
rect 12404 35644 13356 35700
rect 13412 35644 13422 35700
rect 14242 35644 14252 35700
rect 14308 35644 14588 35700
rect 14644 35644 16604 35700
rect 16660 35644 16670 35700
rect 16818 35644 16828 35700
rect 16884 35644 17388 35700
rect 17444 35644 17454 35700
rect 17602 35644 17612 35700
rect 17668 35644 18284 35700
rect 18340 35644 19068 35700
rect 19124 35644 19134 35700
rect 20514 35644 20524 35700
rect 20580 35644 21420 35700
rect 21476 35644 21486 35700
rect 25554 35644 25564 35700
rect 25620 35644 25788 35700
rect 25844 35644 25854 35700
rect 28914 35644 28924 35700
rect 28980 35644 31052 35700
rect 31108 35644 31836 35700
rect 31892 35644 33404 35700
rect 33460 35644 33470 35700
rect 33954 35644 33964 35700
rect 34020 35644 34636 35700
rect 34692 35644 34702 35700
rect 37314 35644 37324 35700
rect 37380 35644 39900 35700
rect 39956 35644 39966 35700
rect 40786 35644 40796 35700
rect 40852 35644 41132 35700
rect 41188 35644 42028 35700
rect 42084 35644 42094 35700
rect 3826 35532 3836 35588
rect 3892 35532 5516 35588
rect 5572 35532 5582 35588
rect 7634 35532 7644 35588
rect 7700 35532 13804 35588
rect 13860 35532 13870 35588
rect 15474 35532 15484 35588
rect 15540 35532 20076 35588
rect 20132 35532 20142 35588
rect 20402 35532 20412 35588
rect 20468 35532 21084 35588
rect 21140 35532 21150 35588
rect 21522 35532 21532 35588
rect 21588 35532 22092 35588
rect 22148 35532 22158 35588
rect 22642 35532 22652 35588
rect 22708 35532 25788 35588
rect 25844 35532 26348 35588
rect 26404 35532 26796 35588
rect 26852 35532 26862 35588
rect 27570 35532 27580 35588
rect 27636 35532 28252 35588
rect 28308 35532 28812 35588
rect 28868 35532 30380 35588
rect 30436 35532 30446 35588
rect 35074 35532 35084 35588
rect 35140 35532 36204 35588
rect 36260 35532 36270 35588
rect 37090 35532 37100 35588
rect 37156 35532 39004 35588
rect 39060 35532 39228 35588
rect 39284 35532 39294 35588
rect 45724 35476 45780 35756
rect 48290 35644 48300 35700
rect 48356 35644 53004 35700
rect 53060 35644 53676 35700
rect 53732 35644 53742 35700
rect 55570 35644 55580 35700
rect 55636 35644 56364 35700
rect 56420 35644 56430 35700
rect 56690 35644 56700 35700
rect 56756 35644 57932 35700
rect 57988 35644 57998 35700
rect 45938 35532 45948 35588
rect 46004 35532 46172 35588
rect 46228 35532 46238 35588
rect 47730 35532 47740 35588
rect 47796 35532 49420 35588
rect 49476 35532 49980 35588
rect 50036 35532 50046 35588
rect 3686 35420 3724 35476
rect 3780 35420 3790 35476
rect 4172 35420 9324 35476
rect 9380 35420 9390 35476
rect 10098 35420 10108 35476
rect 10164 35420 16940 35476
rect 16996 35420 19180 35476
rect 19236 35420 19246 35476
rect 26786 35420 26796 35476
rect 26852 35420 27692 35476
rect 27748 35420 29484 35476
rect 29540 35420 29550 35476
rect 30482 35420 30492 35476
rect 30548 35420 33628 35476
rect 33684 35420 33694 35476
rect 35522 35420 35532 35476
rect 35588 35420 36988 35476
rect 37044 35420 37054 35476
rect 39554 35420 39564 35476
rect 39620 35420 40124 35476
rect 40180 35420 40460 35476
rect 40516 35420 42476 35476
rect 42532 35420 43036 35476
rect 43092 35420 43102 35476
rect 45714 35420 45724 35476
rect 45780 35420 45790 35476
rect 4172 35364 4228 35420
rect 3378 35308 3388 35364
rect 3444 35308 4228 35364
rect 4946 35308 4956 35364
rect 5012 35308 5516 35364
rect 5572 35308 5964 35364
rect 6020 35308 6030 35364
rect 9202 35308 9212 35364
rect 9268 35308 10332 35364
rect 10388 35308 10398 35364
rect 13570 35308 13580 35364
rect 13636 35308 13916 35364
rect 13972 35308 13982 35364
rect 26450 35308 26460 35364
rect 26516 35308 27468 35364
rect 27524 35308 29596 35364
rect 29652 35308 29662 35364
rect 35746 35308 35756 35364
rect 35812 35308 37772 35364
rect 37828 35308 37838 35364
rect 43698 35308 43708 35364
rect 43764 35308 47740 35364
rect 47796 35308 47806 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 2370 35196 2380 35252
rect 2436 35196 3500 35252
rect 3556 35196 3566 35252
rect 6962 35196 6972 35252
rect 7028 35196 9772 35252
rect 9828 35196 9838 35252
rect 10994 35196 11004 35252
rect 11060 35196 11900 35252
rect 11956 35196 11966 35252
rect 13458 35196 13468 35252
rect 13524 35196 13804 35252
rect 13860 35196 13870 35252
rect 17490 35196 17500 35252
rect 17556 35196 18844 35252
rect 18900 35196 18910 35252
rect 25666 35196 25676 35252
rect 25732 35196 26236 35252
rect 26292 35196 26302 35252
rect 31602 35196 31612 35252
rect 31668 35196 33516 35252
rect 33572 35196 33582 35252
rect 47506 35196 47516 35252
rect 47572 35196 53228 35252
rect 53284 35196 53294 35252
rect 1810 35084 1820 35140
rect 1876 35084 3388 35140
rect 3332 35028 3388 35084
rect 4172 35084 6636 35140
rect 6692 35084 6702 35140
rect 7186 35084 7196 35140
rect 7252 35084 8204 35140
rect 8260 35084 8270 35140
rect 12002 35084 12012 35140
rect 12068 35084 14252 35140
rect 14308 35084 14318 35140
rect 15474 35084 15484 35140
rect 15540 35084 16604 35140
rect 16660 35084 18508 35140
rect 18564 35084 18574 35140
rect 19282 35084 19292 35140
rect 19348 35084 20076 35140
rect 20132 35084 20142 35140
rect 27010 35084 27020 35140
rect 27076 35084 34692 35140
rect 36754 35084 36764 35140
rect 36820 35084 36830 35140
rect 37538 35084 37548 35140
rect 37604 35084 38108 35140
rect 38164 35084 38174 35140
rect 41682 35084 41692 35140
rect 41748 35084 43932 35140
rect 43988 35084 43998 35140
rect 49074 35084 49084 35140
rect 49140 35084 49532 35140
rect 49588 35084 49598 35140
rect 4172 35028 4228 35084
rect 6636 35028 6692 35084
rect 34636 35028 34692 35084
rect 36764 35028 36820 35084
rect 37548 35028 37604 35084
rect 3332 34972 4228 35028
rect 4386 34972 4396 35028
rect 4452 34972 5404 35028
rect 5460 34972 5470 35028
rect 6636 34972 8764 35028
rect 8820 34972 9492 35028
rect 9874 34972 9884 35028
rect 9940 34972 12124 35028
rect 12180 34972 12190 35028
rect 13122 34972 13132 35028
rect 13188 34972 16044 35028
rect 16100 34972 17948 35028
rect 18004 34972 18014 35028
rect 18386 34972 18396 35028
rect 18452 34972 20524 35028
rect 20580 34972 20590 35028
rect 25666 34972 25676 35028
rect 25732 34972 31276 35028
rect 31332 34972 31342 35028
rect 32386 34972 32396 35028
rect 32452 34972 33684 35028
rect 34636 34972 37604 35028
rect 38882 34972 38892 35028
rect 38948 34972 40796 35028
rect 40852 34972 40862 35028
rect 47618 34972 47628 35028
rect 47684 34972 48188 35028
rect 48244 34972 48972 35028
rect 49028 34972 49038 35028
rect 9436 34916 9492 34972
rect 33628 34916 33684 34972
rect 3378 34860 3388 34916
rect 3444 34860 3482 34916
rect 5394 34860 5404 34916
rect 5460 34860 5516 34916
rect 5572 34860 5582 34916
rect 6290 34860 6300 34916
rect 6356 34860 7308 34916
rect 7364 34860 7374 34916
rect 9436 34860 10220 34916
rect 10276 34860 11004 34916
rect 11060 34860 11070 34916
rect 14242 34860 14252 34916
rect 14308 34860 15932 34916
rect 15988 34860 15998 34916
rect 17490 34860 17500 34916
rect 17556 34860 18956 34916
rect 19012 34860 19022 34916
rect 19618 34860 19628 34916
rect 19684 34860 20076 34916
rect 20132 34860 20142 34916
rect 30034 34860 30044 34916
rect 30100 34860 31052 34916
rect 31108 34860 31500 34916
rect 31556 34860 32844 34916
rect 32900 34860 33180 34916
rect 33236 34860 33246 34916
rect 33618 34860 33628 34916
rect 33684 34860 34524 34916
rect 34580 34860 34590 34916
rect 34850 34860 34860 34916
rect 34916 34860 35868 34916
rect 35924 34860 35934 34916
rect 37874 34860 37884 34916
rect 37940 34860 39116 34916
rect 39172 34860 39182 34916
rect 42018 34860 42028 34916
rect 42084 34860 42588 34916
rect 42644 34860 42654 34916
rect 50372 34860 51212 34916
rect 51268 34860 51660 34916
rect 51716 34860 52108 34916
rect 52164 34860 52174 34916
rect 52546 34860 52556 34916
rect 52612 34860 53564 34916
rect 53620 34860 54012 34916
rect 54068 34860 54078 34916
rect 34524 34804 34580 34860
rect 50372 34804 50428 34860
rect 1586 34748 1596 34804
rect 1652 34748 4844 34804
rect 4900 34748 4910 34804
rect 6066 34748 6076 34804
rect 6132 34748 7980 34804
rect 8036 34748 8046 34804
rect 14466 34748 14476 34804
rect 14532 34748 17052 34804
rect 17108 34748 19180 34804
rect 19236 34748 20300 34804
rect 20356 34748 20366 34804
rect 21634 34748 21644 34804
rect 21700 34748 24444 34804
rect 24500 34748 24510 34804
rect 29698 34748 29708 34804
rect 29764 34748 31164 34804
rect 31220 34748 32508 34804
rect 32564 34748 32574 34804
rect 34524 34748 36092 34804
rect 36148 34748 36158 34804
rect 42690 34748 42700 34804
rect 42756 34748 50428 34804
rect 50866 34748 50876 34804
rect 50932 34748 53788 34804
rect 53844 34748 53854 34804
rect 2370 34636 2380 34692
rect 2436 34636 2828 34692
rect 2884 34636 4508 34692
rect 4564 34636 5964 34692
rect 6020 34636 7196 34692
rect 7252 34636 7262 34692
rect 8054 34636 8092 34692
rect 8148 34636 8158 34692
rect 10658 34636 10668 34692
rect 10724 34636 12572 34692
rect 12628 34636 13020 34692
rect 13076 34636 13086 34692
rect 15138 34636 15148 34692
rect 15204 34636 15242 34692
rect 16818 34636 16828 34692
rect 16884 34636 17276 34692
rect 17332 34636 17948 34692
rect 18004 34636 19404 34692
rect 19460 34636 20860 34692
rect 20916 34636 21420 34692
rect 21476 34636 21486 34692
rect 21634 34636 21644 34692
rect 21700 34636 21980 34692
rect 22036 34636 22046 34692
rect 26338 34636 26348 34692
rect 26404 34636 27804 34692
rect 27860 34636 27870 34692
rect 28578 34636 28588 34692
rect 28644 34636 34524 34692
rect 34580 34636 35084 34692
rect 35140 34636 35150 34692
rect 38994 34636 39004 34692
rect 39060 34636 39900 34692
rect 39956 34636 42028 34692
rect 42084 34636 42094 34692
rect 43810 34636 43820 34692
rect 43876 34636 44044 34692
rect 44100 34636 44380 34692
rect 44436 34636 44940 34692
rect 44996 34636 45006 34692
rect 5282 34524 5292 34580
rect 5348 34524 5516 34580
rect 5572 34524 5582 34580
rect 6514 34524 6524 34580
rect 6580 34524 11676 34580
rect 11732 34524 11900 34580
rect 11956 34524 16268 34580
rect 16324 34524 16334 34580
rect 32050 34524 32060 34580
rect 32116 34524 38556 34580
rect 38612 34524 38622 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 2034 34412 2044 34468
rect 2100 34412 4284 34468
rect 4340 34412 4350 34468
rect 5366 34412 5404 34468
rect 5460 34412 5470 34468
rect 5730 34412 5740 34468
rect 5796 34412 6412 34468
rect 6468 34412 8540 34468
rect 8596 34412 8606 34468
rect 17602 34412 17612 34468
rect 17668 34412 18620 34468
rect 18676 34412 18686 34468
rect 23538 34412 23548 34468
rect 23604 34412 23884 34468
rect 23940 34412 24332 34468
rect 24388 34412 24398 34468
rect 24770 34412 24780 34468
rect 24836 34412 25340 34468
rect 25396 34412 25406 34468
rect 34290 34412 34300 34468
rect 34356 34412 34860 34468
rect 34916 34412 34926 34468
rect 35186 34412 35196 34468
rect 35252 34412 45836 34468
rect 45892 34412 45902 34468
rect 4096 34300 4172 34356
rect 4228 34300 9212 34356
rect 9268 34300 9278 34356
rect 11330 34300 11340 34356
rect 11396 34300 11900 34356
rect 11956 34300 11966 34356
rect 12226 34300 12236 34356
rect 12292 34300 13692 34356
rect 13748 34300 13758 34356
rect 24098 34300 24108 34356
rect 24164 34300 26012 34356
rect 26068 34300 26078 34356
rect 28914 34300 28924 34356
rect 28980 34300 36652 34356
rect 36708 34300 37324 34356
rect 37380 34300 37390 34356
rect 52098 34300 52108 34356
rect 52164 34300 52668 34356
rect 52724 34300 52734 34356
rect 26012 34244 26068 34300
rect 2258 34188 2268 34244
rect 2324 34188 5180 34244
rect 5236 34188 5964 34244
rect 6020 34188 6030 34244
rect 6514 34188 6524 34244
rect 6580 34188 6860 34244
rect 6916 34188 6926 34244
rect 7074 34188 7084 34244
rect 7140 34188 8092 34244
rect 8148 34188 9100 34244
rect 9156 34188 9996 34244
rect 10052 34188 10062 34244
rect 11778 34188 11788 34244
rect 11844 34188 12796 34244
rect 12852 34188 16828 34244
rect 16884 34188 16894 34244
rect 26012 34188 26460 34244
rect 26516 34188 26526 34244
rect 36194 34188 36204 34244
rect 36260 34188 36270 34244
rect 37538 34188 37548 34244
rect 37604 34188 38220 34244
rect 38276 34188 39900 34244
rect 39956 34188 40796 34244
rect 40852 34188 40862 34244
rect 41234 34188 41244 34244
rect 41300 34188 42588 34244
rect 42644 34188 42812 34244
rect 42868 34188 42878 34244
rect 46946 34188 46956 34244
rect 47012 34188 47404 34244
rect 47460 34188 47852 34244
rect 47908 34188 47918 34244
rect 36204 34132 36260 34188
rect 3714 34076 3724 34132
rect 3780 34076 6412 34132
rect 6468 34076 6478 34132
rect 6738 34076 6748 34132
rect 6804 34076 10108 34132
rect 10164 34076 10174 34132
rect 10742 34076 10780 34132
rect 10836 34076 10846 34132
rect 14802 34076 14812 34132
rect 14868 34076 15820 34132
rect 15876 34076 15886 34132
rect 20626 34076 20636 34132
rect 20692 34076 21644 34132
rect 21700 34076 21710 34132
rect 24434 34076 24444 34132
rect 24500 34076 27468 34132
rect 27524 34076 27534 34132
rect 29922 34076 29932 34132
rect 29988 34076 31724 34132
rect 31780 34076 31790 34132
rect 35074 34076 35084 34132
rect 35140 34076 35756 34132
rect 35812 34076 36764 34132
rect 36820 34076 36830 34132
rect 38322 34076 38332 34132
rect 38388 34076 39452 34132
rect 39508 34076 41468 34132
rect 41524 34076 41534 34132
rect 48962 34076 48972 34132
rect 49028 34076 49420 34132
rect 49476 34076 49980 34132
rect 50036 34076 50046 34132
rect 6412 34020 6468 34076
rect 1922 33964 1932 34020
rect 1988 33964 2156 34020
rect 2212 33964 3612 34020
rect 3668 33964 3678 34020
rect 4060 33964 4172 34020
rect 4228 33964 4238 34020
rect 6412 33964 10668 34020
rect 10724 33964 10734 34020
rect 14018 33964 14028 34020
rect 14084 33964 15148 34020
rect 15204 33964 16044 34020
rect 16100 33964 16110 34020
rect 17378 33964 17388 34020
rect 17444 33964 17836 34020
rect 17892 33964 18732 34020
rect 18788 33964 19180 34020
rect 19236 33964 19246 34020
rect 19730 33964 19740 34020
rect 19796 33964 20524 34020
rect 20580 33964 20590 34020
rect 21298 33964 21308 34020
rect 21364 33964 22764 34020
rect 22820 33964 22830 34020
rect 23062 33964 23100 34020
rect 23156 33964 24220 34020
rect 24276 33964 24286 34020
rect 24882 33964 24892 34020
rect 24948 33964 27244 34020
rect 27300 33964 27310 34020
rect 32274 33964 32284 34020
rect 32340 33964 41916 34020
rect 41972 33964 42364 34020
rect 42420 33964 43820 34020
rect 43876 33964 43886 34020
rect 44482 33964 44492 34020
rect 44548 33964 47628 34020
rect 47684 33964 47694 34020
rect 4060 33908 4116 33964
rect 1026 33852 1036 33908
rect 1092 33852 4116 33908
rect 4274 33852 4284 33908
rect 4340 33852 5292 33908
rect 5348 33852 6412 33908
rect 6468 33852 6478 33908
rect 7970 33852 7980 33908
rect 8036 33852 10108 33908
rect 10164 33852 10174 33908
rect 13010 33852 13020 33908
rect 13076 33852 18508 33908
rect 18564 33852 19516 33908
rect 19572 33852 19582 33908
rect 20178 33852 20188 33908
rect 20244 33852 21644 33908
rect 21700 33852 21710 33908
rect 22614 33852 22652 33908
rect 22708 33852 22718 33908
rect 25526 33852 25564 33908
rect 25620 33852 25630 33908
rect 26450 33852 26460 33908
rect 26516 33852 27132 33908
rect 27188 33852 28476 33908
rect 28532 33852 28542 33908
rect 29810 33852 29820 33908
rect 29876 33852 30604 33908
rect 30660 33852 30670 33908
rect 32498 33852 32508 33908
rect 32564 33852 45500 33908
rect 45556 33852 46060 33908
rect 46116 33852 46126 33908
rect 4844 33740 8428 33796
rect 8484 33740 8988 33796
rect 9044 33740 13244 33796
rect 13300 33740 13468 33796
rect 13524 33740 13692 33796
rect 13748 33740 13758 33796
rect 16930 33740 16940 33796
rect 16996 33740 18396 33796
rect 18452 33740 18462 33796
rect 25638 33740 25676 33796
rect 25732 33740 25742 33796
rect 30370 33740 30380 33796
rect 30436 33740 32172 33796
rect 32228 33740 32732 33796
rect 32788 33740 32798 33796
rect 39330 33740 39340 33796
rect 39396 33740 40012 33796
rect 40068 33740 40460 33796
rect 40516 33740 40526 33796
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 3602 33628 3612 33684
rect 3668 33628 3836 33684
rect 3892 33628 4340 33684
rect 4284 33572 4340 33628
rect 4844 33572 4900 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 5058 33628 5068 33684
rect 5124 33628 10780 33684
rect 10836 33628 12348 33684
rect 12404 33628 12414 33684
rect 20514 33628 20524 33684
rect 20580 33628 23212 33684
rect 23268 33628 23278 33684
rect 23426 33628 23436 33684
rect 23492 33628 23996 33684
rect 24052 33628 24062 33684
rect 31826 33628 31836 33684
rect 31892 33628 32396 33684
rect 32452 33628 32462 33684
rect 37538 33628 37548 33684
rect 37604 33628 37614 33684
rect 38098 33628 38108 33684
rect 38164 33628 41468 33684
rect 41524 33628 41534 33684
rect 3378 33516 3388 33572
rect 3444 33516 4060 33572
rect 4116 33516 4126 33572
rect 4284 33516 4900 33572
rect 5506 33516 5516 33572
rect 5572 33516 6076 33572
rect 6132 33516 6142 33572
rect 8642 33516 8652 33572
rect 8708 33516 12516 33572
rect 12898 33516 12908 33572
rect 12964 33516 16156 33572
rect 16212 33516 16222 33572
rect 17602 33516 17612 33572
rect 17668 33516 17678 33572
rect 19058 33516 19068 33572
rect 19124 33516 21084 33572
rect 21140 33516 21150 33572
rect 26786 33516 26796 33572
rect 26852 33516 27356 33572
rect 27412 33516 27422 33572
rect 12460 33460 12516 33516
rect 17612 33460 17668 33516
rect 37548 33460 37604 33628
rect 39106 33516 39116 33572
rect 39172 33516 41692 33572
rect 41748 33516 41758 33572
rect 3938 33404 3948 33460
rect 4004 33404 6972 33460
rect 7028 33404 7038 33460
rect 8082 33404 8092 33460
rect 8148 33404 8876 33460
rect 8932 33404 8942 33460
rect 12460 33404 15148 33460
rect 15204 33404 15596 33460
rect 15652 33404 15662 33460
rect 16258 33404 16268 33460
rect 16324 33404 17668 33460
rect 18498 33404 18508 33460
rect 18564 33404 19516 33460
rect 19572 33404 19628 33460
rect 19684 33404 19694 33460
rect 20374 33404 20412 33460
rect 20468 33404 22092 33460
rect 22148 33404 22158 33460
rect 22530 33404 22540 33460
rect 22596 33404 37604 33460
rect 38546 33404 38556 33460
rect 38612 33404 40236 33460
rect 40292 33404 40302 33460
rect 54450 33404 54460 33460
rect 54516 33404 56476 33460
rect 56532 33404 56542 33460
rect 3490 33292 3500 33348
rect 3556 33292 5180 33348
rect 5236 33292 5628 33348
rect 5684 33292 7532 33348
rect 7588 33292 7598 33348
rect 7746 33292 7756 33348
rect 7812 33292 9660 33348
rect 9716 33292 9726 33348
rect 12450 33292 12460 33348
rect 12516 33292 15260 33348
rect 15316 33292 15326 33348
rect 16044 33292 16380 33348
rect 16436 33292 16446 33348
rect 17826 33292 17836 33348
rect 17892 33292 18396 33348
rect 18452 33292 18462 33348
rect 22866 33292 22876 33348
rect 22932 33292 32620 33348
rect 32676 33292 32686 33348
rect 35970 33292 35980 33348
rect 36036 33292 37436 33348
rect 37492 33292 37502 33348
rect 16044 33236 16100 33292
rect 4274 33180 4284 33236
rect 4340 33180 4844 33236
rect 4900 33180 4910 33236
rect 6402 33180 6412 33236
rect 6468 33180 7868 33236
rect 7924 33180 7934 33236
rect 13794 33180 13804 33236
rect 13860 33180 14252 33236
rect 14308 33180 14318 33236
rect 16034 33180 16044 33236
rect 16100 33180 16110 33236
rect 18610 33180 18620 33236
rect 18676 33180 24332 33236
rect 24388 33180 24398 33236
rect 26898 33180 26908 33236
rect 26964 33180 29036 33236
rect 29092 33180 29102 33236
rect 30370 33180 30380 33236
rect 30436 33180 36316 33236
rect 36372 33180 39004 33236
rect 39060 33180 39564 33236
rect 39620 33180 39630 33236
rect 39900 33180 40908 33236
rect 40964 33180 40974 33236
rect 39900 33124 39956 33180
rect 2818 33068 2828 33124
rect 2884 33068 5292 33124
rect 5348 33068 6076 33124
rect 6132 33068 6142 33124
rect 9202 33068 9212 33124
rect 9268 33068 16716 33124
rect 16772 33068 16782 33124
rect 17042 33068 17052 33124
rect 17108 33068 17724 33124
rect 17780 33068 17790 33124
rect 18274 33068 18284 33124
rect 18340 33068 18956 33124
rect 19012 33068 19022 33124
rect 19730 33068 19740 33124
rect 19796 33068 21308 33124
rect 21364 33068 21374 33124
rect 22642 33068 22652 33124
rect 22708 33068 23100 33124
rect 23156 33068 23166 33124
rect 31266 33068 31276 33124
rect 31332 33068 33404 33124
rect 33460 33068 33470 33124
rect 36418 33068 36428 33124
rect 36484 33068 39900 33124
rect 39956 33068 39966 33124
rect 40114 33068 40124 33124
rect 40180 33068 41020 33124
rect 41076 33068 41086 33124
rect 46050 33068 46060 33124
rect 46116 33068 46508 33124
rect 46564 33068 47068 33124
rect 47124 33068 47134 33124
rect 22876 33012 22932 33068
rect 3332 32956 12572 33012
rect 12628 32956 12638 33012
rect 14914 32956 14924 33012
rect 14980 32956 19404 33012
rect 19460 32956 19470 33012
rect 22866 32956 22876 33012
rect 22932 32956 22942 33012
rect 32498 32956 32508 33012
rect 32564 32956 44380 33012
rect 44436 32956 44828 33012
rect 44884 32956 44894 33012
rect 3332 32900 3388 32956
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 1474 32844 1484 32900
rect 1540 32844 1932 32900
rect 1988 32844 3388 32900
rect 5292 32844 7700 32900
rect 7858 32844 7868 32900
rect 7924 32844 8540 32900
rect 8596 32844 12124 32900
rect 12180 32844 13916 32900
rect 13972 32844 13982 32900
rect 20626 32844 20636 32900
rect 20692 32844 26236 32900
rect 26292 32844 26302 32900
rect 38882 32844 38892 32900
rect 38948 32844 39116 32900
rect 39172 32844 39676 32900
rect 39732 32844 42140 32900
rect 42196 32844 44044 32900
rect 44100 32844 44110 32900
rect 5292 32788 5348 32844
rect 7644 32788 7700 32844
rect 2482 32732 2492 32788
rect 2548 32732 5348 32788
rect 5506 32732 5516 32788
rect 5572 32732 6972 32788
rect 7028 32732 7038 32788
rect 7644 32732 8428 32788
rect 8484 32732 9548 32788
rect 9604 32732 9614 32788
rect 13794 32732 13804 32788
rect 13860 32732 14364 32788
rect 14420 32732 15036 32788
rect 15092 32732 15102 32788
rect 15810 32732 15820 32788
rect 15876 32732 17388 32788
rect 17444 32732 17454 32788
rect 17714 32732 17724 32788
rect 17780 32732 18396 32788
rect 18452 32732 18462 32788
rect 18946 32732 18956 32788
rect 19012 32732 20860 32788
rect 20916 32732 22092 32788
rect 22148 32732 22158 32788
rect 26534 32732 26572 32788
rect 26628 32732 26638 32788
rect 35522 32732 35532 32788
rect 35588 32732 39340 32788
rect 39396 32732 39406 32788
rect 40226 32732 40236 32788
rect 40292 32732 43820 32788
rect 43876 32732 43886 32788
rect 49186 32732 49196 32788
rect 49252 32732 49868 32788
rect 49924 32732 50428 32788
rect 50372 32676 50428 32732
rect 3602 32620 3612 32676
rect 3668 32620 6188 32676
rect 6244 32620 6254 32676
rect 7634 32620 7644 32676
rect 7700 32620 10780 32676
rect 10836 32620 10846 32676
rect 11442 32620 11452 32676
rect 11508 32620 13468 32676
rect 13524 32620 13534 32676
rect 14354 32620 14364 32676
rect 14420 32620 20300 32676
rect 20356 32620 20366 32676
rect 21298 32620 21308 32676
rect 21364 32620 21756 32676
rect 21812 32620 21822 32676
rect 23436 32620 23548 32676
rect 23604 32620 23614 32676
rect 31378 32620 31388 32676
rect 31444 32620 38332 32676
rect 38388 32620 43036 32676
rect 43092 32620 44492 32676
rect 44548 32620 44558 32676
rect 50372 32620 50820 32676
rect 23436 32564 23492 32620
rect 50764 32564 50820 32620
rect 3826 32508 3836 32564
rect 3892 32508 4284 32564
rect 4340 32508 4350 32564
rect 4498 32508 4508 32564
rect 4564 32508 5628 32564
rect 5684 32508 5694 32564
rect 9090 32508 9100 32564
rect 9156 32508 12684 32564
rect 12740 32508 12750 32564
rect 13542 32508 13580 32564
rect 13636 32508 13646 32564
rect 16258 32508 16268 32564
rect 16324 32508 23492 32564
rect 24322 32508 24332 32564
rect 24388 32508 26012 32564
rect 26068 32508 26078 32564
rect 28130 32508 28140 32564
rect 28196 32508 28700 32564
rect 28756 32508 29596 32564
rect 29652 32508 29662 32564
rect 30818 32508 30828 32564
rect 30884 32508 35308 32564
rect 35364 32508 36988 32564
rect 37044 32508 38388 32564
rect 38546 32508 38556 32564
rect 38612 32508 39228 32564
rect 39284 32508 39294 32564
rect 41906 32508 41916 32564
rect 41972 32508 42924 32564
rect 42980 32508 42990 32564
rect 49970 32508 49980 32564
rect 50036 32508 50428 32564
rect 50484 32508 50494 32564
rect 50754 32508 50764 32564
rect 50820 32508 51212 32564
rect 51268 32508 51278 32564
rect 54786 32508 54796 32564
rect 54852 32508 55356 32564
rect 55412 32508 55422 32564
rect 56914 32508 56924 32564
rect 56980 32508 57820 32564
rect 57876 32508 57886 32564
rect 38332 32452 38388 32508
rect 2930 32396 2940 32452
rect 2996 32396 8092 32452
rect 8148 32396 8158 32452
rect 11218 32396 11228 32452
rect 11284 32396 11676 32452
rect 11732 32396 11742 32452
rect 12338 32396 12348 32452
rect 12404 32396 15708 32452
rect 15764 32396 15820 32452
rect 15876 32396 15886 32452
rect 16146 32396 16156 32452
rect 16212 32396 16492 32452
rect 16548 32396 17948 32452
rect 18004 32396 18014 32452
rect 19394 32396 19404 32452
rect 19460 32396 21868 32452
rect 21924 32396 21934 32452
rect 22082 32396 22092 32452
rect 22148 32396 23212 32452
rect 23268 32396 23278 32452
rect 24098 32396 24108 32452
rect 24164 32396 25116 32452
rect 25172 32396 26908 32452
rect 26964 32396 26974 32452
rect 27906 32396 27916 32452
rect 27972 32396 29932 32452
rect 29988 32396 29998 32452
rect 32610 32396 32620 32452
rect 32676 32396 33628 32452
rect 33684 32396 35644 32452
rect 35700 32396 36316 32452
rect 36372 32396 36382 32452
rect 38332 32396 38444 32452
rect 38500 32396 38510 32452
rect 38658 32396 38668 32452
rect 38724 32396 40012 32452
rect 40068 32396 40078 32452
rect 44930 32396 44940 32452
rect 44996 32396 45500 32452
rect 45556 32396 45566 32452
rect 3378 32284 3388 32340
rect 3444 32284 4284 32340
rect 4340 32284 13580 32340
rect 13636 32284 13646 32340
rect 16818 32284 16828 32340
rect 16884 32284 17724 32340
rect 17780 32284 17790 32340
rect 18050 32284 18060 32340
rect 18116 32284 18620 32340
rect 18676 32284 18686 32340
rect 19954 32284 19964 32340
rect 20020 32284 24556 32340
rect 24612 32284 24622 32340
rect 24994 32284 25004 32340
rect 25060 32284 26908 32340
rect 27010 32284 27020 32340
rect 27076 32284 27580 32340
rect 27636 32284 27692 32340
rect 27748 32284 27758 32340
rect 33506 32284 33516 32340
rect 33572 32284 34524 32340
rect 34580 32284 34590 32340
rect 36082 32284 36092 32340
rect 36148 32284 37436 32340
rect 37492 32284 37502 32340
rect 38546 32284 38556 32340
rect 38612 32284 40684 32340
rect 40740 32284 40750 32340
rect 43810 32284 43820 32340
rect 43876 32284 45164 32340
rect 45220 32284 45230 32340
rect 24556 32228 24612 32284
rect 26852 32228 26908 32284
rect 4834 32172 4844 32228
rect 4900 32172 5516 32228
rect 5572 32172 5582 32228
rect 6962 32172 6972 32228
rect 7028 32172 14700 32228
rect 14756 32172 14766 32228
rect 24556 32172 25900 32228
rect 25956 32172 25966 32228
rect 26852 32172 28252 32228
rect 28308 32172 28318 32228
rect 33394 32172 33404 32228
rect 33460 32172 34412 32228
rect 34468 32172 34478 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 12562 32060 12572 32116
rect 12628 32060 14476 32116
rect 14532 32060 14924 32116
rect 14980 32060 14990 32116
rect 18498 32060 18508 32116
rect 18564 32060 19180 32116
rect 19236 32060 19246 32116
rect 20178 32060 20188 32116
rect 20244 32060 20972 32116
rect 21028 32060 21038 32116
rect 34066 32060 34076 32116
rect 34132 32060 34636 32116
rect 34692 32060 34702 32116
rect 2370 31948 2380 32004
rect 2436 31948 3500 32004
rect 3556 31948 3566 32004
rect 6066 31948 6076 32004
rect 6132 31948 7196 32004
rect 7252 31948 9212 32004
rect 9268 31948 9884 32004
rect 9940 31948 10220 32004
rect 10276 31948 10286 32004
rect 15092 31892 15148 32004
rect 15204 31948 15214 32004
rect 15474 31948 15484 32004
rect 15540 31948 16828 32004
rect 16884 31948 18844 32004
rect 18900 31948 20076 32004
rect 20132 31948 20524 32004
rect 20580 31948 20590 32004
rect 23100 31948 25452 32004
rect 25508 31948 25518 32004
rect 25778 31948 25788 32004
rect 25844 31948 35532 32004
rect 35588 31948 35598 32004
rect 38098 31948 38108 32004
rect 38164 31948 43820 32004
rect 43876 31948 44828 32004
rect 44884 31948 44894 32004
rect 53890 31948 53900 32004
rect 53956 31948 57372 32004
rect 57428 31948 57438 32004
rect 23100 31892 23156 31948
rect 2258 31836 2268 31892
rect 2324 31836 3388 31892
rect 3602 31836 3612 31892
rect 3668 31836 3724 31892
rect 3780 31836 3790 31892
rect 5058 31836 5068 31892
rect 5124 31836 10108 31892
rect 10164 31836 12012 31892
rect 12068 31836 12078 31892
rect 13682 31836 13692 31892
rect 13748 31836 15148 31892
rect 17714 31836 17724 31892
rect 17780 31836 18508 31892
rect 18564 31836 18574 31892
rect 19058 31836 19068 31892
rect 19124 31836 20748 31892
rect 20804 31836 21756 31892
rect 21812 31836 21822 31892
rect 22194 31836 22204 31892
rect 22260 31836 22876 31892
rect 22932 31836 22942 31892
rect 23090 31836 23100 31892
rect 23156 31836 23166 31892
rect 24434 31836 24444 31892
rect 24500 31836 31388 31892
rect 31444 31836 31454 31892
rect 34962 31836 34972 31892
rect 35028 31836 35196 31892
rect 35252 31836 35262 31892
rect 40002 31836 40012 31892
rect 40068 31836 40236 31892
rect 40292 31836 41916 31892
rect 41972 31836 41982 31892
rect 48514 31836 48524 31892
rect 48580 31836 54460 31892
rect 54516 31836 54796 31892
rect 54852 31836 55132 31892
rect 55188 31836 55468 31892
rect 55524 31836 55534 31892
rect 3332 31780 3388 31836
rect 22876 31780 22932 31836
rect 3332 31724 6188 31780
rect 6244 31724 6254 31780
rect 7746 31724 7756 31780
rect 7812 31724 8204 31780
rect 8260 31724 10220 31780
rect 10276 31724 10780 31780
rect 10836 31724 10846 31780
rect 11666 31724 11676 31780
rect 11732 31724 12908 31780
rect 12964 31724 12974 31780
rect 14690 31724 14700 31780
rect 14756 31724 15036 31780
rect 15092 31724 15260 31780
rect 15316 31724 15326 31780
rect 17042 31724 17052 31780
rect 17108 31724 17276 31780
rect 17332 31724 17342 31780
rect 18722 31724 18732 31780
rect 18788 31724 21980 31780
rect 22036 31724 22046 31780
rect 22876 31724 23996 31780
rect 24052 31724 24062 31780
rect 25890 31724 25900 31780
rect 25956 31724 25966 31780
rect 26114 31724 26124 31780
rect 26180 31724 26572 31780
rect 26628 31724 26638 31780
rect 31826 31724 31836 31780
rect 31892 31724 34412 31780
rect 34468 31724 34478 31780
rect 42242 31724 42252 31780
rect 42308 31724 42588 31780
rect 42644 31724 42654 31780
rect 43586 31724 43596 31780
rect 43652 31724 46060 31780
rect 46116 31724 46126 31780
rect 47170 31724 47180 31780
rect 47236 31724 48412 31780
rect 48468 31724 48478 31780
rect 25900 31668 25956 31724
rect 2818 31612 2828 31668
rect 2884 31612 7980 31668
rect 8036 31612 8046 31668
rect 8614 31612 8652 31668
rect 8708 31612 8718 31668
rect 9650 31612 9660 31668
rect 9716 31612 13132 31668
rect 13188 31612 14588 31668
rect 14644 31612 18172 31668
rect 18228 31612 20412 31668
rect 20468 31612 20478 31668
rect 21980 31612 23772 31668
rect 23828 31612 23838 31668
rect 25106 31612 25116 31668
rect 25172 31612 25956 31668
rect 30818 31612 30828 31668
rect 30884 31612 31724 31668
rect 31780 31612 31790 31668
rect 34962 31612 34972 31668
rect 35028 31612 35868 31668
rect 35924 31612 35934 31668
rect 36838 31612 36876 31668
rect 36932 31612 36942 31668
rect 37314 31612 37324 31668
rect 37380 31612 37772 31668
rect 37828 31612 37838 31668
rect 38742 31612 38780 31668
rect 38836 31612 38846 31668
rect 41682 31612 41692 31668
rect 41748 31612 44268 31668
rect 44324 31612 44334 31668
rect 44706 31612 44716 31668
rect 44772 31612 45836 31668
rect 45892 31612 45902 31668
rect 49074 31612 49084 31668
rect 49140 31612 49756 31668
rect 49812 31612 49822 31668
rect 52658 31612 52668 31668
rect 52724 31612 54012 31668
rect 54068 31612 54078 31668
rect 21980 31556 22036 31612
rect 2034 31500 2044 31556
rect 2100 31500 6300 31556
rect 6356 31500 6366 31556
rect 7634 31500 7644 31556
rect 7700 31500 10556 31556
rect 10612 31500 10622 31556
rect 12002 31500 12012 31556
rect 12068 31500 12572 31556
rect 12628 31500 14980 31556
rect 15138 31500 15148 31556
rect 15204 31500 15596 31556
rect 15652 31500 15662 31556
rect 17378 31500 17388 31556
rect 17444 31500 19404 31556
rect 19460 31500 19470 31556
rect 19618 31500 19628 31556
rect 19684 31500 22036 31556
rect 22194 31500 22204 31556
rect 22260 31500 25900 31556
rect 25956 31500 26684 31556
rect 26740 31500 26750 31556
rect 28326 31500 28364 31556
rect 28420 31500 30492 31556
rect 30548 31500 30558 31556
rect 31154 31500 31164 31556
rect 31220 31500 31948 31556
rect 32004 31500 33516 31556
rect 33572 31500 33582 31556
rect 36530 31500 36540 31556
rect 36596 31500 37436 31556
rect 37492 31500 37502 31556
rect 45938 31500 45948 31556
rect 46004 31500 55244 31556
rect 55300 31500 55310 31556
rect 7644 31444 7700 31500
rect 14924 31444 14980 31500
rect 6178 31388 6188 31444
rect 6244 31388 7700 31444
rect 10434 31388 10444 31444
rect 10500 31388 12236 31444
rect 12292 31388 12302 31444
rect 14924 31388 15484 31444
rect 15540 31388 18060 31444
rect 18116 31388 18126 31444
rect 28018 31388 28028 31444
rect 28084 31388 36092 31444
rect 36148 31388 37660 31444
rect 37716 31388 38332 31444
rect 38388 31388 38398 31444
rect 39106 31388 39116 31444
rect 39172 31388 39452 31444
rect 39508 31388 39788 31444
rect 39844 31388 39854 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 3378 31276 3388 31332
rect 3444 31276 4172 31332
rect 4228 31276 6300 31332
rect 6356 31276 6636 31332
rect 6692 31276 8092 31332
rect 8148 31276 9660 31332
rect 9716 31276 9726 31332
rect 12114 31276 12124 31332
rect 12180 31276 12460 31332
rect 12516 31276 17276 31332
rect 17332 31276 17342 31332
rect 22754 31276 22764 31332
rect 22820 31276 22830 31332
rect 26226 31276 26236 31332
rect 26292 31276 38220 31332
rect 38276 31276 40572 31332
rect 40628 31276 40638 31332
rect 8530 31164 8540 31220
rect 8596 31164 10444 31220
rect 10500 31164 11228 31220
rect 11284 31164 11294 31220
rect 17378 31164 17388 31220
rect 17444 31164 17836 31220
rect 17892 31164 19068 31220
rect 19124 31164 19516 31220
rect 19572 31164 19582 31220
rect 21606 31164 21644 31220
rect 21700 31164 21710 31220
rect 8988 31052 9996 31108
rect 10052 31052 10062 31108
rect 16482 31052 16492 31108
rect 16548 31052 16716 31108
rect 16772 31052 21868 31108
rect 21924 31052 21934 31108
rect 8988 30996 9044 31052
rect 4162 30940 4172 30996
rect 4228 30940 5180 30996
rect 5236 30940 5246 30996
rect 5394 30940 5404 30996
rect 5460 30940 7084 30996
rect 7140 30940 7150 30996
rect 8418 30940 8428 30996
rect 8484 30940 8988 30996
rect 9044 30940 9054 30996
rect 9314 30940 9324 30996
rect 9380 30940 10108 30996
rect 10164 30940 10174 30996
rect 10322 30940 10332 30996
rect 10388 30940 10556 30996
rect 10612 30940 11900 30996
rect 11956 30940 11966 30996
rect 15138 30940 15148 30996
rect 15204 30940 15242 30996
rect 16146 30940 16156 30996
rect 16212 30940 16828 30996
rect 16884 30940 16894 30996
rect 19394 30940 19404 30996
rect 19460 30940 21308 30996
rect 21364 30940 22092 30996
rect 22148 30940 22158 30996
rect 22764 30884 22820 31276
rect 23986 31164 23996 31220
rect 24052 31164 26124 31220
rect 26180 31164 26190 31220
rect 28802 31164 28812 31220
rect 28868 31164 29372 31220
rect 29428 31164 32284 31220
rect 32340 31164 32620 31220
rect 32676 31164 33404 31220
rect 33460 31164 33470 31220
rect 33730 31164 33740 31220
rect 33796 31164 38108 31220
rect 38164 31164 38174 31220
rect 42690 31164 42700 31220
rect 42756 31164 43820 31220
rect 43876 31164 43886 31220
rect 47730 31164 47740 31220
rect 47796 31164 48188 31220
rect 48244 31164 48254 31220
rect 48402 31164 48412 31220
rect 48468 31164 50428 31220
rect 52770 31164 52780 31220
rect 52836 31164 53340 31220
rect 53396 31164 53406 31220
rect 50372 31108 50428 31164
rect 25666 31052 25676 31108
rect 25732 31052 26460 31108
rect 26516 31052 26526 31108
rect 30146 31052 30156 31108
rect 30212 31052 32732 31108
rect 32788 31052 34076 31108
rect 34132 31052 34142 31108
rect 34300 31052 36428 31108
rect 36484 31052 36876 31108
rect 36932 31052 36942 31108
rect 39106 31052 39116 31108
rect 39172 31052 42588 31108
rect 42644 31052 42654 31108
rect 47394 31052 47404 31108
rect 47460 31052 49756 31108
rect 49812 31052 49980 31108
rect 50036 31052 50046 31108
rect 50372 31052 51380 31108
rect 51538 31052 51548 31108
rect 51604 31052 52444 31108
rect 52500 31052 52510 31108
rect 34300 30996 34356 31052
rect 51324 30996 51380 31052
rect 24994 30940 25004 30996
rect 25060 30940 25564 30996
rect 25620 30940 25630 30996
rect 27346 30940 27356 30996
rect 27412 30940 27804 30996
rect 27860 30940 28476 30996
rect 28532 30940 28542 30996
rect 30930 30940 30940 30996
rect 30996 30940 31836 30996
rect 31892 30940 32844 30996
rect 32900 30940 34356 30996
rect 35858 30940 35868 30996
rect 35924 30940 36764 30996
rect 36820 30940 36830 30996
rect 51324 30940 52668 30996
rect 52724 30940 52734 30996
rect 3826 30828 3836 30884
rect 3892 30828 3948 30884
rect 4004 30828 4844 30884
rect 4900 30828 6748 30884
rect 6804 30828 6814 30884
rect 7298 30828 7308 30884
rect 7364 30828 11228 30884
rect 11284 30828 14812 30884
rect 14868 30828 16044 30884
rect 16100 30828 16110 30884
rect 21746 30828 21756 30884
rect 21812 30828 22652 30884
rect 22708 30828 24444 30884
rect 24500 30828 25116 30884
rect 25172 30828 25676 30884
rect 25732 30828 25742 30884
rect 34290 30828 34300 30884
rect 34356 30828 36652 30884
rect 36708 30828 36718 30884
rect 39218 30828 39228 30884
rect 39284 30828 40012 30884
rect 40068 30828 40078 30884
rect 40786 30828 40796 30884
rect 40852 30828 42140 30884
rect 42196 30828 42812 30884
rect 42868 30828 42878 30884
rect 43698 30828 43708 30884
rect 43764 30828 51772 30884
rect 51828 30828 52556 30884
rect 52612 30828 53116 30884
rect 53172 30828 53182 30884
rect 1474 30716 1484 30772
rect 1540 30716 4620 30772
rect 4676 30716 4686 30772
rect 13682 30716 13692 30772
rect 13748 30716 20300 30772
rect 20356 30716 20366 30772
rect 26562 30716 26572 30772
rect 26628 30716 27580 30772
rect 27636 30716 27646 30772
rect 29922 30716 29932 30772
rect 29988 30716 31052 30772
rect 31108 30716 31118 30772
rect 32722 30716 32732 30772
rect 32788 30716 35644 30772
rect 35700 30716 36204 30772
rect 36260 30716 36270 30772
rect 46386 30716 46396 30772
rect 46452 30716 56588 30772
rect 56644 30716 56812 30772
rect 56868 30716 57372 30772
rect 57428 30716 57708 30772
rect 57764 30716 57774 30772
rect 10994 30604 11004 30660
rect 11060 30604 11116 30660
rect 11172 30604 11182 30660
rect 19282 30604 19292 30660
rect 19348 30604 19628 30660
rect 19684 30604 19694 30660
rect 23650 30604 23660 30660
rect 23716 30604 25564 30660
rect 25620 30604 25900 30660
rect 25956 30604 25966 30660
rect 38742 30604 38780 30660
rect 38836 30604 38846 30660
rect 45378 30604 45388 30660
rect 45444 30604 46620 30660
rect 46676 30604 46686 30660
rect 48178 30604 48188 30660
rect 48244 30604 51324 30660
rect 51380 30604 51390 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 6626 30492 6636 30548
rect 6692 30492 9772 30548
rect 9828 30492 11116 30548
rect 11172 30492 11788 30548
rect 11844 30492 11854 30548
rect 18386 30492 18396 30548
rect 18452 30492 19404 30548
rect 19460 30492 21644 30548
rect 21700 30492 21710 30548
rect 24546 30492 24556 30548
rect 24612 30492 30380 30548
rect 30436 30492 30446 30548
rect 32946 30492 32956 30548
rect 33012 30492 33292 30548
rect 33348 30492 34972 30548
rect 35028 30492 35038 30548
rect 3378 30380 3388 30436
rect 3444 30380 5628 30436
rect 5684 30380 8428 30436
rect 8484 30380 8494 30436
rect 8866 30380 8876 30436
rect 8932 30380 16940 30436
rect 16996 30380 18172 30436
rect 18228 30380 18238 30436
rect 18992 30380 19068 30436
rect 19124 30380 19628 30436
rect 19684 30380 19694 30436
rect 24434 30380 24444 30436
rect 24500 30380 24780 30436
rect 24836 30380 24846 30436
rect 34738 30380 34748 30436
rect 34804 30380 35532 30436
rect 35588 30380 35598 30436
rect 5058 30268 5068 30324
rect 5124 30268 5404 30324
rect 5460 30268 5470 30324
rect 11106 30268 11116 30324
rect 11172 30268 11676 30324
rect 11732 30268 11742 30324
rect 11890 30268 11900 30324
rect 11956 30268 13132 30324
rect 13188 30268 14140 30324
rect 14196 30268 14206 30324
rect 15698 30268 15708 30324
rect 15764 30268 16604 30324
rect 16660 30268 16670 30324
rect 18722 30268 18732 30324
rect 18788 30268 19180 30324
rect 19236 30268 19246 30324
rect 20850 30268 20860 30324
rect 20916 30268 25676 30324
rect 25732 30268 26012 30324
rect 26068 30268 26078 30324
rect 38322 30268 38332 30324
rect 38388 30268 40348 30324
rect 40404 30268 40414 30324
rect 48402 30268 48412 30324
rect 48468 30268 49868 30324
rect 49924 30268 49934 30324
rect 2706 30156 2716 30212
rect 2772 30156 3276 30212
rect 3332 30156 3342 30212
rect 7186 30156 7196 30212
rect 7252 30156 7756 30212
rect 7812 30156 7822 30212
rect 7970 30156 7980 30212
rect 8036 30156 8876 30212
rect 8932 30156 8942 30212
rect 10658 30156 10668 30212
rect 10724 30156 11004 30212
rect 11060 30156 11070 30212
rect 11330 30156 11340 30212
rect 11396 30156 16380 30212
rect 16436 30156 16446 30212
rect 17266 30156 17276 30212
rect 17332 30156 22652 30212
rect 22708 30156 22718 30212
rect 23202 30156 23212 30212
rect 23268 30156 25340 30212
rect 25396 30156 25676 30212
rect 25732 30156 27132 30212
rect 27188 30156 27198 30212
rect 29250 30156 29260 30212
rect 29316 30156 30828 30212
rect 30884 30156 30894 30212
rect 31938 30156 31948 30212
rect 32004 30156 33628 30212
rect 33684 30156 34300 30212
rect 34356 30156 34366 30212
rect 36082 30156 36092 30212
rect 36148 30156 41804 30212
rect 41860 30156 42924 30212
rect 42980 30156 42990 30212
rect 47506 30156 47516 30212
rect 47572 30156 48524 30212
rect 48580 30156 49084 30212
rect 49140 30156 49150 30212
rect 52658 30156 52668 30212
rect 52724 30156 53676 30212
rect 53732 30156 53742 30212
rect 54898 30156 54908 30212
rect 54964 30156 55468 30212
rect 55524 30156 55534 30212
rect 9202 30044 9212 30100
rect 9268 30044 12348 30100
rect 12404 30044 12908 30100
rect 12964 30044 12974 30100
rect 19282 30044 19292 30100
rect 19348 30044 19740 30100
rect 19796 30044 19806 30100
rect 21970 30044 21980 30100
rect 22036 30044 22316 30100
rect 22372 30044 22988 30100
rect 23044 30044 23436 30100
rect 23492 30044 23502 30100
rect 24210 30044 24220 30100
rect 24276 30044 25396 30100
rect 34514 30044 34524 30100
rect 34580 30044 36988 30100
rect 37044 30044 37054 30100
rect 40002 30044 40012 30100
rect 40068 30044 40572 30100
rect 40628 30044 42028 30100
rect 42084 30044 43484 30100
rect 43540 30044 43550 30100
rect 45602 30044 45612 30100
rect 45668 30044 49196 30100
rect 49252 30044 50092 30100
rect 50148 30044 50158 30100
rect 50754 30044 50764 30100
rect 50820 30044 52108 30100
rect 52164 30044 52174 30100
rect 25340 29988 25396 30044
rect 10368 29932 10444 29988
rect 10500 29932 11228 29988
rect 11284 29932 11294 29988
rect 11788 29932 13580 29988
rect 13636 29932 14028 29988
rect 14084 29932 14094 29988
rect 19842 29932 19852 29988
rect 19908 29932 20244 29988
rect 20402 29932 20412 29988
rect 20468 29932 21532 29988
rect 21588 29932 25116 29988
rect 25172 29932 25182 29988
rect 25340 29932 28924 29988
rect 28980 29932 28990 29988
rect 29586 29932 29596 29988
rect 29652 29932 33852 29988
rect 33908 29932 34636 29988
rect 34692 29932 34702 29988
rect 38882 29932 38892 29988
rect 38948 29932 41692 29988
rect 41748 29932 41758 29988
rect 46050 29932 46060 29988
rect 46116 29932 47292 29988
rect 47348 29932 47740 29988
rect 47796 29932 48300 29988
rect 48356 29932 48366 29988
rect 11788 29876 11844 29932
rect 20188 29876 20244 29932
rect 27580 29876 27636 29932
rect 1922 29820 1932 29876
rect 1988 29820 2380 29876
rect 2436 29820 4620 29876
rect 4676 29820 4686 29876
rect 6402 29820 6412 29876
rect 6468 29820 11844 29876
rect 12786 29820 12796 29876
rect 12852 29820 15036 29876
rect 15092 29820 17164 29876
rect 17220 29820 17724 29876
rect 17780 29820 17790 29876
rect 20188 29820 22428 29876
rect 22484 29820 22494 29876
rect 26114 29820 26124 29876
rect 26180 29820 26796 29876
rect 26852 29820 26862 29876
rect 27570 29820 27580 29876
rect 27636 29820 27646 29876
rect 33852 29820 35420 29876
rect 35476 29820 35980 29876
rect 36036 29820 36046 29876
rect 46274 29820 46284 29876
rect 46340 29820 46956 29876
rect 47012 29820 47022 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 33852 29764 33908 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 4284 29708 11676 29764
rect 11732 29708 11742 29764
rect 12226 29708 12236 29764
rect 12292 29708 14252 29764
rect 14308 29708 14318 29764
rect 18162 29708 18172 29764
rect 18228 29708 19292 29764
rect 19348 29708 19358 29764
rect 22082 29708 22092 29764
rect 22148 29708 25956 29764
rect 33058 29708 33068 29764
rect 33124 29708 33404 29764
rect 33460 29708 33852 29764
rect 33908 29708 33918 29764
rect 35074 29708 35084 29764
rect 35140 29708 37324 29764
rect 37380 29708 38892 29764
rect 38948 29708 38958 29764
rect 44146 29708 44156 29764
rect 44212 29708 45164 29764
rect 45220 29708 46396 29764
rect 46452 29708 46462 29764
rect 4284 29652 4340 29708
rect 25900 29652 25956 29708
rect 3462 29596 3500 29652
rect 3556 29596 3566 29652
rect 4050 29596 4060 29652
rect 4116 29596 4284 29652
rect 4340 29596 4350 29652
rect 5506 29596 5516 29652
rect 5572 29596 6076 29652
rect 6132 29596 6142 29652
rect 10434 29596 10444 29652
rect 10500 29596 11116 29652
rect 11172 29596 11182 29652
rect 11442 29596 11452 29652
rect 11508 29596 12684 29652
rect 12740 29596 14140 29652
rect 14196 29596 14206 29652
rect 16594 29596 16604 29652
rect 16660 29596 17500 29652
rect 17556 29596 18452 29652
rect 25638 29596 25676 29652
rect 25732 29596 25742 29652
rect 25890 29596 25900 29652
rect 25956 29596 26012 29652
rect 26068 29596 26078 29652
rect 29810 29596 29820 29652
rect 29876 29596 33404 29652
rect 33460 29596 33470 29652
rect 34962 29596 34972 29652
rect 35028 29596 37884 29652
rect 37940 29596 37950 29652
rect 46274 29596 46284 29652
rect 46340 29596 47516 29652
rect 47572 29596 48076 29652
rect 48132 29596 48142 29652
rect 18396 29540 18452 29596
rect 4610 29484 4620 29540
rect 4676 29484 4844 29540
rect 4900 29484 6860 29540
rect 6916 29484 6926 29540
rect 8306 29484 8316 29540
rect 8372 29484 10780 29540
rect 10836 29484 11004 29540
rect 11060 29484 11070 29540
rect 11666 29484 11676 29540
rect 11732 29484 12908 29540
rect 12964 29484 13244 29540
rect 13300 29484 13310 29540
rect 15260 29484 15820 29540
rect 15876 29484 17052 29540
rect 17108 29484 18172 29540
rect 18228 29484 18238 29540
rect 18396 29484 21980 29540
rect 22036 29484 22046 29540
rect 25106 29484 25116 29540
rect 25172 29484 27132 29540
rect 27188 29484 27198 29540
rect 29138 29484 29148 29540
rect 29204 29484 30156 29540
rect 30212 29484 30604 29540
rect 30660 29484 30670 29540
rect 33618 29484 33628 29540
rect 33684 29484 37436 29540
rect 37492 29484 37502 29540
rect 52994 29484 53004 29540
rect 53060 29484 54124 29540
rect 54180 29484 54190 29540
rect 56018 29484 56028 29540
rect 56084 29484 57484 29540
rect 57540 29484 57550 29540
rect 15260 29428 15316 29484
rect 34972 29428 35028 29484
rect 9846 29372 9884 29428
rect 9940 29372 13580 29428
rect 13636 29372 13804 29428
rect 13860 29372 13870 29428
rect 14354 29372 14364 29428
rect 14420 29372 14924 29428
rect 14980 29372 14990 29428
rect 15250 29372 15260 29428
rect 15316 29372 15326 29428
rect 16146 29372 16156 29428
rect 16212 29372 21140 29428
rect 26450 29372 26460 29428
rect 26516 29372 26908 29428
rect 26964 29372 26974 29428
rect 31378 29372 31388 29428
rect 31444 29372 31948 29428
rect 32004 29372 32014 29428
rect 34962 29372 34972 29428
rect 35028 29372 35038 29428
rect 35186 29372 35196 29428
rect 35252 29372 35756 29428
rect 35812 29372 35822 29428
rect 40450 29372 40460 29428
rect 40516 29372 41692 29428
rect 41748 29372 41758 29428
rect 55412 29372 55692 29428
rect 55748 29372 55758 29428
rect 21084 29316 21140 29372
rect 10994 29260 11004 29316
rect 11060 29260 11116 29316
rect 11172 29260 11182 29316
rect 13682 29260 13692 29316
rect 13748 29260 16996 29316
rect 19618 29260 19628 29316
rect 19684 29260 20300 29316
rect 20356 29260 20366 29316
rect 21046 29260 21084 29316
rect 21140 29260 21150 29316
rect 28018 29260 28028 29316
rect 28084 29260 28588 29316
rect 28644 29260 28654 29316
rect 29810 29260 29820 29316
rect 29876 29260 30044 29316
rect 30100 29260 30828 29316
rect 30884 29260 30894 29316
rect 34748 29260 38220 29316
rect 38276 29260 38286 29316
rect 44034 29260 44044 29316
rect 44100 29260 45724 29316
rect 45780 29260 46172 29316
rect 46228 29260 46238 29316
rect 54562 29260 54572 29316
rect 54628 29260 55356 29316
rect 55412 29260 55468 29372
rect 16940 29204 16996 29260
rect 5842 29148 5852 29204
rect 5908 29148 8540 29204
rect 8596 29148 9996 29204
rect 10052 29148 11228 29204
rect 11284 29148 11294 29204
rect 14354 29148 14364 29204
rect 14420 29148 14812 29204
rect 14868 29148 14878 29204
rect 16930 29148 16940 29204
rect 16996 29148 23548 29204
rect 23604 29148 23614 29204
rect 23762 29148 23772 29204
rect 23828 29148 25900 29204
rect 25956 29148 25966 29204
rect 26198 29148 26236 29204
rect 26292 29148 26302 29204
rect 30258 29148 30268 29204
rect 30324 29148 30604 29204
rect 30660 29148 30670 29204
rect 3910 29036 3948 29092
rect 4004 29036 4014 29092
rect 8306 29036 8316 29092
rect 8372 29036 14028 29092
rect 14084 29036 17612 29092
rect 17668 29036 17678 29092
rect 25228 29036 30044 29092
rect 30100 29036 30110 29092
rect 34486 29036 34524 29092
rect 34580 29036 34590 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 25228 28980 25284 29036
rect 34748 28980 34804 29260
rect 34962 29148 34972 29204
rect 35028 29148 35084 29204
rect 35140 29148 35150 29204
rect 35410 29148 35420 29204
rect 35476 29148 36092 29204
rect 36148 29148 36158 29204
rect 38322 29148 38332 29204
rect 38388 29148 41580 29204
rect 41636 29148 43148 29204
rect 43204 29148 43214 29204
rect 43362 29148 43372 29204
rect 43428 29148 46060 29204
rect 46116 29148 46126 29204
rect 55682 29148 55692 29204
rect 55748 29148 58044 29204
rect 58100 29148 58110 29204
rect 40562 29036 40572 29092
rect 40628 29036 54348 29092
rect 54404 29036 55132 29092
rect 55188 29036 56140 29092
rect 56196 29036 56206 29092
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 7532 28924 7868 28980
rect 7924 28924 9324 28980
rect 9380 28924 9390 28980
rect 13132 28924 15148 28980
rect 22754 28924 22764 28980
rect 22820 28924 25228 28980
rect 25284 28924 25294 28980
rect 25778 28924 25788 28980
rect 25844 28924 31388 28980
rect 31444 28924 31454 28980
rect 32274 28924 32284 28980
rect 32340 28924 32732 28980
rect 32788 28924 32798 28980
rect 33170 28924 33180 28980
rect 33236 28924 34748 28980
rect 34804 28924 34814 28980
rect 43922 28924 43932 28980
rect 43988 28924 56364 28980
rect 56420 28924 56700 28980
rect 56756 28924 57260 28980
rect 57316 28924 57326 28980
rect 57670 28924 57708 28980
rect 57764 28924 57774 28980
rect 7532 28868 7588 28924
rect 13132 28868 13188 28924
rect 3714 28812 3724 28868
rect 3780 28812 4172 28868
rect 4228 28812 7588 28868
rect 7746 28812 7756 28868
rect 7812 28812 13132 28868
rect 13188 28812 13198 28868
rect 15092 28756 15148 28924
rect 17490 28812 17500 28868
rect 17556 28812 17612 28868
rect 17668 28812 17678 28868
rect 18274 28812 18284 28868
rect 18340 28812 18508 28868
rect 18564 28812 18844 28868
rect 18900 28812 18910 28868
rect 24546 28812 24556 28868
rect 24612 28812 39788 28868
rect 39844 28812 39854 28868
rect 40002 28812 40012 28868
rect 40068 28812 40684 28868
rect 40740 28812 41916 28868
rect 41972 28812 41982 28868
rect 52658 28812 52668 28868
rect 52724 28812 53452 28868
rect 53508 28812 53518 28868
rect 3490 28700 3500 28756
rect 3556 28700 4508 28756
rect 4564 28700 5180 28756
rect 5236 28700 5246 28756
rect 6374 28700 6412 28756
rect 6468 28700 6478 28756
rect 11778 28700 11788 28756
rect 11844 28700 12796 28756
rect 12852 28700 12862 28756
rect 13010 28700 13020 28756
rect 13076 28700 14420 28756
rect 14578 28700 14588 28756
rect 14644 28700 14924 28756
rect 14980 28700 14990 28756
rect 15092 28700 17836 28756
rect 17892 28700 17902 28756
rect 22418 28700 22428 28756
rect 22484 28700 28028 28756
rect 28084 28700 28094 28756
rect 33842 28700 33852 28756
rect 33908 28700 34524 28756
rect 34580 28700 35868 28756
rect 35924 28700 37324 28756
rect 37380 28700 40796 28756
rect 40852 28700 40862 28756
rect 45378 28700 45388 28756
rect 45444 28700 45948 28756
rect 46004 28700 46014 28756
rect 46274 28700 46284 28756
rect 46340 28700 47068 28756
rect 47124 28700 47134 28756
rect 53554 28700 53564 28756
rect 53620 28700 58716 28756
rect 58772 28700 58782 28756
rect 14364 28644 14420 28700
rect 12562 28588 12572 28644
rect 12628 28588 14140 28644
rect 14196 28588 14206 28644
rect 14364 28588 15036 28644
rect 15092 28588 16940 28644
rect 16996 28588 17724 28644
rect 17780 28588 17790 28644
rect 18162 28588 18172 28644
rect 18228 28588 18620 28644
rect 18676 28588 19348 28644
rect 20514 28588 20524 28644
rect 20580 28588 25676 28644
rect 25732 28588 25742 28644
rect 26114 28588 26124 28644
rect 26180 28588 27132 28644
rect 27188 28588 27198 28644
rect 27766 28588 27804 28644
rect 27860 28588 28476 28644
rect 28532 28588 28542 28644
rect 30818 28588 30828 28644
rect 30884 28588 32284 28644
rect 32340 28588 32956 28644
rect 33012 28588 33022 28644
rect 34514 28588 34524 28644
rect 34580 28588 35756 28644
rect 35812 28588 35822 28644
rect 35970 28588 35980 28644
rect 36036 28588 38220 28644
rect 38276 28588 38286 28644
rect 42354 28588 42364 28644
rect 42420 28588 42924 28644
rect 42980 28588 44716 28644
rect 44772 28588 44782 28644
rect 46610 28588 46620 28644
rect 46676 28588 47180 28644
rect 47236 28588 47246 28644
rect 50418 28588 50428 28644
rect 50484 28588 50876 28644
rect 50932 28588 52108 28644
rect 52164 28588 52174 28644
rect 55346 28588 55356 28644
rect 55412 28588 56364 28644
rect 56420 28588 56430 28644
rect 19292 28532 19348 28588
rect 5394 28476 5404 28532
rect 5460 28476 5740 28532
rect 5796 28476 7084 28532
rect 7140 28476 7150 28532
rect 7970 28476 7980 28532
rect 8036 28476 8988 28532
rect 9044 28476 9054 28532
rect 9650 28476 9660 28532
rect 9716 28476 10668 28532
rect 10724 28476 12348 28532
rect 12404 28476 12414 28532
rect 13654 28476 13692 28532
rect 13748 28476 13758 28532
rect 14914 28476 14924 28532
rect 14980 28476 18844 28532
rect 18900 28476 19068 28532
rect 19124 28476 19134 28532
rect 19292 28476 20300 28532
rect 20356 28476 22204 28532
rect 22260 28476 23772 28532
rect 23828 28476 24220 28532
rect 24276 28476 24286 28532
rect 26852 28476 27020 28532
rect 27076 28476 27692 28532
rect 27748 28476 28140 28532
rect 28196 28476 28206 28532
rect 28578 28476 28588 28532
rect 28644 28476 29932 28532
rect 29988 28476 30492 28532
rect 30548 28476 30558 28532
rect 32610 28476 32620 28532
rect 32676 28476 32844 28532
rect 32900 28476 32910 28532
rect 34626 28476 34636 28532
rect 34692 28476 35084 28532
rect 35140 28476 35150 28532
rect 36082 28476 36092 28532
rect 36148 28476 38108 28532
rect 38164 28476 38174 28532
rect 39666 28476 39676 28532
rect 39732 28476 40908 28532
rect 40964 28476 40974 28532
rect 41906 28476 41916 28532
rect 41972 28476 43708 28532
rect 43764 28476 43774 28532
rect 55010 28476 55020 28532
rect 55076 28476 57708 28532
rect 57764 28476 57774 28532
rect 26852 28420 26908 28476
rect 9090 28364 9100 28420
rect 9156 28364 10780 28420
rect 10836 28364 10846 28420
rect 13794 28364 13804 28420
rect 13860 28364 16436 28420
rect 16594 28364 16604 28420
rect 16660 28364 20412 28420
rect 20468 28364 20478 28420
rect 20962 28364 20972 28420
rect 21028 28364 23660 28420
rect 23716 28364 24108 28420
rect 24164 28364 26908 28420
rect 30146 28364 30156 28420
rect 30212 28364 30940 28420
rect 30996 28364 31006 28420
rect 32498 28364 32508 28420
rect 32564 28364 37548 28420
rect 37604 28364 37614 28420
rect 38612 28364 38780 28420
rect 38836 28364 38846 28420
rect 42578 28364 42588 28420
rect 42644 28364 44044 28420
rect 44100 28364 44110 28420
rect 16380 28308 16436 28364
rect 20412 28308 20468 28364
rect 30492 28308 30548 28364
rect 38612 28308 38668 28364
rect 8082 28252 8092 28308
rect 8148 28252 10444 28308
rect 10500 28252 10510 28308
rect 14242 28252 14252 28308
rect 14308 28252 16156 28308
rect 16212 28252 16222 28308
rect 16380 28252 18732 28308
rect 18788 28252 18798 28308
rect 20412 28252 21196 28308
rect 21252 28252 21262 28308
rect 24994 28252 25004 28308
rect 25060 28252 30492 28308
rect 30548 28252 30558 28308
rect 33068 28252 34188 28308
rect 34244 28252 38668 28308
rect 41122 28252 41132 28308
rect 41188 28252 41692 28308
rect 41748 28252 43036 28308
rect 43092 28252 43102 28308
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 33068 28196 33124 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 10098 28140 10108 28196
rect 10164 28140 13244 28196
rect 13300 28140 13692 28196
rect 13748 28140 18396 28196
rect 18452 28140 18462 28196
rect 33058 28140 33068 28196
rect 33124 28140 33134 28196
rect 39890 28140 39900 28196
rect 39956 28140 40236 28196
rect 40292 28140 44604 28196
rect 44660 28140 44670 28196
rect 45826 28140 45836 28196
rect 45892 28140 46508 28196
rect 46564 28140 46574 28196
rect 15698 28028 15708 28084
rect 15764 28028 15932 28084
rect 15988 28028 16380 28084
rect 16436 28028 18620 28084
rect 18676 28028 18686 28084
rect 28354 28028 28364 28084
rect 28420 28028 29372 28084
rect 29428 28028 31388 28084
rect 31444 28028 32396 28084
rect 32452 28028 33180 28084
rect 33236 28028 33246 28084
rect 33842 28028 33852 28084
rect 33908 28028 34188 28084
rect 34244 28028 34254 28084
rect 36306 28028 36316 28084
rect 36372 28028 36764 28084
rect 36820 28028 36830 28084
rect 42354 28028 42364 28084
rect 42420 28028 43596 28084
rect 43652 28028 43662 28084
rect 2034 27916 2044 27972
rect 2100 27916 3388 27972
rect 6514 27916 6524 27972
rect 6580 27916 7532 27972
rect 7588 27916 8988 27972
rect 9044 27916 9772 27972
rect 9828 27916 9838 27972
rect 9986 27916 9996 27972
rect 10052 27916 10108 27972
rect 10164 27916 11004 27972
rect 11060 27916 11070 27972
rect 15138 27916 15148 27972
rect 15204 27916 15214 27972
rect 16146 27916 16156 27972
rect 16212 27916 16492 27972
rect 16548 27916 16558 27972
rect 25442 27916 25452 27972
rect 25508 27916 25900 27972
rect 25956 27916 25966 27972
rect 27010 27916 27020 27972
rect 27076 27916 27580 27972
rect 27636 27916 28476 27972
rect 28532 27916 28542 27972
rect 36530 27916 36540 27972
rect 36596 27916 36652 27972
rect 36708 27916 36718 27972
rect 45602 27916 45612 27972
rect 45668 27916 46732 27972
rect 46788 27916 47404 27972
rect 47460 27916 47964 27972
rect 48020 27916 48636 27972
rect 48692 27916 48702 27972
rect 3332 27860 3388 27916
rect 15148 27860 15204 27916
rect 3332 27804 8092 27860
rect 8148 27804 8158 27860
rect 8418 27804 8428 27860
rect 8484 27804 8876 27860
rect 8932 27804 9996 27860
rect 10052 27804 10062 27860
rect 15092 27804 16716 27860
rect 16772 27804 16782 27860
rect 19282 27804 19292 27860
rect 19348 27804 19852 27860
rect 19908 27804 19918 27860
rect 22754 27804 22764 27860
rect 22820 27804 24556 27860
rect 24612 27804 27804 27860
rect 27860 27804 27870 27860
rect 28018 27804 28028 27860
rect 28084 27804 28700 27860
rect 28756 27804 28766 27860
rect 30604 27804 36988 27860
rect 37044 27804 38556 27860
rect 38612 27804 45500 27860
rect 45556 27804 45566 27860
rect 45938 27804 45948 27860
rect 46004 27804 47740 27860
rect 47796 27804 48972 27860
rect 49028 27804 49038 27860
rect 50642 27804 50652 27860
rect 50708 27804 51100 27860
rect 51156 27804 51166 27860
rect 15092 27748 15148 27804
rect 30604 27748 30660 27804
rect 1922 27692 1932 27748
rect 1988 27692 3500 27748
rect 3556 27692 3836 27748
rect 3892 27692 3902 27748
rect 8978 27692 8988 27748
rect 9044 27692 15148 27748
rect 15362 27692 15372 27748
rect 15428 27692 16268 27748
rect 16324 27692 16334 27748
rect 30258 27692 30268 27748
rect 30324 27692 30604 27748
rect 30660 27692 30670 27748
rect 34738 27692 34748 27748
rect 34804 27692 41244 27748
rect 41300 27692 41310 27748
rect 49634 27692 49644 27748
rect 49700 27692 50092 27748
rect 50148 27692 50158 27748
rect 51100 27692 51772 27748
rect 51828 27692 52444 27748
rect 52500 27692 52510 27748
rect 51100 27636 51156 27692
rect 4162 27580 4172 27636
rect 4228 27580 6972 27636
rect 7028 27580 7038 27636
rect 10322 27580 10332 27636
rect 10388 27580 13356 27636
rect 13412 27580 14588 27636
rect 14644 27580 15596 27636
rect 15652 27580 15662 27636
rect 19954 27580 19964 27636
rect 20020 27580 37100 27636
rect 37156 27580 38668 27636
rect 38724 27580 38734 27636
rect 40002 27580 40012 27636
rect 40068 27580 41020 27636
rect 41076 27580 41086 27636
rect 41346 27580 41356 27636
rect 41412 27580 42924 27636
rect 42980 27580 43596 27636
rect 43652 27580 43662 27636
rect 51090 27580 51100 27636
rect 51156 27580 51166 27636
rect 7970 27468 7980 27524
rect 8036 27468 8316 27524
rect 8372 27468 8382 27524
rect 24546 27468 24556 27524
rect 24612 27468 28588 27524
rect 28644 27468 32508 27524
rect 32564 27468 32574 27524
rect 35634 27468 35644 27524
rect 35700 27468 36876 27524
rect 36932 27468 36942 27524
rect 37650 27468 37660 27524
rect 37716 27468 41468 27524
rect 41524 27468 41804 27524
rect 41860 27468 41870 27524
rect 51202 27468 51212 27524
rect 51268 27468 51772 27524
rect 51828 27468 51838 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 18050 27356 18060 27412
rect 18116 27356 26236 27412
rect 26292 27356 28028 27412
rect 28084 27356 28094 27412
rect 31826 27356 31836 27412
rect 31892 27356 33852 27412
rect 33908 27356 33918 27412
rect 36530 27356 36540 27412
rect 36596 27356 40236 27412
rect 40292 27356 40302 27412
rect 41346 27356 41356 27412
rect 41412 27356 41422 27412
rect 46050 27356 46060 27412
rect 46116 27356 47404 27412
rect 47460 27356 47470 27412
rect 41356 27300 41412 27356
rect 3332 27244 5292 27300
rect 5348 27244 5358 27300
rect 8642 27244 8652 27300
rect 8708 27244 12460 27300
rect 12516 27244 12526 27300
rect 26338 27244 26348 27300
rect 26404 27244 29484 27300
rect 29540 27244 30716 27300
rect 30772 27244 31164 27300
rect 31220 27244 32844 27300
rect 32900 27244 32910 27300
rect 35298 27244 35308 27300
rect 35364 27244 39116 27300
rect 39172 27244 39182 27300
rect 39442 27244 39452 27300
rect 39508 27244 41412 27300
rect 45602 27244 45612 27300
rect 45668 27244 46956 27300
rect 47012 27244 47022 27300
rect 48402 27244 48412 27300
rect 48468 27244 50652 27300
rect 50708 27244 50718 27300
rect 3332 27188 3388 27244
rect 2594 27132 2604 27188
rect 2660 27132 3388 27188
rect 3490 27132 3500 27188
rect 3556 27132 4172 27188
rect 4228 27132 4238 27188
rect 4946 27132 4956 27188
rect 5012 27132 6300 27188
rect 6356 27132 8316 27188
rect 8372 27132 8382 27188
rect 8754 27132 8764 27188
rect 8820 27132 10332 27188
rect 10388 27132 10398 27188
rect 12114 27132 12124 27188
rect 12180 27132 14700 27188
rect 14756 27132 14766 27188
rect 20850 27132 20860 27188
rect 20916 27132 26572 27188
rect 26628 27132 28028 27188
rect 28084 27132 28094 27188
rect 30370 27132 30380 27188
rect 30436 27132 30828 27188
rect 30884 27132 34748 27188
rect 34804 27132 34814 27188
rect 36838 27132 36876 27188
rect 36932 27132 36942 27188
rect 38658 27132 38668 27188
rect 38724 27132 39228 27188
rect 39284 27132 41356 27188
rect 41412 27132 41422 27188
rect 42690 27132 42700 27188
rect 42756 27132 44492 27188
rect 44548 27132 44558 27188
rect 46162 27132 46172 27188
rect 46228 27132 49532 27188
rect 49588 27132 49598 27188
rect 49746 27132 49756 27188
rect 49812 27132 50428 27188
rect 50484 27132 50494 27188
rect 51202 27132 51212 27188
rect 51268 27132 55020 27188
rect 55076 27132 55086 27188
rect 3042 27020 3052 27076
rect 3108 27020 6748 27076
rect 6804 27020 7084 27076
rect 7140 27020 7150 27076
rect 8082 27020 8092 27076
rect 8148 27020 9996 27076
rect 10052 27020 10062 27076
rect 12002 27020 12012 27076
rect 12068 27020 12078 27076
rect 15362 27020 15372 27076
rect 15428 27020 23996 27076
rect 24052 27020 25004 27076
rect 25060 27020 26012 27076
rect 26068 27020 26078 27076
rect 28690 27020 28700 27076
rect 28756 27020 30940 27076
rect 30996 27020 31612 27076
rect 31668 27020 31678 27076
rect 32498 27020 32508 27076
rect 32564 27020 32844 27076
rect 32900 27020 32910 27076
rect 33814 27020 33852 27076
rect 33908 27020 33918 27076
rect 39554 27020 39564 27076
rect 39620 27020 40572 27076
rect 40628 27020 40638 27076
rect 41906 27020 41916 27076
rect 41972 27020 52108 27076
rect 52164 27020 52780 27076
rect 52836 27020 53676 27076
rect 53732 27020 53742 27076
rect 12012 26964 12068 27020
rect 2482 26908 2492 26964
rect 2548 26908 4732 26964
rect 4788 26908 4798 26964
rect 4946 26908 4956 26964
rect 5012 26908 5292 26964
rect 5348 26908 6524 26964
rect 6580 26908 6590 26964
rect 10546 26908 10556 26964
rect 10612 26908 10892 26964
rect 10948 26908 11452 26964
rect 11508 26908 12068 26964
rect 15810 26908 15820 26964
rect 15876 26908 16940 26964
rect 16996 26908 18172 26964
rect 18228 26908 18238 26964
rect 19170 26908 19180 26964
rect 19236 26908 20860 26964
rect 20916 26908 20926 26964
rect 27234 26908 27244 26964
rect 27300 26908 28812 26964
rect 28868 26908 28878 26964
rect 34402 26908 34412 26964
rect 34468 26908 34972 26964
rect 35028 26908 35038 26964
rect 39330 26908 39340 26964
rect 39396 26908 40908 26964
rect 40964 26908 42252 26964
rect 42308 26908 43148 26964
rect 43204 26908 43214 26964
rect 43652 26908 44044 26964
rect 44100 26908 44268 26964
rect 44324 26908 44334 26964
rect 46498 26908 46508 26964
rect 46564 26908 47516 26964
rect 47572 26908 48188 26964
rect 48244 26908 48254 26964
rect 50530 26908 50540 26964
rect 50596 26908 51324 26964
rect 51380 26908 51996 26964
rect 52052 26908 52668 26964
rect 52724 26908 52734 26964
rect 43652 26852 43708 26908
rect 1922 26796 1932 26852
rect 1988 26796 2380 26852
rect 2436 26796 2446 26852
rect 5058 26796 5068 26852
rect 5124 26796 8540 26852
rect 8596 26796 9436 26852
rect 9492 26796 11228 26852
rect 11284 26796 11676 26852
rect 11732 26796 11742 26852
rect 12450 26796 12460 26852
rect 12516 26796 12796 26852
rect 12852 26796 12862 26852
rect 13010 26796 13020 26852
rect 13076 26796 15708 26852
rect 15764 26796 15774 26852
rect 19628 26796 25116 26852
rect 25172 26796 25182 26852
rect 32498 26796 32508 26852
rect 32564 26796 35532 26852
rect 35588 26796 35598 26852
rect 36502 26796 36540 26852
rect 36596 26796 36606 26852
rect 38994 26796 39004 26852
rect 39060 26796 40460 26852
rect 40516 26796 40526 26852
rect 40786 26796 40796 26852
rect 40852 26796 41244 26852
rect 41300 26796 43708 26852
rect 45938 26796 45948 26852
rect 46004 26796 47628 26852
rect 47684 26796 48412 26852
rect 48468 26796 48478 26852
rect 53666 26796 53676 26852
rect 53732 26796 56476 26852
rect 56532 26796 57932 26852
rect 57988 26796 57998 26852
rect 19628 26740 19684 26796
rect 4834 26684 4844 26740
rect 4900 26684 5292 26740
rect 5348 26684 5358 26740
rect 11554 26684 11564 26740
rect 11620 26684 19684 26740
rect 33954 26684 33964 26740
rect 34020 26684 34972 26740
rect 35028 26684 35038 26740
rect 36642 26684 36652 26740
rect 36708 26684 38780 26740
rect 38836 26684 38846 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 39004 26628 39060 26796
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 4050 26572 4060 26628
rect 4116 26572 4284 26628
rect 4340 26572 4350 26628
rect 11554 26572 11564 26628
rect 11620 26572 14028 26628
rect 14084 26572 14700 26628
rect 14756 26572 18956 26628
rect 19012 26572 19022 26628
rect 23874 26572 23884 26628
rect 23940 26572 39060 26628
rect 45378 26572 45388 26628
rect 45444 26572 46620 26628
rect 46676 26572 46686 26628
rect 1698 26460 1708 26516
rect 1764 26460 1932 26516
rect 1988 26460 2268 26516
rect 2324 26460 2334 26516
rect 2930 26460 2940 26516
rect 2996 26460 4172 26516
rect 4228 26460 4238 26516
rect 10322 26460 10332 26516
rect 10388 26460 14476 26516
rect 14532 26460 14542 26516
rect 18722 26460 18732 26516
rect 18788 26460 19964 26516
rect 20020 26460 20030 26516
rect 20850 26460 20860 26516
rect 20916 26460 26012 26516
rect 26068 26460 26078 26516
rect 26226 26460 26236 26516
rect 26292 26460 26796 26516
rect 26852 26460 26862 26516
rect 34626 26460 34636 26516
rect 34692 26460 35196 26516
rect 35252 26460 37212 26516
rect 37268 26460 38556 26516
rect 38612 26460 38622 26516
rect 38770 26460 38780 26516
rect 38836 26460 40460 26516
rect 40516 26460 40526 26516
rect 43698 26460 43708 26516
rect 43764 26460 48300 26516
rect 48356 26460 48860 26516
rect 48916 26460 48926 26516
rect 4834 26348 4844 26404
rect 4900 26348 6524 26404
rect 6580 26348 6590 26404
rect 9650 26348 9660 26404
rect 9716 26348 11452 26404
rect 11508 26348 12124 26404
rect 12180 26348 13244 26404
rect 13300 26348 14140 26404
rect 14196 26348 14206 26404
rect 22530 26348 22540 26404
rect 22596 26348 22764 26404
rect 22820 26348 24892 26404
rect 24948 26348 24958 26404
rect 28466 26348 28476 26404
rect 28532 26348 29484 26404
rect 29540 26348 30156 26404
rect 30212 26348 30222 26404
rect 33954 26348 33964 26404
rect 34020 26348 40348 26404
rect 40404 26348 40414 26404
rect 43586 26348 43596 26404
rect 43652 26348 45500 26404
rect 45556 26348 46060 26404
rect 46116 26348 46126 26404
rect 3378 26236 3388 26292
rect 3444 26236 4284 26292
rect 4340 26236 5404 26292
rect 5460 26236 5470 26292
rect 9762 26236 9772 26292
rect 9828 26236 11004 26292
rect 11060 26236 13468 26292
rect 13524 26236 13534 26292
rect 18722 26236 18732 26292
rect 18788 26236 19068 26292
rect 19124 26236 20972 26292
rect 21028 26236 21038 26292
rect 22082 26236 22092 26292
rect 22148 26236 23548 26292
rect 23604 26236 23614 26292
rect 26002 26236 26012 26292
rect 26068 26236 26908 26292
rect 26964 26236 26974 26292
rect 27346 26236 27356 26292
rect 27412 26236 29372 26292
rect 29428 26236 29438 26292
rect 29698 26236 29708 26292
rect 29764 26236 30156 26292
rect 30212 26236 30222 26292
rect 31938 26236 31948 26292
rect 32004 26236 33740 26292
rect 33796 26236 33806 26292
rect 35410 26236 35420 26292
rect 35476 26236 36988 26292
rect 37044 26236 37054 26292
rect 38994 26236 39004 26292
rect 39060 26236 39788 26292
rect 39844 26236 40124 26292
rect 40180 26236 40190 26292
rect 41010 26236 41020 26292
rect 41076 26236 41916 26292
rect 41972 26236 41982 26292
rect 45602 26236 45612 26292
rect 45668 26236 45948 26292
rect 46004 26236 46732 26292
rect 46788 26236 48300 26292
rect 48356 26236 48366 26292
rect 56690 26236 56700 26292
rect 56756 26236 56924 26292
rect 56980 26236 57596 26292
rect 57652 26236 57662 26292
rect 29708 26180 29764 26236
rect 2482 26124 2492 26180
rect 2548 26124 2828 26180
rect 2884 26124 3276 26180
rect 3332 26124 3342 26180
rect 4946 26124 4956 26180
rect 5012 26124 5964 26180
rect 6020 26124 7308 26180
rect 7364 26124 8540 26180
rect 8596 26124 8606 26180
rect 9202 26124 9212 26180
rect 9268 26124 11452 26180
rect 11508 26124 11518 26180
rect 12450 26124 12460 26180
rect 12516 26124 12908 26180
rect 12964 26124 13916 26180
rect 13972 26124 13982 26180
rect 20066 26124 20076 26180
rect 20132 26124 20524 26180
rect 20580 26124 20590 26180
rect 27570 26124 27580 26180
rect 27636 26124 28476 26180
rect 28532 26124 28542 26180
rect 29138 26124 29148 26180
rect 29204 26124 29764 26180
rect 34962 26124 34972 26180
rect 35028 26124 36652 26180
rect 36708 26124 36718 26180
rect 39890 26124 39900 26180
rect 39956 26124 42364 26180
rect 42420 26124 43036 26180
rect 43092 26124 43876 26180
rect 49410 26124 49420 26180
rect 49476 26124 49868 26180
rect 49924 26124 50540 26180
rect 50596 26124 50606 26180
rect 3276 26068 3332 26124
rect 43820 26068 43876 26124
rect 3276 26012 6748 26068
rect 6804 26012 10220 26068
rect 10276 26012 10668 26068
rect 10724 26012 10734 26068
rect 14242 26012 14252 26068
rect 14308 26012 16492 26068
rect 16548 26012 16558 26068
rect 25666 26012 25676 26068
rect 25732 26012 27132 26068
rect 27188 26012 27524 26068
rect 34850 26012 34860 26068
rect 34916 26012 40684 26068
rect 40740 26012 41692 26068
rect 41748 26012 41758 26068
rect 43810 26012 43820 26068
rect 43876 26012 43886 26068
rect 53666 26012 53676 26068
rect 53732 26012 54348 26068
rect 54404 26012 54414 26068
rect 27468 25956 27524 26012
rect 10434 25900 10444 25956
rect 10500 25900 10892 25956
rect 10948 25900 10958 25956
rect 22978 25900 22988 25956
rect 23044 25900 26908 25956
rect 27458 25900 27468 25956
rect 27524 25900 27534 25956
rect 28354 25900 28364 25956
rect 28420 25900 29372 25956
rect 29428 25900 29596 25956
rect 29652 25900 30380 25956
rect 30436 25900 30446 25956
rect 38882 25900 38892 25956
rect 38948 25900 43148 25956
rect 43204 25900 44268 25956
rect 44324 25900 44334 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 26852 25844 26908 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 2930 25788 2940 25844
rect 2996 25788 3500 25844
rect 3556 25788 4060 25844
rect 4116 25788 4126 25844
rect 7858 25788 7868 25844
rect 7924 25788 12236 25844
rect 12292 25788 12572 25844
rect 12628 25788 12638 25844
rect 22754 25788 22764 25844
rect 22820 25788 24668 25844
rect 24724 25788 24734 25844
rect 26852 25788 28476 25844
rect 28532 25788 28542 25844
rect 35858 25788 35868 25844
rect 35924 25788 36428 25844
rect 36484 25788 36494 25844
rect 39666 25788 39676 25844
rect 39732 25788 40236 25844
rect 40292 25788 40302 25844
rect 4274 25676 4284 25732
rect 4340 25676 6300 25732
rect 6356 25676 9100 25732
rect 9156 25676 9166 25732
rect 19618 25676 19628 25732
rect 19684 25676 21868 25732
rect 21924 25676 23660 25732
rect 23716 25676 23726 25732
rect 26450 25676 26460 25732
rect 26516 25676 39228 25732
rect 39284 25676 40124 25732
rect 40180 25676 40190 25732
rect 1810 25564 1820 25620
rect 1876 25564 9660 25620
rect 9716 25564 9726 25620
rect 11666 25564 11676 25620
rect 11732 25564 18620 25620
rect 18676 25564 18686 25620
rect 23538 25564 23548 25620
rect 23604 25564 29148 25620
rect 29204 25564 29214 25620
rect 33170 25564 33180 25620
rect 33236 25564 33964 25620
rect 34020 25564 34030 25620
rect 34290 25564 34300 25620
rect 34356 25564 34748 25620
rect 34804 25564 34814 25620
rect 36978 25564 36988 25620
rect 37044 25564 37436 25620
rect 37492 25564 37502 25620
rect 41458 25564 41468 25620
rect 41524 25564 42364 25620
rect 42420 25564 42430 25620
rect 50530 25564 50540 25620
rect 50596 25564 51324 25620
rect 51380 25564 51390 25620
rect 2258 25452 2268 25508
rect 2324 25452 7868 25508
rect 7924 25452 7934 25508
rect 11778 25452 11788 25508
rect 11844 25452 12348 25508
rect 12404 25452 12414 25508
rect 12562 25452 12572 25508
rect 12628 25452 13132 25508
rect 13188 25452 13198 25508
rect 14018 25452 14028 25508
rect 14084 25452 15372 25508
rect 15428 25452 18396 25508
rect 18452 25452 18462 25508
rect 24658 25452 24668 25508
rect 24724 25452 25116 25508
rect 25172 25452 25182 25508
rect 27234 25452 27244 25508
rect 27300 25452 28476 25508
rect 28532 25452 30268 25508
rect 30324 25452 30334 25508
rect 32834 25452 32844 25508
rect 32900 25452 33068 25508
rect 33124 25452 33516 25508
rect 33572 25452 33582 25508
rect 42802 25452 42812 25508
rect 42868 25452 43932 25508
rect 43988 25452 43998 25508
rect 49186 25452 49196 25508
rect 49252 25452 49420 25508
rect 49476 25452 49486 25508
rect 50754 25452 50764 25508
rect 50820 25452 53900 25508
rect 53956 25452 54572 25508
rect 54628 25452 54638 25508
rect 4050 25340 4060 25396
rect 4116 25340 4956 25396
rect 5012 25340 5022 25396
rect 9314 25340 9324 25396
rect 9380 25340 9996 25396
rect 10052 25340 11620 25396
rect 25778 25340 25788 25396
rect 25844 25340 28364 25396
rect 28420 25340 30380 25396
rect 30436 25340 31836 25396
rect 31892 25340 31902 25396
rect 32050 25340 32060 25396
rect 32116 25340 33292 25396
rect 33348 25340 37884 25396
rect 37940 25340 37950 25396
rect 44930 25340 44940 25396
rect 44996 25340 45500 25396
rect 45556 25340 45566 25396
rect 46610 25340 46620 25396
rect 46676 25340 47180 25396
rect 47236 25340 47740 25396
rect 47796 25340 47806 25396
rect 48402 25340 48412 25396
rect 48468 25340 50876 25396
rect 50932 25340 50942 25396
rect 56018 25340 56028 25396
rect 56084 25340 57260 25396
rect 57316 25340 57326 25396
rect 11564 25284 11620 25340
rect 2370 25228 2380 25284
rect 2436 25228 3164 25284
rect 3220 25228 3612 25284
rect 3668 25228 3678 25284
rect 4274 25228 4284 25284
rect 4340 25228 4844 25284
rect 4900 25228 4910 25284
rect 10434 25228 10444 25284
rect 10500 25228 11340 25284
rect 11396 25228 11406 25284
rect 11554 25228 11564 25284
rect 11620 25228 11630 25284
rect 20738 25228 20748 25284
rect 20804 25228 22316 25284
rect 22372 25228 22382 25284
rect 23538 25228 23548 25284
rect 23604 25228 26460 25284
rect 26516 25228 26526 25284
rect 31154 25228 31164 25284
rect 31220 25228 32284 25284
rect 32340 25228 32508 25284
rect 32564 25228 32574 25284
rect 35298 25228 35308 25284
rect 35364 25228 35756 25284
rect 35812 25228 39228 25284
rect 39284 25228 39294 25284
rect 42130 25228 42140 25284
rect 42196 25228 42364 25284
rect 42420 25228 43260 25284
rect 43316 25228 44044 25284
rect 44100 25228 44380 25284
rect 44436 25228 44604 25284
rect 44660 25228 44670 25284
rect 45602 25228 45612 25284
rect 45668 25228 52780 25284
rect 52836 25228 52846 25284
rect 4284 25172 4340 25228
rect 2706 25116 2716 25172
rect 2772 25116 4340 25172
rect 5618 25116 5628 25172
rect 5684 25116 5740 25172
rect 5796 25116 5806 25172
rect 10210 25116 10220 25172
rect 10276 25116 10780 25172
rect 10836 25116 16268 25172
rect 16324 25116 16334 25172
rect 20178 25116 20188 25172
rect 20244 25116 21420 25172
rect 21476 25116 21486 25172
rect 29810 25116 29820 25172
rect 29876 25116 31052 25172
rect 31108 25116 31948 25172
rect 32004 25116 32014 25172
rect 32946 25116 32956 25172
rect 33012 25116 33964 25172
rect 34020 25116 34030 25172
rect 34290 25116 34300 25172
rect 34356 25116 35084 25172
rect 35140 25116 35150 25172
rect 36082 25116 36092 25172
rect 36148 25116 41132 25172
rect 41188 25116 41198 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 6066 25004 6076 25060
rect 6132 25004 13692 25060
rect 13748 25004 13758 25060
rect 18946 25004 18956 25060
rect 19012 25004 19404 25060
rect 19460 25004 19470 25060
rect 28242 25004 28252 25060
rect 28308 25004 32172 25060
rect 32228 25004 32238 25060
rect 32722 25004 32732 25060
rect 32788 25004 42252 25060
rect 42308 25004 42318 25060
rect 3714 24892 3724 24948
rect 3780 24892 3836 24948
rect 3892 24892 3902 24948
rect 12226 24892 12236 24948
rect 12292 24892 14140 24948
rect 14196 24892 14924 24948
rect 14980 24892 14990 24948
rect 15698 24892 15708 24948
rect 15764 24892 16604 24948
rect 16660 24892 16670 24948
rect 18722 24892 18732 24948
rect 18788 24892 20860 24948
rect 20916 24892 20926 24948
rect 31826 24892 31836 24948
rect 31892 24892 32060 24948
rect 32116 24892 32126 24948
rect 33842 24892 33852 24948
rect 33908 24892 38668 24948
rect 47842 24892 47852 24948
rect 47908 24892 48636 24948
rect 48692 24892 49980 24948
rect 50036 24892 50046 24948
rect 56242 24892 56252 24948
rect 56308 24892 57484 24948
rect 57540 24892 57550 24948
rect 38612 24836 38668 24892
rect 7410 24780 7420 24836
rect 7476 24780 8876 24836
rect 8932 24780 10444 24836
rect 10500 24780 10510 24836
rect 27570 24780 27580 24836
rect 27636 24780 29484 24836
rect 29540 24780 29932 24836
rect 29988 24780 32844 24836
rect 32900 24780 34860 24836
rect 34916 24780 34926 24836
rect 38612 24780 51884 24836
rect 51940 24780 51950 24836
rect 55122 24780 55132 24836
rect 55188 24780 55580 24836
rect 55636 24780 55646 24836
rect 3938 24668 3948 24724
rect 4004 24668 4732 24724
rect 4788 24668 6972 24724
rect 7028 24668 8092 24724
rect 8148 24668 8158 24724
rect 9986 24668 9996 24724
rect 10052 24668 11676 24724
rect 11732 24668 11742 24724
rect 24658 24668 24668 24724
rect 24724 24668 26236 24724
rect 26292 24668 26302 24724
rect 31266 24668 31276 24724
rect 31332 24668 31724 24724
rect 31780 24668 34188 24724
rect 34244 24668 34254 24724
rect 34962 24668 34972 24724
rect 35028 24668 36316 24724
rect 36372 24668 38780 24724
rect 38836 24668 38846 24724
rect 45378 24668 45388 24724
rect 45444 24668 47964 24724
rect 48020 24668 48030 24724
rect 48738 24668 48748 24724
rect 48804 24668 49756 24724
rect 49812 24668 49822 24724
rect 57138 24668 57148 24724
rect 57204 24668 57820 24724
rect 57876 24668 57886 24724
rect 19282 24556 19292 24612
rect 19348 24556 20524 24612
rect 20580 24556 21868 24612
rect 21924 24556 21934 24612
rect 31378 24556 31388 24612
rect 31444 24556 34524 24612
rect 34580 24556 34590 24612
rect 53218 24556 53228 24612
rect 53284 24556 58044 24612
rect 58100 24556 58110 24612
rect 13990 24444 14028 24500
rect 14084 24444 14094 24500
rect 26198 24444 26236 24500
rect 26292 24444 26302 24500
rect 28018 24444 28028 24500
rect 28084 24444 28588 24500
rect 28644 24444 28654 24500
rect 37762 24444 37772 24500
rect 37828 24444 39900 24500
rect 39956 24444 39966 24500
rect 46050 24444 46060 24500
rect 46116 24444 46844 24500
rect 46900 24444 46910 24500
rect 8372 24332 10220 24388
rect 10276 24332 11452 24388
rect 11508 24332 11518 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 6300 24220 7924 24276
rect 8306 24220 8316 24276
rect 8372 24220 8428 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 38612 24220 47516 24276
rect 47572 24220 47582 24276
rect 6300 24164 6356 24220
rect 7868 24164 7924 24220
rect 38612 24164 38668 24220
rect 3490 24108 3500 24164
rect 3556 24108 6356 24164
rect 6514 24108 6524 24164
rect 6580 24108 7308 24164
rect 7364 24108 7644 24164
rect 7700 24108 7710 24164
rect 7868 24108 9884 24164
rect 9940 24108 10556 24164
rect 10612 24108 10622 24164
rect 17154 24108 17164 24164
rect 17220 24108 19572 24164
rect 25890 24108 25900 24164
rect 25956 24108 25966 24164
rect 26852 24108 38668 24164
rect 39442 24108 39452 24164
rect 39508 24108 41132 24164
rect 41188 24108 41692 24164
rect 41748 24108 41758 24164
rect 19516 24052 19572 24108
rect 25900 24052 25956 24108
rect 1586 23996 1596 24052
rect 1652 23996 3724 24052
rect 3780 23996 3790 24052
rect 5730 23996 5740 24052
rect 5796 23996 9772 24052
rect 9828 23996 9838 24052
rect 10434 23996 10444 24052
rect 10500 23996 13020 24052
rect 13076 23996 13086 24052
rect 18274 23996 18284 24052
rect 18340 23996 19068 24052
rect 19124 23996 19134 24052
rect 19506 23996 19516 24052
rect 19572 23996 20524 24052
rect 20580 23996 25956 24052
rect 26786 23996 26796 24052
rect 26852 23996 26908 24108
rect 32386 23996 32396 24052
rect 32452 23996 36092 24052
rect 36148 23996 37772 24052
rect 37828 23996 37838 24052
rect 38210 23996 38220 24052
rect 38276 23996 43932 24052
rect 43988 23996 44380 24052
rect 44436 23996 45052 24052
rect 45108 23996 45118 24052
rect 7074 23884 7084 23940
rect 7140 23884 8652 23940
rect 8708 23884 8718 23940
rect 11218 23884 11228 23940
rect 11284 23884 14252 23940
rect 14308 23884 14318 23940
rect 16146 23884 16156 23940
rect 16212 23884 20188 23940
rect 20244 23884 20254 23940
rect 21410 23884 21420 23940
rect 21476 23884 24444 23940
rect 24500 23884 25452 23940
rect 25508 23884 25518 23940
rect 28466 23884 28476 23940
rect 28532 23884 29596 23940
rect 29652 23884 29662 23940
rect 30930 23884 30940 23940
rect 30996 23884 31276 23940
rect 31332 23884 31342 23940
rect 36194 23884 36204 23940
rect 36260 23884 37548 23940
rect 37604 23884 37614 23940
rect 38322 23884 38332 23940
rect 38388 23884 40908 23940
rect 40964 23884 42028 23940
rect 42084 23884 42094 23940
rect 42914 23884 42924 23940
rect 42980 23884 45836 23940
rect 45892 23884 45902 23940
rect 4946 23772 4956 23828
rect 5012 23772 8204 23828
rect 8260 23772 8270 23828
rect 10546 23772 10556 23828
rect 10612 23772 11004 23828
rect 11060 23772 11676 23828
rect 11732 23772 12460 23828
rect 12516 23772 12526 23828
rect 17602 23772 17612 23828
rect 17668 23772 19404 23828
rect 19460 23772 22540 23828
rect 22596 23772 22606 23828
rect 26562 23772 26572 23828
rect 26628 23772 26796 23828
rect 26852 23772 26862 23828
rect 36754 23772 36764 23828
rect 36820 23772 38220 23828
rect 38276 23772 38286 23828
rect 38994 23772 39004 23828
rect 39060 23772 40572 23828
rect 40628 23772 40638 23828
rect 41458 23772 41468 23828
rect 41524 23772 42476 23828
rect 42532 23772 42542 23828
rect 46498 23772 46508 23828
rect 46564 23772 52668 23828
rect 52724 23772 53004 23828
rect 53060 23772 53070 23828
rect 55122 23772 55132 23828
rect 55188 23772 56364 23828
rect 56420 23772 56430 23828
rect 8092 23660 8988 23716
rect 9044 23660 9054 23716
rect 10770 23660 10780 23716
rect 10836 23660 11900 23716
rect 11956 23660 11966 23716
rect 16034 23660 16044 23716
rect 16100 23660 16492 23716
rect 16548 23660 16828 23716
rect 16884 23660 18060 23716
rect 18116 23660 18126 23716
rect 19618 23660 19628 23716
rect 19684 23660 20748 23716
rect 20804 23660 22204 23716
rect 22260 23660 22270 23716
rect 22978 23660 22988 23716
rect 23044 23660 24220 23716
rect 24276 23660 25676 23716
rect 25732 23660 25742 23716
rect 30146 23660 30156 23716
rect 30212 23660 32396 23716
rect 32452 23660 32462 23716
rect 34066 23660 34076 23716
rect 34132 23660 34636 23716
rect 34692 23660 34702 23716
rect 36866 23660 36876 23716
rect 36932 23660 38444 23716
rect 38500 23660 38510 23716
rect 47170 23660 47180 23716
rect 47236 23660 47516 23716
rect 47572 23660 48972 23716
rect 49028 23660 49038 23716
rect 3602 23548 3612 23604
rect 3668 23548 6972 23604
rect 7028 23548 7868 23604
rect 7924 23548 7934 23604
rect 8092 23492 8148 23660
rect 34076 23604 34132 23660
rect 1474 23436 1484 23492
rect 1540 23436 8148 23492
rect 8316 23548 8764 23604
rect 8820 23548 13916 23604
rect 13972 23548 13982 23604
rect 23650 23548 23660 23604
rect 23716 23548 24668 23604
rect 24724 23548 24734 23604
rect 24882 23548 24892 23604
rect 24948 23548 30940 23604
rect 30996 23548 34132 23604
rect 34738 23548 34748 23604
rect 34804 23548 35868 23604
rect 35924 23548 36764 23604
rect 36820 23548 36830 23604
rect 46386 23548 46396 23604
rect 46452 23548 46956 23604
rect 47012 23548 47022 23604
rect 8316 23380 8372 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 13458 23436 13468 23492
rect 13524 23436 15148 23492
rect 15204 23436 15596 23492
rect 15652 23436 15662 23492
rect 20514 23436 20524 23492
rect 20580 23436 22428 23492
rect 22484 23436 22494 23492
rect 26898 23436 26908 23492
rect 26964 23436 27356 23492
rect 27412 23436 27422 23492
rect 30342 23436 30380 23492
rect 30436 23436 32060 23492
rect 32116 23436 32126 23492
rect 32386 23436 32396 23492
rect 32452 23436 35196 23492
rect 35252 23436 35262 23492
rect 35522 23436 35532 23492
rect 35588 23436 37324 23492
rect 37380 23436 37390 23492
rect 43810 23436 43820 23492
rect 43876 23436 45724 23492
rect 45780 23436 46284 23492
rect 46340 23436 46350 23492
rect 1026 23324 1036 23380
rect 1092 23324 5628 23380
rect 5684 23324 5694 23380
rect 7858 23324 7868 23380
rect 7924 23324 8372 23380
rect 8978 23324 8988 23380
rect 9044 23324 11228 23380
rect 11284 23324 11294 23380
rect 11778 23324 11788 23380
rect 11844 23324 13580 23380
rect 13636 23324 13646 23380
rect 14466 23324 14476 23380
rect 14532 23324 15484 23380
rect 15540 23324 15550 23380
rect 17602 23324 17612 23380
rect 17668 23324 17678 23380
rect 26562 23324 26572 23380
rect 26628 23324 32732 23380
rect 32788 23324 32798 23380
rect 32956 23324 38668 23380
rect 40002 23324 40012 23380
rect 40068 23324 49308 23380
rect 49364 23324 49374 23380
rect 17612 23268 17668 23324
rect 32956 23268 33012 23324
rect 38612 23268 38668 23324
rect 2258 23212 2268 23268
rect 2324 23212 4620 23268
rect 4676 23212 5068 23268
rect 5124 23212 5516 23268
rect 5572 23212 5582 23268
rect 8306 23212 8316 23268
rect 8372 23212 10892 23268
rect 10948 23212 10958 23268
rect 12786 23212 12796 23268
rect 12852 23212 13804 23268
rect 13860 23212 17668 23268
rect 18498 23212 18508 23268
rect 18564 23212 18956 23268
rect 19012 23212 19022 23268
rect 21970 23212 21980 23268
rect 22036 23212 22316 23268
rect 22372 23212 23100 23268
rect 23156 23212 23166 23268
rect 24546 23212 24556 23268
rect 24612 23212 24780 23268
rect 24836 23212 26124 23268
rect 26180 23212 26348 23268
rect 26404 23212 27356 23268
rect 27412 23212 27422 23268
rect 30566 23212 30604 23268
rect 30660 23212 30670 23268
rect 32162 23212 32172 23268
rect 32228 23212 33012 23268
rect 33394 23212 33404 23268
rect 33460 23212 33470 23268
rect 35074 23212 35084 23268
rect 35140 23212 35644 23268
rect 35700 23212 35710 23268
rect 36978 23212 36988 23268
rect 37044 23212 37054 23268
rect 38612 23212 44940 23268
rect 44996 23212 45006 23268
rect 51314 23212 51324 23268
rect 51380 23212 54012 23268
rect 54068 23212 54460 23268
rect 54516 23212 54526 23268
rect 6626 23100 6636 23156
rect 6692 23100 9548 23156
rect 9604 23100 9614 23156
rect 10770 23100 10780 23156
rect 10836 23100 11228 23156
rect 11284 23100 11294 23156
rect 13010 23100 13020 23156
rect 13076 23100 15484 23156
rect 15540 23100 15550 23156
rect 16930 23100 16940 23156
rect 16996 23100 18172 23156
rect 18228 23100 20636 23156
rect 20692 23100 21308 23156
rect 21364 23100 21374 23156
rect 24882 23100 24892 23156
rect 24948 23100 27468 23156
rect 27524 23100 27534 23156
rect 30678 23100 30716 23156
rect 30772 23100 30782 23156
rect 32172 23044 32228 23212
rect 23650 22988 23660 23044
rect 23716 22988 26908 23044
rect 26964 22988 26974 23044
rect 30146 22988 30156 23044
rect 30212 22988 31164 23044
rect 31220 22988 32228 23044
rect 17938 22876 17948 22932
rect 18004 22876 18732 22932
rect 18788 22876 18798 22932
rect 20738 22876 20748 22932
rect 20804 22876 24108 22932
rect 24164 22876 25900 22932
rect 25956 22876 25966 22932
rect 30146 22876 30156 22932
rect 30212 22876 32620 22932
rect 32676 22876 32686 22932
rect 20748 22820 20804 22876
rect 33404 22820 33460 23212
rect 34626 23100 34636 23156
rect 34692 23100 35532 23156
rect 35588 23100 35598 23156
rect 36988 23044 37044 23212
rect 39666 23100 39676 23156
rect 39732 23100 40348 23156
rect 40404 23100 40414 23156
rect 42578 23100 42588 23156
rect 42644 23100 43484 23156
rect 43540 23100 43550 23156
rect 53554 23100 53564 23156
rect 53620 23100 54348 23156
rect 54404 23100 54414 23156
rect 34962 22988 34972 23044
rect 35028 22988 35644 23044
rect 35700 22988 37996 23044
rect 38052 22988 38062 23044
rect 38770 22988 38780 23044
rect 38836 22988 45612 23044
rect 45668 22988 46732 23044
rect 46788 22988 46798 23044
rect 48290 22988 48300 23044
rect 48356 22988 49196 23044
rect 49252 22988 49262 23044
rect 53442 22988 53452 23044
rect 53508 22988 53788 23044
rect 53844 22988 54460 23044
rect 54516 22988 54526 23044
rect 34178 22876 34188 22932
rect 34244 22876 34636 22932
rect 34692 22876 34702 22932
rect 39778 22876 39788 22932
rect 39844 22876 40124 22932
rect 40180 22876 40796 22932
rect 40852 22876 41692 22932
rect 41748 22876 45388 22932
rect 45444 22876 45454 22932
rect 16370 22764 16380 22820
rect 16436 22764 17612 22820
rect 17668 22764 18396 22820
rect 18452 22764 20804 22820
rect 32274 22764 32284 22820
rect 32340 22764 32844 22820
rect 32900 22764 32910 22820
rect 33404 22764 33740 22820
rect 33796 22764 33806 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 28802 22652 28812 22708
rect 28868 22652 30604 22708
rect 30660 22652 31164 22708
rect 31220 22652 33852 22708
rect 33908 22652 33918 22708
rect 3714 22540 3724 22596
rect 3780 22540 23100 22596
rect 23156 22540 23166 22596
rect 2146 22428 2156 22484
rect 2212 22428 2828 22484
rect 2884 22428 2894 22484
rect 4050 22428 4060 22484
rect 4116 22428 5740 22484
rect 5796 22428 6748 22484
rect 6804 22428 6814 22484
rect 10182 22428 10220 22484
rect 10276 22428 10286 22484
rect 20178 22428 20188 22484
rect 20244 22428 21644 22484
rect 21700 22428 21710 22484
rect 32050 22428 32060 22484
rect 32116 22428 35644 22484
rect 35700 22428 35710 22484
rect 39330 22428 39340 22484
rect 39396 22428 39900 22484
rect 39956 22428 39966 22484
rect 46386 22428 46396 22484
rect 46452 22428 46732 22484
rect 46788 22428 48188 22484
rect 48244 22428 48254 22484
rect 2828 22372 2884 22428
rect 2828 22316 4844 22372
rect 4900 22316 4910 22372
rect 19506 22316 19516 22372
rect 19572 22316 19582 22372
rect 20850 22316 20860 22372
rect 20916 22316 21420 22372
rect 21476 22316 21980 22372
rect 22036 22316 22046 22372
rect 30818 22316 30828 22372
rect 30884 22316 31388 22372
rect 31444 22316 31454 22372
rect 33842 22316 33852 22372
rect 33908 22316 36540 22372
rect 36596 22316 36606 22372
rect 4060 22260 4116 22316
rect 19516 22260 19572 22316
rect 39340 22260 39396 22428
rect 44818 22316 44828 22372
rect 44884 22316 45500 22372
rect 45556 22316 45566 22372
rect 46050 22316 46060 22372
rect 46116 22316 50540 22372
rect 50596 22316 51100 22372
rect 51156 22316 51166 22372
rect 4050 22204 4060 22260
rect 4116 22204 4126 22260
rect 5058 22204 5068 22260
rect 5124 22204 5292 22260
rect 5348 22204 6412 22260
rect 6468 22204 6478 22260
rect 8372 22204 11116 22260
rect 11172 22204 11452 22260
rect 11508 22204 12012 22260
rect 12068 22204 12078 22260
rect 19516 22204 26012 22260
rect 26068 22204 26236 22260
rect 26292 22204 27580 22260
rect 27636 22204 27646 22260
rect 27906 22204 27916 22260
rect 27972 22204 39396 22260
rect 45714 22204 45724 22260
rect 45780 22204 47740 22260
rect 47796 22204 47806 22260
rect 51202 22204 51212 22260
rect 51268 22204 51996 22260
rect 52052 22204 52062 22260
rect 52210 22204 52220 22260
rect 52276 22204 53564 22260
rect 53620 22204 53630 22260
rect 8372 22148 8428 22204
rect 4162 22092 4172 22148
rect 4228 22092 8428 22148
rect 9874 22092 9884 22148
rect 9940 22092 12236 22148
rect 12292 22092 12302 22148
rect 12674 22092 12684 22148
rect 12740 22092 13132 22148
rect 13188 22092 15148 22148
rect 15204 22092 15214 22148
rect 19730 22092 19740 22148
rect 19796 22092 20636 22148
rect 20692 22092 20702 22148
rect 21644 22036 21700 22204
rect 23538 22092 23548 22148
rect 23604 22092 23772 22148
rect 23828 22092 24220 22148
rect 24276 22092 24286 22148
rect 26852 22092 28812 22148
rect 28868 22092 29372 22148
rect 29428 22092 29438 22148
rect 32722 22092 32732 22148
rect 32788 22092 33068 22148
rect 33124 22092 33134 22148
rect 35186 22092 35196 22148
rect 35252 22092 37324 22148
rect 37380 22092 37390 22148
rect 40450 22092 40460 22148
rect 40516 22092 41468 22148
rect 41524 22092 42364 22148
rect 42420 22092 42430 22148
rect 46162 22092 46172 22148
rect 46228 22092 47628 22148
rect 47684 22092 47694 22148
rect 56354 22092 56364 22148
rect 56420 22092 58156 22148
rect 58212 22092 58222 22148
rect 1810 21980 1820 22036
rect 1876 21980 12348 22036
rect 12404 21980 12414 22036
rect 17826 21980 17836 22036
rect 17892 21980 18172 22036
rect 18228 21980 18238 22036
rect 21074 21980 21084 22036
rect 21140 21980 21150 22036
rect 21634 21980 21644 22036
rect 21700 21980 21710 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 21084 21924 21140 21980
rect 2706 21868 2716 21924
rect 2772 21868 6636 21924
rect 6692 21868 6702 21924
rect 20514 21868 20524 21924
rect 20580 21868 20590 21924
rect 21084 21868 21532 21924
rect 21588 21868 21598 21924
rect 23314 21868 23324 21924
rect 23380 21868 23660 21924
rect 23716 21868 23726 21924
rect 20524 21812 20580 21868
rect 26852 21812 26908 22092
rect 35634 21980 35644 22036
rect 35700 21980 39228 22036
rect 39284 21980 39294 22036
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 33282 21868 33292 21924
rect 33348 21868 34972 21924
rect 35028 21868 35308 21924
rect 35364 21868 35374 21924
rect 36306 21868 36316 21924
rect 36372 21868 37884 21924
rect 37940 21868 39116 21924
rect 39172 21868 39182 21924
rect 2258 21756 2268 21812
rect 2324 21756 3052 21812
rect 3108 21756 6412 21812
rect 6468 21756 6860 21812
rect 6916 21756 8820 21812
rect 8978 21756 8988 21812
rect 9044 21756 9660 21812
rect 9716 21756 9726 21812
rect 15810 21756 15820 21812
rect 15876 21756 16828 21812
rect 16884 21756 18172 21812
rect 18228 21756 19516 21812
rect 19572 21756 19582 21812
rect 20300 21756 20580 21812
rect 22530 21756 22540 21812
rect 22596 21756 22876 21812
rect 22932 21756 22942 21812
rect 24658 21756 24668 21812
rect 24724 21756 25116 21812
rect 25172 21756 25182 21812
rect 25666 21756 25676 21812
rect 25732 21756 26908 21812
rect 27682 21756 27692 21812
rect 27748 21756 29148 21812
rect 29204 21756 29214 21812
rect 30818 21756 30828 21812
rect 30884 21756 32172 21812
rect 32228 21756 32238 21812
rect 35522 21756 35532 21812
rect 35588 21756 36204 21812
rect 36260 21756 37212 21812
rect 37268 21756 38220 21812
rect 38276 21756 38780 21812
rect 38836 21756 38846 21812
rect 40114 21756 40124 21812
rect 40180 21756 40572 21812
rect 40628 21756 42812 21812
rect 42868 21756 42878 21812
rect 44146 21756 44156 21812
rect 44212 21756 46676 21812
rect 46834 21756 46844 21812
rect 46900 21756 47404 21812
rect 47460 21756 47470 21812
rect 8764 21700 8820 21756
rect 20300 21700 20356 21756
rect 46620 21700 46676 21756
rect 1810 21644 1820 21700
rect 1876 21644 3948 21700
rect 4004 21644 4014 21700
rect 6178 21644 6188 21700
rect 6244 21644 7420 21700
rect 7476 21644 7486 21700
rect 8082 21644 8092 21700
rect 8148 21644 8540 21700
rect 8596 21644 8606 21700
rect 8764 21644 9100 21700
rect 9156 21644 9436 21700
rect 9492 21644 9502 21700
rect 16930 21644 16940 21700
rect 16996 21644 17724 21700
rect 17780 21644 17790 21700
rect 18834 21644 18844 21700
rect 18900 21644 20356 21700
rect 20514 21644 20524 21700
rect 20580 21644 20748 21700
rect 20804 21644 21756 21700
rect 21812 21644 23100 21700
rect 23156 21644 23166 21700
rect 26786 21644 26796 21700
rect 26852 21644 27468 21700
rect 27524 21644 27534 21700
rect 29250 21644 29260 21700
rect 29316 21644 29326 21700
rect 30566 21644 30604 21700
rect 30660 21644 30670 21700
rect 31938 21644 31948 21700
rect 32004 21644 32732 21700
rect 32788 21644 33740 21700
rect 33796 21644 33806 21700
rect 34178 21644 34188 21700
rect 34244 21644 36764 21700
rect 36820 21644 36830 21700
rect 45042 21644 45052 21700
rect 45108 21644 45948 21700
rect 46004 21644 46014 21700
rect 46620 21644 49308 21700
rect 49364 21644 49644 21700
rect 49700 21644 49710 21700
rect 50530 21644 50540 21700
rect 50596 21644 52332 21700
rect 52388 21644 52398 21700
rect 29260 21588 29316 21644
rect 2146 21532 2156 21588
rect 2212 21532 3052 21588
rect 3108 21532 4844 21588
rect 4900 21532 4910 21588
rect 5954 21532 5964 21588
rect 6020 21532 6636 21588
rect 6692 21532 6702 21588
rect 10658 21532 10668 21588
rect 10724 21532 12236 21588
rect 12292 21532 12302 21588
rect 15586 21532 15596 21588
rect 15652 21532 17836 21588
rect 17892 21532 17902 21588
rect 18274 21532 18284 21588
rect 18340 21532 20076 21588
rect 20132 21532 23212 21588
rect 23268 21532 23278 21588
rect 26310 21532 26348 21588
rect 26404 21532 26414 21588
rect 29260 21532 32956 21588
rect 33012 21532 33022 21588
rect 35858 21532 35868 21588
rect 35924 21532 37100 21588
rect 37156 21532 37166 21588
rect 39218 21532 39228 21588
rect 39284 21532 41468 21588
rect 41524 21532 41534 21588
rect 47282 21532 47292 21588
rect 47348 21532 49868 21588
rect 49924 21532 51100 21588
rect 51156 21532 51166 21588
rect 57250 21532 57260 21588
rect 57316 21532 57708 21588
rect 57764 21532 58492 21588
rect 58548 21532 58558 21588
rect 4844 21476 4900 21532
rect 18284 21476 18340 21532
rect 3154 21420 3164 21476
rect 3220 21420 3724 21476
rect 3780 21420 3948 21476
rect 4004 21420 4396 21476
rect 4452 21420 4462 21476
rect 4844 21420 5068 21476
rect 5124 21420 8988 21476
rect 9044 21420 9054 21476
rect 11666 21420 11676 21476
rect 11732 21420 15820 21476
rect 15876 21420 15886 21476
rect 17154 21420 17164 21476
rect 17220 21420 18340 21476
rect 21298 21420 21308 21476
rect 21364 21420 21756 21476
rect 21812 21420 26684 21476
rect 26740 21420 26750 21476
rect 28690 21420 28700 21476
rect 28756 21420 39788 21476
rect 39844 21420 39854 21476
rect 43922 21420 43932 21476
rect 43988 21420 44716 21476
rect 44772 21420 44782 21476
rect 56578 21420 56588 21476
rect 56644 21420 57596 21476
rect 57652 21420 57662 21476
rect 8194 21308 8204 21364
rect 8260 21308 8540 21364
rect 8596 21308 12124 21364
rect 12180 21308 12572 21364
rect 12628 21308 13692 21364
rect 13748 21308 13758 21364
rect 22194 21308 22204 21364
rect 22260 21308 26908 21364
rect 30034 21308 30044 21364
rect 30100 21308 30492 21364
rect 30548 21308 30558 21364
rect 34066 21308 34076 21364
rect 34132 21308 36372 21364
rect 38882 21308 38892 21364
rect 38948 21308 40348 21364
rect 40404 21308 40414 21364
rect 40674 21308 40684 21364
rect 40740 21308 42028 21364
rect 42084 21308 43484 21364
rect 43540 21308 44492 21364
rect 44548 21308 44558 21364
rect 49634 21308 49644 21364
rect 49700 21308 51324 21364
rect 51380 21308 52108 21364
rect 52164 21308 52174 21364
rect 54338 21308 54348 21364
rect 54404 21308 54796 21364
rect 54852 21308 55356 21364
rect 55412 21308 56476 21364
rect 56532 21308 57652 21364
rect 8194 21196 8204 21252
rect 8260 21196 8428 21252
rect 8484 21196 8494 21252
rect 12124 21196 13132 21252
rect 13188 21196 13198 21252
rect 21970 21196 21980 21252
rect 22036 21196 22652 21252
rect 22708 21196 22718 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 12124 21140 12180 21196
rect 26852 21140 26908 21308
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 7970 21084 7980 21140
rect 8036 21084 8428 21140
rect 8530 21084 8540 21140
rect 8596 21084 12124 21140
rect 12180 21084 12190 21140
rect 12338 21084 12348 21140
rect 12404 21084 18284 21140
rect 18340 21084 18350 21140
rect 22418 21084 22428 21140
rect 22484 21084 22494 21140
rect 26852 21084 28756 21140
rect 8372 21028 8428 21084
rect 4946 20972 4956 21028
rect 5012 20972 5516 21028
rect 5572 20972 7308 21028
rect 7364 20972 7374 21028
rect 8372 20972 12404 21028
rect 13458 20972 13468 21028
rect 13524 20972 13916 21028
rect 13972 20972 13982 21028
rect 16146 20972 16156 21028
rect 16212 20972 18732 21028
rect 18788 20972 18798 21028
rect 12348 20916 12404 20972
rect 2706 20860 2716 20916
rect 2772 20860 4060 20916
rect 4116 20860 4126 20916
rect 5618 20860 5628 20916
rect 5684 20860 6412 20916
rect 6468 20860 6478 20916
rect 9762 20860 9772 20916
rect 9828 20860 10332 20916
rect 10388 20860 10398 20916
rect 12338 20860 12348 20916
rect 12404 20860 14140 20916
rect 14196 20860 15260 20916
rect 15316 20860 15326 20916
rect 18050 20860 18060 20916
rect 18116 20860 20188 20916
rect 20244 20860 20254 20916
rect 22428 20804 22484 21084
rect 28700 21028 28756 21084
rect 36316 21028 36372 21308
rect 57596 21252 57652 21308
rect 39218 21196 39228 21252
rect 39284 21196 41916 21252
rect 41972 21196 42588 21252
rect 42644 21196 43148 21252
rect 43204 21196 43214 21252
rect 57586 21196 57596 21252
rect 57652 21196 57662 21252
rect 36754 21084 36764 21140
rect 36820 21084 43708 21140
rect 43764 21084 43774 21140
rect 46610 21084 46620 21140
rect 46676 21084 47180 21140
rect 47236 21084 47852 21140
rect 47908 21084 47918 21140
rect 26002 20972 26012 21028
rect 26068 20972 27132 21028
rect 27188 20972 27804 21028
rect 27860 20972 27870 21028
rect 28690 20972 28700 21028
rect 28756 20972 28766 21028
rect 31602 20972 31612 21028
rect 31668 20972 34188 21028
rect 34244 20972 34254 21028
rect 34738 20972 34748 21028
rect 34804 20972 35756 21028
rect 35812 20972 35822 21028
rect 36316 20972 38668 21028
rect 39778 20972 39788 21028
rect 39844 20972 40012 21028
rect 40068 20972 40236 21028
rect 40292 20972 40684 21028
rect 40740 20972 40750 21028
rect 24322 20860 24332 20916
rect 24388 20860 28700 20916
rect 28756 20860 28766 20916
rect 29026 20860 29036 20916
rect 29092 20860 29708 20916
rect 29764 20860 32508 20916
rect 32564 20860 34860 20916
rect 34916 20860 34926 20916
rect 36082 20860 36092 20916
rect 36148 20860 38108 20916
rect 38164 20860 38174 20916
rect 38612 20860 38668 20972
rect 38724 20860 38734 20916
rect 6850 20748 6860 20804
rect 6916 20748 7308 20804
rect 7364 20748 7980 20804
rect 8036 20748 8046 20804
rect 8866 20748 8876 20804
rect 8932 20748 9436 20804
rect 9492 20748 10892 20804
rect 10948 20748 10958 20804
rect 11778 20748 11788 20804
rect 11844 20748 12236 20804
rect 12292 20748 12302 20804
rect 17714 20748 17724 20804
rect 17780 20748 22092 20804
rect 22148 20748 22158 20804
rect 22428 20748 27188 20804
rect 27318 20748 27356 20804
rect 27412 20748 27422 20804
rect 28578 20748 28588 20804
rect 28644 20748 29260 20804
rect 29316 20748 29326 20804
rect 33394 20748 33404 20804
rect 33460 20748 33628 20804
rect 33684 20748 33694 20804
rect 34178 20748 34188 20804
rect 34244 20748 34636 20804
rect 34692 20748 34702 20804
rect 36642 20748 36652 20804
rect 36708 20748 37548 20804
rect 37604 20748 37614 20804
rect 41010 20748 41020 20804
rect 41076 20748 42364 20804
rect 42420 20748 43036 20804
rect 43092 20748 43102 20804
rect 27132 20692 27188 20748
rect 6178 20636 6188 20692
rect 6244 20636 8988 20692
rect 9044 20636 9054 20692
rect 10556 20636 21980 20692
rect 22036 20636 22046 20692
rect 23202 20636 23212 20692
rect 23268 20636 23660 20692
rect 23716 20636 23726 20692
rect 24994 20636 25004 20692
rect 25060 20636 26796 20692
rect 26852 20636 26862 20692
rect 27122 20636 27132 20692
rect 27188 20636 33908 20692
rect 54674 20636 54684 20692
rect 54740 20636 56028 20692
rect 56084 20636 58044 20692
rect 58100 20636 58110 20692
rect 8418 20524 8428 20580
rect 8484 20524 10332 20580
rect 10388 20524 10398 20580
rect 10556 20356 10612 20636
rect 33852 20580 33908 20636
rect 13346 20524 13356 20580
rect 13412 20524 13804 20580
rect 13860 20524 13870 20580
rect 18274 20524 18284 20580
rect 18340 20524 21756 20580
rect 21812 20524 21822 20580
rect 23314 20524 23324 20580
rect 23380 20524 24220 20580
rect 24276 20524 24286 20580
rect 25442 20524 25452 20580
rect 25508 20524 26012 20580
rect 26068 20524 26078 20580
rect 26898 20524 26908 20580
rect 26964 20524 28364 20580
rect 28420 20524 28430 20580
rect 33842 20524 33852 20580
rect 33908 20524 35868 20580
rect 35924 20524 35934 20580
rect 36530 20524 36540 20580
rect 36596 20524 38556 20580
rect 38612 20524 39452 20580
rect 39508 20524 39518 20580
rect 25106 20412 25116 20468
rect 25172 20412 26796 20468
rect 26852 20412 31836 20468
rect 31892 20412 33404 20468
rect 33460 20412 34076 20468
rect 34132 20412 34142 20468
rect 53666 20412 53676 20468
rect 53732 20412 55020 20468
rect 55076 20412 58380 20468
rect 58436 20412 58446 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 1922 20300 1932 20356
rect 1988 20300 4508 20356
rect 4564 20300 4574 20356
rect 4946 20300 4956 20356
rect 5012 20300 6636 20356
rect 6692 20300 6702 20356
rect 7970 20300 7980 20356
rect 8036 20300 10612 20356
rect 22082 20300 22092 20356
rect 22148 20300 22988 20356
rect 23044 20300 23054 20356
rect 23650 20300 23660 20356
rect 23716 20300 24444 20356
rect 24500 20300 24510 20356
rect 26898 20300 26908 20356
rect 26964 20300 27244 20356
rect 27300 20300 27310 20356
rect 28130 20300 28140 20356
rect 28196 20300 28364 20356
rect 28420 20300 28756 20356
rect 34626 20300 34636 20356
rect 34692 20300 39004 20356
rect 39060 20300 39070 20356
rect 40562 20300 40572 20356
rect 40628 20300 40796 20356
rect 40852 20300 40862 20356
rect 6066 20188 6076 20244
rect 6132 20188 7196 20244
rect 7252 20188 11116 20244
rect 11172 20188 11182 20244
rect 20178 20188 20188 20244
rect 20244 20188 23548 20244
rect 23604 20188 24668 20244
rect 24724 20188 24734 20244
rect 27468 20188 28084 20244
rect 27468 20132 27524 20188
rect 28028 20132 28084 20188
rect 28700 20132 28756 20300
rect 28914 20188 28924 20244
rect 28980 20188 29820 20244
rect 29876 20188 29886 20244
rect 32722 20188 32732 20244
rect 32788 20188 33516 20244
rect 33572 20188 35532 20244
rect 35588 20188 35598 20244
rect 37986 20188 37996 20244
rect 38052 20188 46060 20244
rect 46116 20188 46508 20244
rect 46564 20188 48300 20244
rect 48356 20188 48366 20244
rect 56466 20188 56476 20244
rect 56532 20188 56542 20244
rect 56476 20132 56532 20188
rect 2370 20076 2380 20132
rect 2436 20076 6860 20132
rect 6916 20076 6926 20132
rect 16706 20076 16716 20132
rect 16772 20076 19180 20132
rect 19236 20076 19246 20132
rect 27234 20076 27244 20132
rect 27300 20076 27524 20132
rect 27682 20076 27692 20132
rect 27748 20076 27804 20132
rect 27860 20076 27870 20132
rect 28018 20076 28028 20132
rect 28084 20076 28476 20132
rect 28532 20076 28542 20132
rect 28700 20076 31388 20132
rect 31444 20076 31836 20132
rect 31892 20076 31902 20132
rect 32946 20076 32956 20132
rect 33012 20076 33852 20132
rect 33908 20076 35084 20132
rect 35140 20076 35150 20132
rect 35970 20076 35980 20132
rect 36036 20076 36540 20132
rect 36596 20076 36606 20132
rect 36754 20076 36764 20132
rect 36820 20076 37548 20132
rect 37604 20076 37614 20132
rect 40114 20076 40124 20132
rect 40180 20076 40460 20132
rect 40516 20076 40526 20132
rect 50306 20076 50316 20132
rect 50372 20076 53788 20132
rect 53844 20076 53854 20132
rect 56476 20076 57932 20132
rect 57988 20076 57998 20132
rect 3042 19964 3052 20020
rect 3108 19964 3500 20020
rect 3556 19964 4284 20020
rect 4340 19964 7084 20020
rect 7140 19964 7150 20020
rect 10658 19964 10668 20020
rect 10724 19964 11564 20020
rect 11620 19964 11630 20020
rect 12002 19964 12012 20020
rect 12068 19964 12572 20020
rect 12628 19964 12638 20020
rect 15586 19964 15596 20020
rect 15652 19964 16492 20020
rect 16548 19964 16558 20020
rect 22642 19964 22652 20020
rect 22708 19964 28700 20020
rect 28756 19964 30156 20020
rect 30212 19964 30222 20020
rect 31714 19964 31724 20020
rect 31780 19964 32284 20020
rect 32340 19964 32350 20020
rect 32834 19964 32844 20020
rect 32900 19964 36876 20020
rect 36932 19964 42588 20020
rect 42644 19964 42654 20020
rect 54460 19964 55692 20020
rect 55748 19964 56812 20020
rect 56868 19964 57820 20020
rect 57876 19964 57886 20020
rect 54460 19908 54516 19964
rect 1810 19852 1820 19908
rect 1876 19852 3612 19908
rect 3668 19852 3678 19908
rect 14018 19852 14028 19908
rect 14084 19852 16268 19908
rect 16324 19852 16334 19908
rect 17042 19852 17052 19908
rect 17108 19852 18508 19908
rect 18564 19852 19068 19908
rect 19124 19852 19404 19908
rect 19460 19852 19470 19908
rect 23090 19852 23100 19908
rect 23156 19852 27692 19908
rect 27748 19852 28028 19908
rect 28084 19852 28094 19908
rect 52882 19852 52892 19908
rect 52948 19852 54460 19908
rect 54516 19852 54526 19908
rect 55010 19852 55020 19908
rect 55076 19852 56028 19908
rect 56084 19852 58156 19908
rect 58212 19852 58222 19908
rect 1138 19740 1148 19796
rect 1204 19740 22204 19796
rect 22260 19740 23212 19796
rect 23268 19740 23278 19796
rect 23762 19740 23772 19796
rect 23828 19740 26460 19796
rect 26516 19740 26526 19796
rect 29250 19740 29260 19796
rect 29316 19740 29820 19796
rect 29876 19740 29886 19796
rect 32050 19740 32060 19796
rect 32116 19740 32508 19796
rect 32564 19740 34524 19796
rect 34580 19740 34590 19796
rect 34962 19740 34972 19796
rect 35028 19740 35756 19796
rect 35812 19740 36092 19796
rect 36148 19740 36428 19796
rect 36484 19740 36494 19796
rect 53778 19740 53788 19796
rect 53844 19740 54012 19796
rect 54068 19740 57260 19796
rect 57316 19740 57326 19796
rect 5170 19628 5180 19684
rect 5236 19628 6636 19684
rect 6692 19628 6702 19684
rect 15250 19628 15260 19684
rect 15316 19628 18396 19684
rect 18452 19628 18462 19684
rect 19058 19628 19068 19684
rect 19124 19628 19292 19684
rect 19348 19628 19358 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 25666 19516 25676 19572
rect 25732 19516 26348 19572
rect 26404 19516 27804 19572
rect 27860 19516 27870 19572
rect 34402 19516 34412 19572
rect 34468 19516 35028 19572
rect 4162 19404 4172 19460
rect 4228 19404 7532 19460
rect 7588 19404 7598 19460
rect 31126 19404 31164 19460
rect 31220 19404 31230 19460
rect 5058 19292 5068 19348
rect 5124 19292 5852 19348
rect 5908 19292 5918 19348
rect 6514 19292 6524 19348
rect 6580 19292 7980 19348
rect 8036 19292 10108 19348
rect 10164 19292 10174 19348
rect 10966 19292 11004 19348
rect 11060 19292 11070 19348
rect 11890 19292 11900 19348
rect 11956 19292 12572 19348
rect 12628 19292 14364 19348
rect 14420 19292 14430 19348
rect 28774 19292 28812 19348
rect 28868 19292 28878 19348
rect 29474 19292 29484 19348
rect 29540 19292 30268 19348
rect 30324 19292 30334 19348
rect 30930 19292 30940 19348
rect 30996 19292 32396 19348
rect 32452 19292 33964 19348
rect 34020 19292 34748 19348
rect 34804 19292 34814 19348
rect 34972 19236 35028 19516
rect 39442 19404 39452 19460
rect 39508 19404 46060 19460
rect 46116 19404 46126 19460
rect 39330 19292 39340 19348
rect 39396 19292 39676 19348
rect 39732 19292 41020 19348
rect 41076 19292 41244 19348
rect 41300 19292 41310 19348
rect 3602 19180 3612 19236
rect 3668 19180 4956 19236
rect 5012 19180 5022 19236
rect 7522 19180 7532 19236
rect 7588 19180 12180 19236
rect 22306 19180 22316 19236
rect 22372 19180 23100 19236
rect 23156 19180 23166 19236
rect 24882 19180 24892 19236
rect 24948 19180 26460 19236
rect 26516 19180 27020 19236
rect 27076 19180 27086 19236
rect 34850 19180 34860 19236
rect 34916 19180 35028 19236
rect 36194 19180 36204 19236
rect 36260 19180 37884 19236
rect 37940 19180 37950 19236
rect 40338 19180 40348 19236
rect 40404 19180 40908 19236
rect 40964 19180 41468 19236
rect 41524 19180 41534 19236
rect 42914 19180 42924 19236
rect 42980 19180 44044 19236
rect 44100 19180 44110 19236
rect 48626 19180 48636 19236
rect 48692 19180 49084 19236
rect 49140 19180 50092 19236
rect 50148 19180 50158 19236
rect 51426 19180 51436 19236
rect 51492 19180 53788 19236
rect 53844 19180 53854 19236
rect 54338 19180 54348 19236
rect 54404 19180 55468 19236
rect 55524 19180 56140 19236
rect 56196 19180 56206 19236
rect 12124 19124 12180 19180
rect 8194 19068 8204 19124
rect 8260 19068 10220 19124
rect 10276 19068 10286 19124
rect 11554 19068 11564 19124
rect 11620 19068 11788 19124
rect 11844 19068 11854 19124
rect 12114 19068 12124 19124
rect 12180 19068 12190 19124
rect 23202 19068 23212 19124
rect 23268 19068 23772 19124
rect 23828 19068 23838 19124
rect 24546 19068 24556 19124
rect 24612 19068 25676 19124
rect 25732 19068 25742 19124
rect 29586 19068 29596 19124
rect 29652 19068 30156 19124
rect 30212 19068 31668 19124
rect 42802 19068 42812 19124
rect 42868 19068 44156 19124
rect 44212 19068 44716 19124
rect 44772 19068 44782 19124
rect 47394 19068 47404 19124
rect 47460 19068 49196 19124
rect 49252 19068 49980 19124
rect 50036 19068 50046 19124
rect 52210 19068 52220 19124
rect 52276 19068 52668 19124
rect 52724 19068 53452 19124
rect 53508 19068 53900 19124
rect 53956 19068 55356 19124
rect 55412 19068 55580 19124
rect 55636 19068 55646 19124
rect 31612 19012 31668 19068
rect 6626 18956 6636 19012
rect 6692 18956 8428 19012
rect 8484 18956 11340 19012
rect 11396 18956 11406 19012
rect 12898 18956 12908 19012
rect 12964 18956 13916 19012
rect 13972 18956 14700 19012
rect 14756 18956 15596 19012
rect 15652 18956 15662 19012
rect 26562 18956 26572 19012
rect 26628 18956 27244 19012
rect 27300 18956 27310 19012
rect 29362 18956 29372 19012
rect 29428 18956 30492 19012
rect 30548 18956 30558 19012
rect 30678 18956 30716 19012
rect 30772 18956 30782 19012
rect 31602 18956 31612 19012
rect 31668 18956 31678 19012
rect 39442 18956 39452 19012
rect 39508 18956 40236 19012
rect 40292 18956 40302 19012
rect 46498 18956 46508 19012
rect 46564 18956 47292 19012
rect 47348 18956 47358 19012
rect 50418 18956 50428 19012
rect 50484 18956 51436 19012
rect 51492 18956 51502 19012
rect 30268 18844 33068 18900
rect 33124 18844 34748 18900
rect 34804 18844 34814 18900
rect 40898 18844 40908 18900
rect 40964 18844 41580 18900
rect 41636 18844 41646 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 30268 18788 30324 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 28466 18732 28476 18788
rect 28532 18732 30268 18788
rect 30324 18732 30334 18788
rect 30594 18732 30604 18788
rect 30660 18732 31164 18788
rect 31220 18732 31230 18788
rect 31490 18732 31500 18788
rect 31556 18732 32060 18788
rect 32116 18732 40796 18788
rect 40852 18732 40862 18788
rect 56690 18732 56700 18788
rect 56756 18732 57372 18788
rect 57428 18732 57438 18788
rect 57698 18732 57708 18788
rect 57764 18732 58604 18788
rect 58660 18732 58670 18788
rect 4162 18620 4172 18676
rect 4228 18620 4508 18676
rect 4564 18620 6076 18676
rect 6132 18620 6142 18676
rect 10210 18620 10220 18676
rect 10276 18620 10556 18676
rect 10612 18620 10622 18676
rect 24994 18620 25004 18676
rect 25060 18620 25676 18676
rect 25732 18620 26572 18676
rect 26628 18620 26638 18676
rect 27010 18620 27020 18676
rect 27076 18620 27916 18676
rect 27972 18620 27982 18676
rect 29474 18620 29484 18676
rect 29540 18620 31276 18676
rect 31332 18620 31612 18676
rect 31668 18620 31678 18676
rect 33506 18620 33516 18676
rect 33572 18620 34636 18676
rect 34692 18620 34702 18676
rect 37314 18620 37324 18676
rect 37380 18620 41356 18676
rect 41412 18620 41580 18676
rect 41636 18620 41646 18676
rect 42242 18620 42252 18676
rect 42308 18620 45500 18676
rect 45556 18620 45566 18676
rect 53554 18620 53564 18676
rect 53620 18620 54012 18676
rect 54068 18620 54078 18676
rect 56578 18620 56588 18676
rect 56644 18620 57596 18676
rect 57652 18620 57662 18676
rect 3714 18508 3724 18564
rect 3780 18508 7084 18564
rect 7140 18508 7150 18564
rect 12114 18508 12124 18564
rect 12180 18508 13468 18564
rect 13524 18508 13534 18564
rect 20188 18508 23548 18564
rect 23604 18508 23614 18564
rect 23874 18508 23884 18564
rect 23940 18508 24332 18564
rect 24388 18508 24398 18564
rect 24770 18508 24780 18564
rect 24836 18508 25900 18564
rect 25956 18508 25966 18564
rect 26898 18508 26908 18564
rect 26964 18508 27468 18564
rect 27524 18508 27534 18564
rect 29558 18508 29596 18564
rect 29652 18508 29662 18564
rect 29932 18508 31052 18564
rect 31108 18508 32172 18564
rect 32228 18508 32238 18564
rect 20188 18452 20244 18508
rect 3378 18396 3388 18452
rect 3444 18396 7980 18452
rect 8036 18396 8540 18452
rect 8596 18396 8606 18452
rect 9650 18396 9660 18452
rect 9716 18396 12572 18452
rect 12628 18396 13356 18452
rect 13412 18396 13422 18452
rect 16146 18396 16156 18452
rect 16212 18396 20244 18452
rect 26338 18396 26348 18452
rect 26404 18396 27580 18452
rect 27636 18396 27646 18452
rect 28354 18396 28364 18452
rect 28420 18396 28812 18452
rect 28868 18396 29036 18452
rect 29092 18396 29102 18452
rect 29932 18340 29988 18508
rect 34188 18452 34244 18620
rect 34402 18508 34412 18564
rect 34468 18508 35644 18564
rect 35700 18508 37436 18564
rect 37492 18508 37502 18564
rect 38994 18508 39004 18564
rect 39060 18508 45612 18564
rect 45668 18508 45678 18564
rect 52770 18508 52780 18564
rect 52836 18508 53452 18564
rect 53508 18508 53518 18564
rect 56018 18508 56028 18564
rect 56084 18508 57820 18564
rect 57876 18508 57886 18564
rect 30594 18396 30604 18452
rect 30660 18396 31500 18452
rect 31556 18396 33628 18452
rect 33684 18396 33694 18452
rect 34178 18396 34188 18452
rect 34244 18396 36092 18452
rect 36148 18396 36158 18452
rect 39778 18396 39788 18452
rect 39844 18396 40236 18452
rect 40292 18396 43148 18452
rect 43204 18396 43214 18452
rect 43586 18396 43596 18452
rect 43652 18396 48076 18452
rect 48132 18396 48142 18452
rect 54114 18396 54124 18452
rect 54180 18396 55916 18452
rect 55972 18396 55982 18452
rect 56242 18396 56252 18452
rect 56308 18396 56476 18452
rect 56532 18396 56542 18452
rect 34748 18340 34804 18396
rect 4050 18284 4060 18340
rect 4116 18284 4620 18340
rect 4676 18284 6748 18340
rect 6804 18284 6814 18340
rect 15698 18284 15708 18340
rect 15764 18284 17948 18340
rect 18004 18284 19180 18340
rect 19236 18284 19246 18340
rect 19618 18284 19628 18340
rect 19684 18284 21644 18340
rect 21700 18284 24332 18340
rect 24388 18284 24398 18340
rect 29922 18284 29932 18340
rect 29988 18284 29998 18340
rect 32722 18284 32732 18340
rect 32788 18284 33292 18340
rect 33348 18284 33358 18340
rect 34738 18284 34748 18340
rect 34804 18284 34814 18340
rect 44482 18284 44492 18340
rect 44548 18284 45948 18340
rect 46004 18284 46014 18340
rect 18498 18172 18508 18228
rect 18564 18172 20076 18228
rect 20132 18172 20142 18228
rect 28802 18172 28812 18228
rect 28868 18172 31836 18228
rect 31892 18172 32284 18228
rect 32340 18172 32350 18228
rect 40450 18172 40460 18228
rect 40516 18172 41804 18228
rect 41860 18172 42812 18228
rect 42868 18172 42878 18228
rect 50306 18172 50316 18228
rect 50372 18172 50876 18228
rect 50932 18172 50942 18228
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 36642 17836 36652 17892
rect 36708 17836 37436 17892
rect 37492 17836 37660 17892
rect 37716 17836 37726 17892
rect 48962 17836 48972 17892
rect 49028 17836 52108 17892
rect 52164 17836 52332 17892
rect 52388 17836 52398 17892
rect 2258 17724 2268 17780
rect 2324 17724 4508 17780
rect 4564 17724 4844 17780
rect 4900 17724 6524 17780
rect 6580 17724 7532 17780
rect 7588 17724 7868 17780
rect 7924 17724 8428 17780
rect 8484 17724 8494 17780
rect 19618 17724 19628 17780
rect 19684 17724 20188 17780
rect 20244 17724 20524 17780
rect 20580 17724 20972 17780
rect 21028 17724 21038 17780
rect 38322 17724 38332 17780
rect 38388 17724 38892 17780
rect 38948 17724 39116 17780
rect 39172 17724 39182 17780
rect 41346 17724 41356 17780
rect 41412 17724 42476 17780
rect 42532 17724 42542 17780
rect 43474 17724 43484 17780
rect 43540 17724 43820 17780
rect 43876 17724 43886 17780
rect 44482 17724 44492 17780
rect 44548 17724 46620 17780
rect 46676 17724 47516 17780
rect 47572 17724 47582 17780
rect 48738 17724 48748 17780
rect 48804 17724 49980 17780
rect 50036 17724 50046 17780
rect 19170 17612 19180 17668
rect 19236 17612 19740 17668
rect 19796 17612 22764 17668
rect 22820 17612 22830 17668
rect 23090 17612 23100 17668
rect 23156 17612 25340 17668
rect 25396 17612 25406 17668
rect 25666 17612 25676 17668
rect 25732 17612 27132 17668
rect 27188 17612 27198 17668
rect 31714 17612 31724 17668
rect 31780 17612 32284 17668
rect 32340 17612 32620 17668
rect 32676 17612 32686 17668
rect 33394 17612 33404 17668
rect 33460 17612 33852 17668
rect 33908 17612 34188 17668
rect 34244 17612 34254 17668
rect 34626 17612 34636 17668
rect 34692 17612 35868 17668
rect 35924 17612 35934 17668
rect 43026 17612 43036 17668
rect 43092 17612 43708 17668
rect 43764 17612 43774 17668
rect 47842 17612 47852 17668
rect 47908 17612 48860 17668
rect 48916 17612 48926 17668
rect 26572 17556 26628 17612
rect 19842 17500 19852 17556
rect 19908 17500 20972 17556
rect 21028 17500 21038 17556
rect 26562 17500 26572 17556
rect 26628 17500 26638 17556
rect 30258 17500 30268 17556
rect 30324 17500 30604 17556
rect 30660 17500 30670 17556
rect 30818 17500 30828 17556
rect 30884 17500 32732 17556
rect 32788 17500 33180 17556
rect 33236 17500 33246 17556
rect 35298 17500 35308 17556
rect 35364 17500 35644 17556
rect 35700 17500 35868 17556
rect 35924 17500 36764 17556
rect 36820 17500 37772 17556
rect 37828 17500 37838 17556
rect 42802 17500 42812 17556
rect 42868 17500 44380 17556
rect 44436 17500 44446 17556
rect 48066 17500 48076 17556
rect 48132 17500 48972 17556
rect 49028 17500 49038 17556
rect 16258 17388 16268 17444
rect 16324 17388 18508 17444
rect 18564 17388 18574 17444
rect 20178 17388 20188 17444
rect 20244 17388 21980 17444
rect 22036 17388 22046 17444
rect 28130 17388 28140 17444
rect 28196 17388 28476 17444
rect 28532 17388 28542 17444
rect 31154 17388 31164 17444
rect 31220 17388 31500 17444
rect 31556 17388 31566 17444
rect 35970 17388 35980 17444
rect 36036 17388 37884 17444
rect 37940 17388 37950 17444
rect 40338 17388 40348 17444
rect 40404 17388 40908 17444
rect 40964 17388 40974 17444
rect 21298 17276 21308 17332
rect 21364 17276 21868 17332
rect 21924 17276 22316 17332
rect 22372 17276 22382 17332
rect 28690 17276 28700 17332
rect 28756 17276 29148 17332
rect 29204 17276 44044 17332
rect 44100 17276 44110 17332
rect 53778 17276 53788 17332
rect 53844 17276 57260 17332
rect 57316 17276 57326 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 20300 17164 20860 17220
rect 20916 17164 21420 17220
rect 21476 17164 23548 17220
rect 23604 17164 23614 17220
rect 31826 17164 31836 17220
rect 31892 17164 33964 17220
rect 34020 17164 34030 17220
rect 34850 17164 34860 17220
rect 34916 17164 39004 17220
rect 39060 17164 40348 17220
rect 40404 17164 41468 17220
rect 41524 17164 41534 17220
rect 42130 17164 42140 17220
rect 42196 17164 42588 17220
rect 42644 17164 45668 17220
rect 4610 17052 4620 17108
rect 4676 17052 7644 17108
rect 7700 17052 7710 17108
rect 10210 17052 10220 17108
rect 10276 17052 12012 17108
rect 12068 17052 12078 17108
rect 14914 17052 14924 17108
rect 14980 17052 16828 17108
rect 16884 17052 18060 17108
rect 18116 17052 19180 17108
rect 19236 17052 19246 17108
rect 5292 16884 5348 17052
rect 20300 16996 20356 17164
rect 45612 17108 45668 17164
rect 20514 17052 20524 17108
rect 20580 17052 21644 17108
rect 21700 17052 23212 17108
rect 23268 17052 23278 17108
rect 24994 17052 25004 17108
rect 25060 17052 26348 17108
rect 26404 17052 26414 17108
rect 27010 17052 27020 17108
rect 27076 17052 28364 17108
rect 28420 17052 28430 17108
rect 29362 17052 29372 17108
rect 29428 17052 31164 17108
rect 31220 17052 31230 17108
rect 34066 17052 34076 17108
rect 34132 17052 34524 17108
rect 34580 17052 35084 17108
rect 35140 17052 36092 17108
rect 36148 17052 36158 17108
rect 39554 17052 39564 17108
rect 39620 17052 40572 17108
rect 40628 17052 40638 17108
rect 42914 17052 42924 17108
rect 42980 17052 43260 17108
rect 43316 17052 44268 17108
rect 44324 17052 45164 17108
rect 45220 17052 45230 17108
rect 45602 17052 45612 17108
rect 45668 17052 45948 17108
rect 46004 17052 46284 17108
rect 46340 17052 46350 17108
rect 55412 17052 56476 17108
rect 56532 17052 58380 17108
rect 58436 17052 58446 17108
rect 55412 16996 55468 17052
rect 11228 16940 17052 16996
rect 17108 16940 18844 16996
rect 18900 16940 20356 16996
rect 21074 16940 21084 16996
rect 21140 16940 22204 16996
rect 22260 16940 22270 16996
rect 22978 16940 22988 16996
rect 23044 16940 24108 16996
rect 24164 16940 24444 16996
rect 24500 16940 24510 16996
rect 33170 16940 33180 16996
rect 33236 16940 34188 16996
rect 34244 16940 36540 16996
rect 36596 16940 36606 16996
rect 43138 16940 43148 16996
rect 43204 16940 43484 16996
rect 43540 16940 44716 16996
rect 44772 16940 44782 16996
rect 53890 16940 53900 16996
rect 53956 16940 55468 16996
rect 56354 16940 56364 16996
rect 56420 16940 57036 16996
rect 57092 16940 57102 16996
rect 11228 16884 11284 16940
rect 5282 16828 5292 16884
rect 5348 16828 5358 16884
rect 7746 16828 7756 16884
rect 7812 16828 8540 16884
rect 8596 16828 8606 16884
rect 11218 16828 11228 16884
rect 11284 16828 11294 16884
rect 12226 16828 12236 16884
rect 12292 16828 13916 16884
rect 13972 16828 16268 16884
rect 16324 16828 16334 16884
rect 17938 16828 17948 16884
rect 18004 16828 21868 16884
rect 21924 16828 21934 16884
rect 26002 16828 26012 16884
rect 26068 16828 26684 16884
rect 26740 16828 26750 16884
rect 29026 16828 29036 16884
rect 29092 16828 30212 16884
rect 32946 16828 32956 16884
rect 33012 16828 35532 16884
rect 35588 16828 35756 16884
rect 35812 16828 35822 16884
rect 42690 16828 42700 16884
rect 42756 16828 42924 16884
rect 42980 16828 43820 16884
rect 43876 16828 43886 16884
rect 53666 16828 53676 16884
rect 53732 16828 54012 16884
rect 54068 16828 54078 16884
rect 55010 16828 55020 16884
rect 55076 16828 55580 16884
rect 55636 16828 56028 16884
rect 56084 16828 56094 16884
rect 30156 16772 30212 16828
rect 14018 16716 14028 16772
rect 14084 16716 15148 16772
rect 15204 16716 15214 16772
rect 25666 16716 25676 16772
rect 25732 16716 26124 16772
rect 26180 16716 26190 16772
rect 30156 16716 30380 16772
rect 30436 16716 30446 16772
rect 30594 16716 30604 16772
rect 30660 16716 37548 16772
rect 37604 16716 37614 16772
rect 18610 16604 18620 16660
rect 18676 16604 26908 16660
rect 27346 16604 27356 16660
rect 27412 16604 28476 16660
rect 28532 16604 29036 16660
rect 29092 16604 29102 16660
rect 29698 16604 29708 16660
rect 29764 16604 30660 16660
rect 34178 16604 34188 16660
rect 34244 16604 36204 16660
rect 36260 16604 36270 16660
rect 40674 16604 40684 16660
rect 40740 16604 43708 16660
rect 43764 16604 43774 16660
rect 56802 16604 56812 16660
rect 56868 16604 57596 16660
rect 57652 16604 57662 16660
rect 26852 16548 26908 16604
rect 30604 16548 30660 16604
rect 26852 16492 30380 16548
rect 30436 16492 30446 16548
rect 30594 16492 30604 16548
rect 30660 16492 30670 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 28802 16380 28812 16436
rect 28868 16380 30492 16436
rect 30548 16380 30558 16436
rect 39106 16380 39116 16436
rect 39172 16380 40236 16436
rect 40292 16380 40302 16436
rect 18386 16268 18396 16324
rect 18452 16268 18956 16324
rect 19012 16268 20412 16324
rect 20468 16268 20860 16324
rect 20916 16268 22652 16324
rect 22708 16268 22718 16324
rect 26786 16268 26796 16324
rect 26852 16268 39452 16324
rect 39508 16268 39518 16324
rect 6402 16156 6412 16212
rect 6468 16156 6972 16212
rect 7028 16156 8428 16212
rect 13010 16156 13020 16212
rect 13076 16156 13692 16212
rect 13748 16156 14588 16212
rect 14644 16156 14654 16212
rect 18274 16156 18284 16212
rect 18340 16156 19628 16212
rect 19684 16156 19852 16212
rect 19908 16156 19918 16212
rect 21746 16156 21756 16212
rect 21812 16156 23324 16212
rect 23380 16156 23390 16212
rect 24882 16156 24892 16212
rect 24948 16156 25676 16212
rect 25732 16156 25742 16212
rect 29558 16156 29596 16212
rect 29652 16156 29662 16212
rect 30678 16156 30716 16212
rect 30772 16156 30782 16212
rect 32386 16156 32396 16212
rect 32452 16156 32732 16212
rect 32788 16156 33068 16212
rect 33124 16156 34748 16212
rect 34804 16156 34814 16212
rect 35410 16156 35420 16212
rect 35476 16156 35868 16212
rect 35924 16156 37436 16212
rect 37492 16156 37884 16212
rect 37940 16156 37950 16212
rect 38434 16156 38444 16212
rect 38500 16156 39116 16212
rect 39172 16156 39564 16212
rect 39620 16156 39630 16212
rect 8372 15876 8428 16156
rect 23874 16044 23884 16100
rect 23940 16044 24332 16100
rect 24388 16044 24398 16100
rect 31238 16044 31276 16100
rect 31332 16044 31342 16100
rect 34066 16044 34076 16100
rect 34132 16044 35756 16100
rect 35812 16044 35822 16100
rect 38994 16044 39004 16100
rect 39060 16044 40124 16100
rect 40180 16044 40190 16100
rect 42914 16044 42924 16100
rect 42980 16044 43372 16100
rect 43428 16044 43438 16100
rect 10210 15932 10220 15988
rect 10276 15932 20188 15988
rect 20244 15932 20254 15988
rect 21410 15932 21420 15988
rect 21476 15932 22204 15988
rect 22260 15932 22540 15988
rect 22596 15932 22606 15988
rect 32834 15932 32844 15988
rect 32900 15932 33628 15988
rect 33684 15932 34188 15988
rect 34244 15932 36428 15988
rect 36484 15932 36494 15988
rect 42802 15932 42812 15988
rect 42868 15932 44604 15988
rect 44660 15932 44670 15988
rect 52434 15932 52444 15988
rect 52500 15932 52668 15988
rect 52724 15932 53452 15988
rect 53508 15932 54460 15988
rect 54516 15932 54526 15988
rect 55234 15932 55244 15988
rect 55300 15932 55692 15988
rect 55748 15932 55758 15988
rect 8372 15820 13468 15876
rect 13524 15820 14028 15876
rect 14084 15820 14094 15876
rect 28466 15820 28476 15876
rect 28532 15820 28924 15876
rect 28980 15820 29372 15876
rect 29428 15820 29438 15876
rect 35634 15820 35644 15876
rect 35700 15820 35756 15876
rect 35812 15820 35822 15876
rect 43698 15820 43708 15876
rect 43764 15820 48636 15876
rect 48692 15820 49756 15876
rect 49812 15820 49822 15876
rect 52546 15820 52556 15876
rect 52612 15820 53676 15876
rect 53732 15820 54236 15876
rect 54292 15820 54302 15876
rect 28578 15708 28588 15764
rect 28644 15708 28812 15764
rect 28868 15708 28878 15764
rect 31042 15708 31052 15764
rect 31108 15708 32172 15764
rect 32228 15708 32238 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 27010 15596 27020 15652
rect 27076 15596 27356 15652
rect 27412 15596 27422 15652
rect 24546 15484 24556 15540
rect 24612 15484 25900 15540
rect 25956 15484 25966 15540
rect 26226 15484 26236 15540
rect 26292 15484 26908 15540
rect 26964 15484 26974 15540
rect 31266 15484 31276 15540
rect 31332 15484 31388 15540
rect 31444 15484 31454 15540
rect 35970 15484 35980 15540
rect 36036 15484 36204 15540
rect 36260 15484 36764 15540
rect 36820 15484 38108 15540
rect 38164 15484 38174 15540
rect 56354 15484 56364 15540
rect 56420 15484 58716 15540
rect 58772 15484 58782 15540
rect 15362 15372 15372 15428
rect 15428 15372 16604 15428
rect 16660 15372 17612 15428
rect 17668 15372 17678 15428
rect 24434 15372 24444 15428
rect 24500 15372 24892 15428
rect 24948 15372 27020 15428
rect 27076 15372 27086 15428
rect 32610 15372 32620 15428
rect 32676 15372 32686 15428
rect 34850 15372 34860 15428
rect 34916 15372 35140 15428
rect 35858 15372 35868 15428
rect 35924 15372 37436 15428
rect 37492 15372 37996 15428
rect 38052 15372 38062 15428
rect 39218 15372 39228 15428
rect 39284 15372 40236 15428
rect 40292 15372 41804 15428
rect 41860 15372 42364 15428
rect 42420 15372 43148 15428
rect 43204 15372 43708 15428
rect 43764 15372 43774 15428
rect 45042 15372 45052 15428
rect 45108 15372 45948 15428
rect 46004 15372 46014 15428
rect 49186 15372 49196 15428
rect 49252 15372 49980 15428
rect 50036 15372 50046 15428
rect 57250 15372 57260 15428
rect 57316 15372 57932 15428
rect 57988 15372 57998 15428
rect 32620 15316 32676 15372
rect 35084 15316 35140 15372
rect 7298 15260 7308 15316
rect 7364 15260 8316 15316
rect 8372 15260 11788 15316
rect 11844 15260 15260 15316
rect 15316 15260 18508 15316
rect 18564 15260 18574 15316
rect 21186 15260 21196 15316
rect 21252 15260 22204 15316
rect 22260 15260 22270 15316
rect 22866 15260 22876 15316
rect 22932 15260 23772 15316
rect 23828 15260 23838 15316
rect 24098 15260 24108 15316
rect 24164 15260 25676 15316
rect 25732 15260 27132 15316
rect 27188 15260 27198 15316
rect 28578 15260 28588 15316
rect 28644 15260 29596 15316
rect 29652 15260 29662 15316
rect 31378 15260 31388 15316
rect 31444 15260 32172 15316
rect 32228 15260 33516 15316
rect 33572 15260 33964 15316
rect 34020 15260 34030 15316
rect 35074 15260 35084 15316
rect 35140 15260 35150 15316
rect 36194 15260 36204 15316
rect 36260 15260 37212 15316
rect 37268 15260 38332 15316
rect 38388 15260 38398 15316
rect 39330 15260 39340 15316
rect 39396 15260 39900 15316
rect 39956 15260 39966 15316
rect 40786 15260 40796 15316
rect 40852 15260 42588 15316
rect 42644 15260 43484 15316
rect 43540 15260 43550 15316
rect 49634 15260 49644 15316
rect 49700 15260 52668 15316
rect 52724 15260 52734 15316
rect 54786 15260 54796 15316
rect 54852 15260 55580 15316
rect 55636 15260 55646 15316
rect 56690 15260 56700 15316
rect 56756 15260 57596 15316
rect 57652 15260 57662 15316
rect 6738 15148 6748 15204
rect 6804 15148 8652 15204
rect 8708 15148 9660 15204
rect 9716 15148 9726 15204
rect 9986 15148 9996 15204
rect 10052 15148 11564 15204
rect 11620 15148 11630 15204
rect 47282 15148 47292 15204
rect 47348 15148 48412 15204
rect 48468 15148 49532 15204
rect 49588 15148 49598 15204
rect 6290 15036 6300 15092
rect 6356 15036 18620 15092
rect 18676 15036 18686 15092
rect 24210 15036 24220 15092
rect 24276 15036 27468 15092
rect 27524 15036 28588 15092
rect 28644 15036 28654 15092
rect 29586 15036 29596 15092
rect 29652 15036 30268 15092
rect 30324 15036 30334 15092
rect 30818 15036 30828 15092
rect 30884 15036 31724 15092
rect 31780 15036 31790 15092
rect 32498 15036 32508 15092
rect 32564 15036 35420 15092
rect 35476 15036 35812 15092
rect 35756 14980 35812 15036
rect 38612 15036 43708 15092
rect 35746 14924 35756 14980
rect 35812 14924 35822 14980
rect 36306 14924 36316 14980
rect 36372 14924 37772 14980
rect 37828 14924 37838 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 8754 14700 8764 14756
rect 8820 14700 14140 14756
rect 14196 14700 14206 14756
rect 27906 14700 27916 14756
rect 27972 14700 30156 14756
rect 30212 14700 35308 14756
rect 35364 14700 35644 14756
rect 35700 14700 36764 14756
rect 36820 14700 36830 14756
rect 38612 14644 38668 15036
rect 40450 14924 40460 14980
rect 40516 14924 41356 14980
rect 41412 14924 42700 14980
rect 42756 14924 42766 14980
rect 43652 14868 43708 15036
rect 43652 14812 53564 14868
rect 53620 14812 53630 14868
rect 50866 14700 50876 14756
rect 50932 14700 51884 14756
rect 51940 14700 52332 14756
rect 52388 14700 52398 14756
rect 5618 14588 5628 14644
rect 5684 14588 6412 14644
rect 6468 14588 6860 14644
rect 6916 14588 8092 14644
rect 8148 14588 9548 14644
rect 9604 14588 9614 14644
rect 30482 14588 30492 14644
rect 30548 14588 30716 14644
rect 30772 14588 38668 14644
rect 44706 14588 44716 14644
rect 44772 14588 46508 14644
rect 46564 14588 46956 14644
rect 47012 14588 47022 14644
rect 48738 14588 48748 14644
rect 48804 14588 49644 14644
rect 49700 14588 49710 14644
rect 54674 14588 54684 14644
rect 54740 14588 56476 14644
rect 56532 14588 56542 14644
rect 16034 14476 16044 14532
rect 16100 14476 17948 14532
rect 18004 14476 18014 14532
rect 31490 14476 31500 14532
rect 31556 14476 32284 14532
rect 32340 14476 32732 14532
rect 32788 14476 32798 14532
rect 34514 14476 34524 14532
rect 34580 14476 35084 14532
rect 35140 14476 35308 14532
rect 35252 14420 35308 14476
rect 22978 14364 22988 14420
rect 23044 14364 25564 14420
rect 25620 14364 25630 14420
rect 26114 14364 26124 14420
rect 26180 14364 27244 14420
rect 27300 14364 27310 14420
rect 29474 14364 29484 14420
rect 29540 14364 29932 14420
rect 29988 14364 30380 14420
rect 30436 14364 30446 14420
rect 35252 14364 36316 14420
rect 36372 14364 36382 14420
rect 16034 14252 16044 14308
rect 16100 14252 21644 14308
rect 21700 14252 21710 14308
rect 25890 14252 25900 14308
rect 25956 14252 26796 14308
rect 26852 14252 27356 14308
rect 27412 14252 27422 14308
rect 27234 14140 27244 14196
rect 27300 14140 27692 14196
rect 27748 14140 28812 14196
rect 28868 14140 28878 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 29586 14028 29596 14084
rect 29652 14028 33628 14084
rect 33684 14028 34300 14084
rect 34356 14028 34366 14084
rect 40002 14028 40012 14084
rect 40068 14028 45724 14084
rect 45780 14028 46060 14084
rect 46116 14028 46620 14084
rect 46676 14028 47740 14084
rect 47796 14028 48188 14084
rect 48244 14028 48254 14084
rect 31490 13916 31500 13972
rect 31556 13916 32508 13972
rect 32564 13916 32574 13972
rect 39778 13916 39788 13972
rect 39844 13916 40124 13972
rect 40180 13916 41132 13972
rect 41188 13916 41198 13972
rect 56578 13916 56588 13972
rect 56644 13916 57820 13972
rect 57876 13916 57886 13972
rect 26450 13804 26460 13860
rect 26516 13804 27580 13860
rect 27636 13804 27646 13860
rect 30818 13804 30828 13860
rect 30884 13804 31164 13860
rect 31220 13804 31556 13860
rect 33954 13804 33964 13860
rect 34020 13804 34636 13860
rect 34692 13804 35420 13860
rect 35476 13804 35486 13860
rect 38322 13804 38332 13860
rect 38388 13804 39564 13860
rect 39620 13804 39630 13860
rect 43026 13804 43036 13860
rect 43092 13804 43708 13860
rect 43764 13804 44156 13860
rect 44212 13804 44222 13860
rect 52322 13804 52332 13860
rect 52388 13804 53788 13860
rect 53844 13804 53854 13860
rect 31500 13748 31556 13804
rect 10098 13692 10108 13748
rect 10164 13692 10556 13748
rect 10612 13692 10892 13748
rect 10948 13692 10958 13748
rect 11218 13692 11228 13748
rect 11284 13692 16268 13748
rect 16324 13692 24780 13748
rect 24836 13692 24846 13748
rect 26338 13692 26348 13748
rect 26404 13692 27692 13748
rect 27748 13692 31164 13748
rect 31220 13692 31230 13748
rect 31490 13692 31500 13748
rect 31556 13692 31566 13748
rect 32386 13692 32396 13748
rect 32452 13692 33740 13748
rect 33796 13692 33806 13748
rect 32834 13580 32844 13636
rect 32900 13580 33852 13636
rect 33908 13580 34076 13636
rect 34132 13580 34636 13636
rect 34692 13580 34702 13636
rect 38210 13580 38220 13636
rect 38276 13580 45612 13636
rect 45668 13580 45948 13636
rect 46004 13580 46396 13636
rect 46452 13580 46844 13636
rect 46900 13580 47628 13636
rect 47684 13580 47694 13636
rect 14242 13468 14252 13524
rect 14308 13468 24220 13524
rect 24276 13468 24286 13524
rect 24882 13468 24892 13524
rect 24948 13468 25452 13524
rect 25508 13468 26124 13524
rect 26180 13468 26348 13524
rect 26404 13468 26414 13524
rect 28018 13468 28028 13524
rect 28084 13468 31724 13524
rect 31780 13468 32396 13524
rect 32452 13468 32620 13524
rect 32676 13468 32956 13524
rect 33012 13468 33022 13524
rect 54786 13468 54796 13524
rect 54852 13468 55468 13524
rect 55524 13468 55534 13524
rect 10098 13356 10108 13412
rect 10164 13356 11116 13412
rect 11172 13356 11900 13412
rect 11956 13356 11966 13412
rect 18274 13356 18284 13412
rect 18340 13356 19180 13412
rect 19236 13356 19246 13412
rect 37762 13356 37772 13412
rect 37828 13356 38892 13412
rect 38948 13356 40796 13412
rect 40852 13356 41244 13412
rect 41300 13356 41468 13412
rect 41524 13356 41534 13412
rect 42018 13356 42028 13412
rect 42084 13356 42252 13412
rect 42308 13356 43260 13412
rect 43316 13356 43326 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 11330 13132 11340 13188
rect 11396 13132 17500 13188
rect 17556 13132 17566 13188
rect 19058 13132 19068 13188
rect 19124 13132 23436 13188
rect 23492 13132 23502 13188
rect 26674 13132 26684 13188
rect 26740 13132 26750 13188
rect 26684 13076 26740 13132
rect 4274 13020 4284 13076
rect 4340 13020 5740 13076
rect 5796 13020 5806 13076
rect 13682 13020 13692 13076
rect 13748 13020 13916 13076
rect 13972 13020 14588 13076
rect 14644 13020 14654 13076
rect 18722 13020 18732 13076
rect 18788 13020 19628 13076
rect 19684 13020 20188 13076
rect 20244 13020 20254 13076
rect 26450 13020 26460 13076
rect 26516 13020 26740 13076
rect 39666 13020 39676 13076
rect 39732 13020 46060 13076
rect 46116 13020 46126 13076
rect 47282 13020 47292 13076
rect 47348 13020 49308 13076
rect 49364 13020 49374 13076
rect 51202 13020 51212 13076
rect 51268 13020 52108 13076
rect 52164 13020 52174 13076
rect 18732 12964 18788 13020
rect 8082 12908 8092 12964
rect 8148 12908 8764 12964
rect 8820 12908 8830 12964
rect 10434 12908 10444 12964
rect 10500 12908 11116 12964
rect 11172 12908 11340 12964
rect 11396 12908 11406 12964
rect 11890 12908 11900 12964
rect 11956 12908 12460 12964
rect 12516 12908 12908 12964
rect 12964 12908 18788 12964
rect 19282 12908 19292 12964
rect 19348 12908 19740 12964
rect 19796 12908 20524 12964
rect 20580 12908 20590 12964
rect 29026 12908 29036 12964
rect 29092 12908 29820 12964
rect 29876 12908 29886 12964
rect 39778 12908 39788 12964
rect 39844 12908 41244 12964
rect 41300 12908 41310 12964
rect 50306 12908 50316 12964
rect 50372 12908 50988 12964
rect 51044 12908 51054 12964
rect 3490 12796 3500 12852
rect 3556 12796 4284 12852
rect 4340 12796 9884 12852
rect 9940 12796 9950 12852
rect 23174 12796 23212 12852
rect 23268 12796 24780 12852
rect 24836 12796 24846 12852
rect 30146 12796 30156 12852
rect 30212 12796 30716 12852
rect 30772 12796 30782 12852
rect 49634 12796 49644 12852
rect 49700 12796 50764 12852
rect 50820 12796 50830 12852
rect 8754 12684 8764 12740
rect 8820 12684 10108 12740
rect 10164 12684 10174 12740
rect 14130 12684 14140 12740
rect 14196 12684 14924 12740
rect 14980 12684 15372 12740
rect 15428 12684 15438 12740
rect 28354 12684 28364 12740
rect 28420 12684 30044 12740
rect 30100 12684 30110 12740
rect 37314 12684 37324 12740
rect 37380 12684 38556 12740
rect 38612 12684 39452 12740
rect 39508 12684 39518 12740
rect 50194 12684 50204 12740
rect 50260 12684 51324 12740
rect 51380 12684 51390 12740
rect 22642 12572 22652 12628
rect 22708 12572 23324 12628
rect 23380 12572 23390 12628
rect 28578 12572 28588 12628
rect 28644 12572 28812 12628
rect 28868 12572 29484 12628
rect 29540 12572 29550 12628
rect 32946 12572 32956 12628
rect 33012 12572 33516 12628
rect 33572 12572 33582 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 6178 12348 6188 12404
rect 6244 12348 8092 12404
rect 8148 12348 8158 12404
rect 17042 12348 17052 12404
rect 17108 12348 24220 12404
rect 24276 12348 24286 12404
rect 30492 12348 30940 12404
rect 30996 12348 31006 12404
rect 35410 12348 35420 12404
rect 35476 12348 35644 12404
rect 35700 12348 35710 12404
rect 41570 12348 41580 12404
rect 41636 12348 42028 12404
rect 42084 12348 42094 12404
rect 43586 12348 43596 12404
rect 43652 12348 43932 12404
rect 43988 12348 43998 12404
rect 47618 12348 47628 12404
rect 47684 12348 49756 12404
rect 49812 12348 49822 12404
rect 30492 12292 30548 12348
rect 16034 12236 16044 12292
rect 16100 12236 21420 12292
rect 21476 12236 21486 12292
rect 22866 12236 22876 12292
rect 22932 12236 23660 12292
rect 23716 12236 24332 12292
rect 24388 12236 24398 12292
rect 30146 12236 30156 12292
rect 30212 12236 30492 12292
rect 30548 12236 30558 12292
rect 34962 12236 34972 12292
rect 35028 12236 35532 12292
rect 35588 12236 35868 12292
rect 35924 12236 36988 12292
rect 37044 12236 37054 12292
rect 39442 12236 39452 12292
rect 39508 12236 40236 12292
rect 40292 12236 40302 12292
rect 40562 12236 40572 12292
rect 40628 12236 41804 12292
rect 41860 12236 42588 12292
rect 42644 12236 42654 12292
rect 56018 12236 56028 12292
rect 56084 12236 56924 12292
rect 56980 12236 57596 12292
rect 57652 12236 57662 12292
rect 3602 12124 3612 12180
rect 3668 12124 4172 12180
rect 4228 12124 4508 12180
rect 4564 12124 5404 12180
rect 5460 12124 5470 12180
rect 6962 12124 6972 12180
rect 7028 12124 8428 12180
rect 8484 12124 8494 12180
rect 20132 12124 31052 12180
rect 31108 12124 31118 12180
rect 34626 12124 34636 12180
rect 34692 12124 35644 12180
rect 35700 12124 36652 12180
rect 36708 12124 37548 12180
rect 37604 12124 37614 12180
rect 55570 12124 55580 12180
rect 55636 12124 57708 12180
rect 57764 12124 57774 12180
rect 19170 12012 19180 12068
rect 19236 12012 19628 12068
rect 19684 12012 19694 12068
rect 16482 11900 16492 11956
rect 16548 11900 18284 11956
rect 18340 11900 18350 11956
rect 20132 11844 20188 12124
rect 27570 12012 27580 12068
rect 27636 12012 28588 12068
rect 28644 12012 30380 12068
rect 30436 12012 30446 12068
rect 36866 11900 36876 11956
rect 36932 11900 37884 11956
rect 37940 11900 38332 11956
rect 38388 11900 39228 11956
rect 39284 11900 40348 11956
rect 40404 11900 41132 11956
rect 41188 11900 42252 11956
rect 42308 11900 42318 11956
rect 57138 11900 57148 11956
rect 57204 11900 58492 11956
rect 58548 11900 58558 11956
rect 16828 11788 20188 11844
rect 23436 11788 27132 11844
rect 27188 11788 27198 11844
rect 40450 11788 40460 11844
rect 40516 11788 40796 11844
rect 40852 11788 41580 11844
rect 41636 11788 41646 11844
rect 55412 11788 56140 11844
rect 56196 11788 56206 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 16828 11732 16884 11788
rect 13122 11676 13132 11732
rect 13188 11676 16884 11732
rect 23436 11620 23492 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 38770 11676 38780 11732
rect 38836 11676 39340 11732
rect 39396 11676 40012 11732
rect 40068 11676 42364 11732
rect 42420 11676 42812 11732
rect 42868 11676 43596 11732
rect 43652 11676 43662 11732
rect 55346 11676 55356 11732
rect 55412 11676 55468 11788
rect 43596 11620 43652 11676
rect 18498 11564 18508 11620
rect 18564 11564 23492 11620
rect 30594 11564 30604 11620
rect 30660 11564 31276 11620
rect 31332 11564 31342 11620
rect 43596 11564 43932 11620
rect 43988 11564 43998 11620
rect 19058 11452 19068 11508
rect 19124 11452 21644 11508
rect 21700 11452 22652 11508
rect 22708 11452 23212 11508
rect 23268 11452 23278 11508
rect 28354 11452 28364 11508
rect 28420 11452 30268 11508
rect 30324 11452 30828 11508
rect 30884 11452 30894 11508
rect 43474 11452 43484 11508
rect 43540 11452 44044 11508
rect 44100 11452 45164 11508
rect 45220 11452 45500 11508
rect 45556 11452 45566 11508
rect 4834 11340 4844 11396
rect 4900 11340 6636 11396
rect 6692 11340 6702 11396
rect 10322 11340 10332 11396
rect 10388 11340 11116 11396
rect 11172 11340 12908 11396
rect 12964 11340 12974 11396
rect 25330 11340 25340 11396
rect 25396 11340 26124 11396
rect 26180 11340 26190 11396
rect 30482 11340 30492 11396
rect 30548 11340 31388 11396
rect 31444 11340 31454 11396
rect 34178 11340 34188 11396
rect 34244 11340 34748 11396
rect 34804 11340 34814 11396
rect 40562 11340 40572 11396
rect 40628 11340 40638 11396
rect 44594 11340 44604 11396
rect 44660 11340 45724 11396
rect 45780 11340 45790 11396
rect 40572 11284 40628 11340
rect 31042 11228 31052 11284
rect 31108 11228 31500 11284
rect 31556 11228 32172 11284
rect 32228 11228 32238 11284
rect 40572 11228 41020 11284
rect 41076 11228 41086 11284
rect 45826 11228 45836 11284
rect 45892 11228 47068 11284
rect 47124 11228 47134 11284
rect 51650 11228 51660 11284
rect 51716 11228 53116 11284
rect 53172 11228 53676 11284
rect 53732 11228 53742 11284
rect 54674 11228 54684 11284
rect 54740 11228 56252 11284
rect 56308 11228 56588 11284
rect 56644 11228 56654 11284
rect 53676 11172 53732 11228
rect 5058 11116 5068 11172
rect 5124 11116 8540 11172
rect 8596 11116 8606 11172
rect 24444 11116 24780 11172
rect 24836 11116 25900 11172
rect 25956 11116 27244 11172
rect 27300 11116 28028 11172
rect 28084 11116 28094 11172
rect 28914 11116 28924 11172
rect 28980 11116 29932 11172
rect 29988 11116 33628 11172
rect 33684 11116 33694 11172
rect 42914 11116 42924 11172
rect 42980 11116 43708 11172
rect 43764 11116 43774 11172
rect 46722 11116 46732 11172
rect 46788 11116 49532 11172
rect 49588 11116 49598 11172
rect 53676 11116 54796 11172
rect 54852 11116 54862 11172
rect 56018 11116 56028 11172
rect 56084 11116 56364 11172
rect 56420 11116 57708 11172
rect 57764 11116 57774 11172
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 24444 10948 24500 11116
rect 43708 11060 43764 11116
rect 26002 11004 26012 11060
rect 26068 11004 26348 11060
rect 26404 11004 27804 11060
rect 27860 11004 27870 11060
rect 33730 11004 33740 11060
rect 33796 11004 34188 11060
rect 34244 11004 34254 11060
rect 43708 11004 46844 11060
rect 46900 11004 46910 11060
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 24434 10892 24444 10948
rect 24500 10892 24510 10948
rect 25890 10780 25900 10836
rect 25956 10780 26460 10836
rect 26516 10780 26526 10836
rect 32386 10780 32396 10836
rect 32452 10780 32956 10836
rect 33012 10780 33022 10836
rect 40114 10780 40124 10836
rect 40180 10780 40684 10836
rect 40740 10780 40750 10836
rect 48738 10780 48748 10836
rect 48804 10780 49196 10836
rect 49252 10780 49756 10836
rect 49812 10780 49822 10836
rect 9650 10668 9660 10724
rect 9716 10668 10332 10724
rect 10388 10668 10398 10724
rect 15922 10668 15932 10724
rect 15988 10668 19628 10724
rect 19684 10668 19694 10724
rect 23538 10668 23548 10724
rect 23604 10668 23772 10724
rect 23828 10668 23838 10724
rect 26114 10668 26124 10724
rect 26180 10668 27132 10724
rect 27188 10668 27198 10724
rect 32162 10668 32172 10724
rect 32228 10668 32620 10724
rect 32676 10668 32686 10724
rect 34290 10668 34300 10724
rect 34356 10668 35420 10724
rect 35476 10668 35486 10724
rect 13570 10556 13580 10612
rect 13636 10556 14140 10612
rect 14196 10556 17612 10612
rect 17668 10556 17678 10612
rect 19954 10556 19964 10612
rect 20020 10556 20524 10612
rect 20580 10556 20590 10612
rect 21186 10556 21196 10612
rect 21252 10556 22092 10612
rect 22148 10556 22158 10612
rect 22642 10556 22652 10612
rect 22708 10556 23660 10612
rect 23716 10556 23726 10612
rect 31490 10556 31500 10612
rect 31556 10556 32508 10612
rect 32564 10556 32574 10612
rect 33506 10556 33516 10612
rect 33572 10556 35308 10612
rect 35364 10556 36540 10612
rect 36596 10556 36606 10612
rect 14018 10444 14028 10500
rect 14084 10444 18508 10500
rect 18564 10444 18574 10500
rect 21410 10444 21420 10500
rect 21476 10444 21980 10500
rect 22036 10444 22540 10500
rect 22596 10444 22606 10500
rect 22978 10444 22988 10500
rect 23044 10444 24332 10500
rect 24388 10444 24398 10500
rect 53330 10444 53340 10500
rect 53396 10444 53900 10500
rect 53956 10444 54572 10500
rect 54628 10444 54638 10500
rect 20132 10332 30156 10388
rect 30212 10332 30222 10388
rect 49858 10332 49868 10388
rect 49924 10332 51660 10388
rect 51716 10332 54124 10388
rect 54180 10332 54460 10388
rect 54516 10332 54526 10388
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 20132 10164 20188 10332
rect 54002 10220 54012 10276
rect 54068 10220 54796 10276
rect 54852 10220 54862 10276
rect 55412 10220 56364 10276
rect 56420 10220 56430 10276
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 55412 10164 55468 10220
rect 16828 10108 20188 10164
rect 36306 10108 36316 10164
rect 36372 10108 37100 10164
rect 37156 10108 37166 10164
rect 48514 10108 48524 10164
rect 48580 10108 49532 10164
rect 49588 10108 49598 10164
rect 55122 10108 55132 10164
rect 55188 10108 55468 10164
rect 16828 10052 16884 10108
rect 13010 9996 13020 10052
rect 13076 9996 16884 10052
rect 26674 9996 26684 10052
rect 26740 9996 27020 10052
rect 27076 9996 27086 10052
rect 38098 9996 38108 10052
rect 38164 9996 38892 10052
rect 38948 9996 38958 10052
rect 39330 9996 39340 10052
rect 39396 9996 40348 10052
rect 40404 9996 41916 10052
rect 41972 9996 41982 10052
rect 44258 9996 44268 10052
rect 44324 9996 45612 10052
rect 45668 9996 45678 10052
rect 55458 9996 55468 10052
rect 55524 9996 55804 10052
rect 55860 9996 56924 10052
rect 56980 9996 56990 10052
rect 24994 9884 25004 9940
rect 25060 9884 28588 9940
rect 28644 9884 29596 9940
rect 29652 9884 29662 9940
rect 33506 9884 33516 9940
rect 33572 9884 34076 9940
rect 34132 9884 34636 9940
rect 34692 9884 35084 9940
rect 35140 9884 35150 9940
rect 37426 9884 37436 9940
rect 37492 9884 37884 9940
rect 37940 9884 38556 9940
rect 38612 9884 40460 9940
rect 40516 9884 40526 9940
rect 48290 9884 48300 9940
rect 48356 9884 49196 9940
rect 49252 9884 49262 9940
rect 9874 9772 9884 9828
rect 9940 9772 13132 9828
rect 13188 9772 13198 9828
rect 25778 9772 25788 9828
rect 25844 9772 26908 9828
rect 26964 9772 26974 9828
rect 31378 9772 31388 9828
rect 31444 9772 32172 9828
rect 32228 9772 32238 9828
rect 34402 9772 34412 9828
rect 34468 9772 35308 9828
rect 35364 9772 37996 9828
rect 38052 9772 38062 9828
rect 40002 9772 40012 9828
rect 40068 9772 40908 9828
rect 40964 9772 40974 9828
rect 43026 9772 43036 9828
rect 43092 9772 44604 9828
rect 44660 9772 45164 9828
rect 45220 9772 47068 9828
rect 47124 9772 47134 9828
rect 51538 9772 51548 9828
rect 51604 9772 52108 9828
rect 52164 9772 52780 9828
rect 52836 9772 52846 9828
rect 56018 9772 56028 9828
rect 56084 9772 58044 9828
rect 58100 9772 58110 9828
rect 4946 9660 4956 9716
rect 5012 9660 5740 9716
rect 5796 9660 5806 9716
rect 18946 9660 18956 9716
rect 19012 9660 23548 9716
rect 23604 9660 23614 9716
rect 27122 9660 27132 9716
rect 27188 9660 27692 9716
rect 27748 9660 28476 9716
rect 28532 9660 28542 9716
rect 34962 9660 34972 9716
rect 35028 9660 37548 9716
rect 37604 9660 37614 9716
rect 40674 9660 40684 9716
rect 40740 9660 41692 9716
rect 41748 9660 41758 9716
rect 43250 9660 43260 9716
rect 43316 9660 44268 9716
rect 44324 9660 44334 9716
rect 49858 9660 49868 9716
rect 49924 9660 50428 9716
rect 50484 9660 50494 9716
rect 12450 9548 12460 9604
rect 12516 9548 13916 9604
rect 13972 9548 13982 9604
rect 18386 9548 18396 9604
rect 18452 9548 18732 9604
rect 18788 9548 19292 9604
rect 19348 9548 19358 9604
rect 26898 9548 26908 9604
rect 26964 9548 27468 9604
rect 27524 9548 27916 9604
rect 27972 9548 28700 9604
rect 28756 9548 28766 9604
rect 29698 9548 29708 9604
rect 29764 9548 30268 9604
rect 30324 9548 30716 9604
rect 30772 9548 30782 9604
rect 32834 9548 32844 9604
rect 32900 9548 43036 9604
rect 43092 9548 43102 9604
rect 43652 9548 44156 9604
rect 44212 9548 45388 9604
rect 45444 9548 45454 9604
rect 50866 9548 50876 9604
rect 50932 9548 51548 9604
rect 51604 9548 54572 9604
rect 54628 9548 54638 9604
rect 43652 9492 43708 9548
rect 42018 9436 42028 9492
rect 42084 9436 43708 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 25788 9324 35644 9380
rect 35700 9324 36204 9380
rect 36260 9324 36270 9380
rect 42242 9324 42252 9380
rect 42308 9324 43148 9380
rect 43204 9324 43214 9380
rect 25788 9268 25844 9324
rect 4834 9212 4844 9268
rect 4900 9212 8428 9268
rect 8484 9212 8494 9268
rect 21298 9212 21308 9268
rect 21364 9212 21868 9268
rect 21924 9212 23100 9268
rect 23156 9212 23548 9268
rect 23604 9212 24668 9268
rect 24724 9212 25116 9268
rect 25172 9212 25182 9268
rect 25666 9212 25676 9268
rect 25732 9212 25788 9268
rect 25844 9212 25854 9268
rect 34850 9212 34860 9268
rect 34916 9212 43260 9268
rect 43316 9212 43326 9268
rect 54674 9212 54684 9268
rect 54740 9212 55692 9268
rect 55748 9212 55758 9268
rect 4844 9044 4900 9212
rect 7634 9100 7644 9156
rect 7700 9100 8316 9156
rect 8372 9100 11004 9156
rect 11060 9100 11070 9156
rect 31602 9100 31612 9156
rect 31668 9100 31678 9156
rect 41906 9100 41916 9156
rect 41972 9100 42588 9156
rect 42644 9100 42654 9156
rect 43698 9100 43708 9156
rect 43764 9100 44156 9156
rect 44212 9100 44716 9156
rect 44772 9100 44782 9156
rect 44930 9100 44940 9156
rect 44996 9100 46508 9156
rect 46564 9100 46574 9156
rect 46946 9100 46956 9156
rect 47012 9100 47404 9156
rect 47460 9100 47470 9156
rect 47618 9100 47628 9156
rect 47684 9100 49084 9156
rect 49140 9100 49756 9156
rect 49812 9100 49822 9156
rect 50418 9100 50428 9156
rect 50484 9100 51660 9156
rect 51716 9100 51726 9156
rect 53666 9100 53676 9156
rect 53732 9100 54348 9156
rect 54404 9100 54414 9156
rect 55346 9100 55356 9156
rect 55412 9100 55916 9156
rect 55972 9100 55982 9156
rect 4274 8988 4284 9044
rect 4340 8988 4900 9044
rect 9538 8988 9548 9044
rect 9604 8988 10556 9044
rect 10612 8988 13580 9044
rect 13636 8988 13646 9044
rect 15026 8988 15036 9044
rect 15092 8988 15484 9044
rect 15540 8988 17052 9044
rect 17108 8988 17612 9044
rect 17668 8988 17678 9044
rect 27570 8988 27580 9044
rect 27636 8988 29932 9044
rect 29988 8988 29998 9044
rect 31612 8932 31668 9100
rect 37874 8988 37884 9044
rect 37940 8988 38780 9044
rect 38836 8988 38846 9044
rect 40450 8988 40460 9044
rect 40516 8988 42028 9044
rect 42084 8988 42094 9044
rect 46610 8988 46620 9044
rect 46676 8988 47180 9044
rect 47236 8988 47246 9044
rect 50642 8988 50652 9044
rect 50708 8988 51548 9044
rect 51604 8988 51614 9044
rect 53554 8988 53564 9044
rect 53620 8988 54236 9044
rect 54292 8988 54302 9044
rect 13346 8876 13356 8932
rect 13412 8876 29148 8932
rect 29204 8876 30940 8932
rect 30996 8876 31668 8932
rect 21970 8764 21980 8820
rect 22036 8764 22652 8820
rect 22708 8764 23436 8820
rect 23492 8764 28140 8820
rect 28196 8764 28206 8820
rect 51090 8764 51100 8820
rect 51156 8764 53004 8820
rect 53060 8764 53070 8820
rect 8978 8652 8988 8708
rect 9044 8652 9772 8708
rect 9828 8652 9838 8708
rect 16482 8652 16492 8708
rect 16548 8652 18620 8708
rect 18676 8652 32396 8708
rect 32452 8652 32462 8708
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 17938 8540 17948 8596
rect 18004 8540 18732 8596
rect 18788 8540 18798 8596
rect 17602 8428 17612 8484
rect 17668 8428 19124 8484
rect 28578 8428 28588 8484
rect 28644 8428 29036 8484
rect 29092 8428 29932 8484
rect 29988 8428 33292 8484
rect 33348 8428 33358 8484
rect 35970 8428 35980 8484
rect 36036 8428 37324 8484
rect 37380 8428 38108 8484
rect 38164 8428 38174 8484
rect 19068 8372 19124 8428
rect 5282 8316 5292 8372
rect 5348 8316 6748 8372
rect 6804 8316 7756 8372
rect 7812 8316 7822 8372
rect 19058 8316 19068 8372
rect 19124 8316 19134 8372
rect 20132 8316 26012 8372
rect 26068 8316 26078 8372
rect 28466 8316 28476 8372
rect 28532 8316 29708 8372
rect 29764 8316 29774 8372
rect 30258 8316 30268 8372
rect 30324 8316 31164 8372
rect 31220 8316 31230 8372
rect 33618 8316 33628 8372
rect 33684 8316 34076 8372
rect 34132 8316 34972 8372
rect 35028 8316 35308 8372
rect 35364 8316 35374 8372
rect 43138 8316 43148 8372
rect 43204 8316 43932 8372
rect 43988 8316 43998 8372
rect 47058 8316 47068 8372
rect 47124 8316 47740 8372
rect 47796 8316 47806 8372
rect 51874 8316 51884 8372
rect 51940 8316 53228 8372
rect 53284 8316 53452 8372
rect 53508 8316 53518 8372
rect 20132 8260 20188 8316
rect 18610 8204 18620 8260
rect 18676 8204 20188 8260
rect 23314 8204 23324 8260
rect 23380 8204 23884 8260
rect 23940 8204 23950 8260
rect 33730 8204 33740 8260
rect 33796 8204 34300 8260
rect 34356 8204 35532 8260
rect 35588 8204 35980 8260
rect 36036 8204 36046 8260
rect 39778 8204 39788 8260
rect 39844 8204 40124 8260
rect 40180 8204 40796 8260
rect 40852 8204 40862 8260
rect 42018 8204 42028 8260
rect 42084 8204 42700 8260
rect 42756 8204 43036 8260
rect 43092 8204 43102 8260
rect 50866 8204 50876 8260
rect 50932 8204 50942 8260
rect 52658 8204 52668 8260
rect 52724 8204 54684 8260
rect 54740 8204 54750 8260
rect 50876 8148 50932 8204
rect 20626 8092 20636 8148
rect 20692 8092 23996 8148
rect 24052 8092 24062 8148
rect 28802 8092 28812 8148
rect 28868 8092 36316 8148
rect 36372 8092 36382 8148
rect 50876 8092 53116 8148
rect 53172 8092 53676 8148
rect 53732 8092 53742 8148
rect 7186 7980 7196 8036
rect 7252 7980 7980 8036
rect 8036 7980 8046 8036
rect 15698 7980 15708 8036
rect 15764 7980 21644 8036
rect 21700 7980 21710 8036
rect 24882 7980 24892 8036
rect 24948 7980 25676 8036
rect 25732 7980 27244 8036
rect 27300 7980 27310 8036
rect 28914 7980 28924 8036
rect 28980 7980 29708 8036
rect 29764 7980 30492 8036
rect 30548 7980 32844 8036
rect 32900 7980 32910 8036
rect 39890 7980 39900 8036
rect 39956 7980 40572 8036
rect 40628 7980 40638 8036
rect 49746 7980 49756 8036
rect 49812 7980 50652 8036
rect 50708 7980 50876 8036
rect 50932 7980 50942 8036
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 27122 7756 27132 7812
rect 27188 7756 27748 7812
rect 27692 7700 27748 7756
rect 13346 7644 13356 7700
rect 13412 7644 13804 7700
rect 13860 7644 13870 7700
rect 22988 7644 23324 7700
rect 23380 7644 23390 7700
rect 26674 7644 26684 7700
rect 26740 7644 27468 7700
rect 27524 7644 27534 7700
rect 27682 7644 27692 7700
rect 27748 7644 29820 7700
rect 29876 7644 30268 7700
rect 30324 7644 30334 7700
rect 43922 7644 43932 7700
rect 43988 7644 44492 7700
rect 44548 7644 44558 7700
rect 49634 7644 49644 7700
rect 49700 7644 57708 7700
rect 57764 7644 57774 7700
rect 22988 7588 23044 7644
rect 20132 7532 20860 7588
rect 20916 7532 22988 7588
rect 23044 7532 23054 7588
rect 24658 7532 24668 7588
rect 24724 7532 25788 7588
rect 25844 7532 25854 7588
rect 27346 7532 27356 7588
rect 27412 7532 28252 7588
rect 28308 7532 28318 7588
rect 20132 7476 20188 7532
rect 19618 7420 19628 7476
rect 19684 7420 20188 7476
rect 22194 7420 22204 7476
rect 22260 7420 22540 7476
rect 22596 7420 24444 7476
rect 24500 7420 24510 7476
rect 30370 7420 30380 7476
rect 30436 7420 31612 7476
rect 31668 7420 32620 7476
rect 32676 7420 32686 7476
rect 38546 7420 38556 7476
rect 38612 7420 39900 7476
rect 39956 7420 41020 7476
rect 41076 7420 41086 7476
rect 43138 7420 43148 7476
rect 43204 7420 43820 7476
rect 43876 7420 43886 7476
rect 30258 7308 30268 7364
rect 30324 7308 31276 7364
rect 31332 7308 31836 7364
rect 31892 7308 31902 7364
rect 8306 7196 8316 7252
rect 8372 7196 8540 7252
rect 8596 7196 13356 7252
rect 13412 7196 13422 7252
rect 26786 7196 26796 7252
rect 26852 7196 28812 7252
rect 28868 7196 30156 7252
rect 30212 7196 31164 7252
rect 31220 7196 31230 7252
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 18722 6860 18732 6916
rect 18788 6860 19628 6916
rect 19684 6860 19694 6916
rect 7634 6636 7644 6692
rect 7700 6636 8316 6692
rect 8372 6636 8382 6692
rect 8866 6636 8876 6692
rect 8932 6636 9548 6692
rect 9604 6636 9614 6692
rect 9986 6636 9996 6692
rect 10052 6636 14476 6692
rect 14532 6636 14542 6692
rect 21746 6636 21756 6692
rect 21812 6636 22540 6692
rect 22596 6636 22606 6692
rect 23090 6636 23100 6692
rect 23156 6636 24668 6692
rect 24724 6636 25788 6692
rect 25844 6636 25854 6692
rect 28018 6636 28028 6692
rect 28084 6636 28588 6692
rect 28644 6636 28654 6692
rect 32946 6636 32956 6692
rect 33012 6636 34188 6692
rect 34244 6636 34860 6692
rect 34916 6636 35084 6692
rect 35140 6636 35980 6692
rect 36036 6636 36046 6692
rect 4834 6524 4844 6580
rect 4900 6524 5628 6580
rect 5684 6524 7196 6580
rect 7252 6524 7262 6580
rect 8876 6468 8932 6636
rect 15362 6524 15372 6580
rect 15428 6524 20300 6580
rect 20356 6524 20366 6580
rect 21970 6524 21980 6580
rect 22036 6524 24780 6580
rect 24836 6524 24846 6580
rect 27010 6524 27020 6580
rect 27076 6524 27580 6580
rect 27636 6524 29596 6580
rect 29652 6524 29932 6580
rect 29988 6524 29998 6580
rect 53778 6524 53788 6580
rect 53844 6524 56700 6580
rect 56756 6524 56766 6580
rect 55468 6468 55524 6524
rect 5506 6412 5516 6468
rect 5572 6412 7980 6468
rect 8036 6412 8932 6468
rect 18162 6412 18172 6468
rect 18228 6412 19404 6468
rect 19460 6412 19470 6468
rect 22978 6412 22988 6468
rect 23044 6412 23436 6468
rect 23492 6412 24220 6468
rect 24276 6412 24286 6468
rect 25442 6412 25452 6468
rect 25508 6412 26348 6468
rect 26404 6412 26414 6468
rect 33058 6412 33068 6468
rect 33124 6412 33740 6468
rect 33796 6412 33806 6468
rect 48626 6412 48636 6468
rect 48692 6412 55020 6468
rect 55076 6412 55086 6468
rect 55458 6412 55468 6468
rect 55524 6412 55534 6468
rect 22530 6300 22540 6356
rect 22596 6300 23212 6356
rect 23268 6300 23548 6356
rect 23604 6300 23996 6356
rect 24052 6300 24062 6356
rect 29362 6300 29372 6356
rect 29428 6300 29708 6356
rect 29764 6300 30604 6356
rect 30660 6300 30670 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 44482 6188 44492 6244
rect 44548 6188 48748 6244
rect 48804 6188 48814 6244
rect 6626 6076 6636 6132
rect 6692 6076 7308 6132
rect 7364 6076 8652 6132
rect 8708 6076 9100 6132
rect 9156 6076 9166 6132
rect 10210 6076 10220 6132
rect 10276 6076 12796 6132
rect 12852 6076 13244 6132
rect 13300 6076 14028 6132
rect 14084 6076 14364 6132
rect 14420 6076 18060 6132
rect 18116 6076 18126 6132
rect 26002 6076 26012 6132
rect 26068 6076 26572 6132
rect 26628 6076 29372 6132
rect 29428 6076 29438 6132
rect 30594 6076 30604 6132
rect 30660 6076 33180 6132
rect 33236 6076 33246 6132
rect 44034 6076 44044 6132
rect 44100 6076 45276 6132
rect 45332 6076 45342 6132
rect 47954 6076 47964 6132
rect 48020 6076 53788 6132
rect 53844 6076 53854 6132
rect 10220 6020 10276 6076
rect 8306 5964 8316 6020
rect 8372 5964 10276 6020
rect 24210 5964 24220 6020
rect 24276 5964 25900 6020
rect 25956 5964 26460 6020
rect 26516 5964 26526 6020
rect 35522 5964 35532 6020
rect 35588 5964 36988 6020
rect 37044 5964 42476 6020
rect 42532 5964 42542 6020
rect 45490 5964 45500 6020
rect 45556 5964 46284 6020
rect 46340 5964 47068 6020
rect 47124 5964 47134 6020
rect 15698 5852 15708 5908
rect 15764 5852 16716 5908
rect 16772 5852 17948 5908
rect 18004 5852 18014 5908
rect 18274 5852 18284 5908
rect 18340 5852 21980 5908
rect 22036 5852 22046 5908
rect 23090 5852 23100 5908
rect 23156 5852 23548 5908
rect 23604 5852 23614 5908
rect 32498 5852 32508 5908
rect 32564 5852 33852 5908
rect 33908 5852 33918 5908
rect 34738 5852 34748 5908
rect 34804 5852 35308 5908
rect 35364 5852 35374 5908
rect 37650 5852 37660 5908
rect 37716 5852 39452 5908
rect 39508 5852 39518 5908
rect 43922 5852 43932 5908
rect 43988 5852 44604 5908
rect 44660 5852 45388 5908
rect 45444 5852 45454 5908
rect 46162 5852 46172 5908
rect 46228 5852 46956 5908
rect 47012 5852 47022 5908
rect 20178 5740 20188 5796
rect 20244 5740 30828 5796
rect 30884 5740 30894 5796
rect 35634 5740 35644 5796
rect 35700 5740 43260 5796
rect 43316 5740 44044 5796
rect 44100 5740 44110 5796
rect 10770 5628 10780 5684
rect 10836 5628 14252 5684
rect 14308 5628 16604 5684
rect 16660 5628 16670 5684
rect 19842 5628 19852 5684
rect 19908 5628 20300 5684
rect 20356 5628 20366 5684
rect 26226 5628 26236 5684
rect 26292 5628 26908 5684
rect 26964 5628 27580 5684
rect 27636 5628 27646 5684
rect 46274 5628 46284 5684
rect 46340 5628 47292 5684
rect 47348 5628 47358 5684
rect 13794 5516 13804 5572
rect 13860 5516 30268 5572
rect 30324 5516 31612 5572
rect 31668 5516 31678 5572
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 13122 5404 13132 5460
rect 13188 5404 20188 5460
rect 20244 5404 20254 5460
rect 25890 5404 25900 5460
rect 25956 5404 26348 5460
rect 26404 5404 27020 5460
rect 27076 5404 27468 5460
rect 27524 5404 28476 5460
rect 28532 5404 28542 5460
rect 16034 5292 16044 5348
rect 16100 5292 21644 5348
rect 21700 5292 21710 5348
rect 24546 5292 24556 5348
rect 24612 5292 27132 5348
rect 27188 5292 27804 5348
rect 27860 5292 27870 5348
rect 40898 5292 40908 5348
rect 40964 5292 41468 5348
rect 41524 5292 41534 5348
rect 48514 5292 48524 5348
rect 48580 5292 48748 5348
rect 48804 5292 48814 5348
rect 5058 5180 5068 5236
rect 5124 5180 5964 5236
rect 6020 5180 6030 5236
rect 13020 5180 13580 5236
rect 13636 5180 15484 5236
rect 15540 5180 16380 5236
rect 16436 5180 16446 5236
rect 16594 5180 16604 5236
rect 16660 5180 33628 5236
rect 33684 5180 33694 5236
rect 36642 5180 36652 5236
rect 36708 5180 38220 5236
rect 38276 5180 38286 5236
rect 42914 5180 42924 5236
rect 42980 5180 43820 5236
rect 43876 5180 43886 5236
rect 45826 5180 45836 5236
rect 45892 5180 48076 5236
rect 48132 5180 49196 5236
rect 49252 5180 49262 5236
rect 13020 5124 13076 5180
rect 8306 5068 8316 5124
rect 8372 5068 13076 5124
rect 15362 5068 15372 5124
rect 15428 5068 16828 5124
rect 16884 5068 17612 5124
rect 17668 5068 17678 5124
rect 19058 5068 19068 5124
rect 19124 5068 20188 5124
rect 20290 5068 20300 5124
rect 20356 5068 22876 5124
rect 22932 5068 23212 5124
rect 23268 5068 23278 5124
rect 25442 5068 25452 5124
rect 25508 5068 26012 5124
rect 26068 5068 27692 5124
rect 27748 5068 27758 5124
rect 28914 5068 28924 5124
rect 28980 5068 29708 5124
rect 29764 5068 29774 5124
rect 35634 5068 35644 5124
rect 35700 5068 36428 5124
rect 36484 5068 37660 5124
rect 37716 5068 37726 5124
rect 38546 5068 38556 5124
rect 38612 5068 39228 5124
rect 39284 5068 39294 5124
rect 41794 5068 41804 5124
rect 41860 5068 44156 5124
rect 44212 5068 44222 5124
rect 48178 5068 48188 5124
rect 48244 5068 48972 5124
rect 49028 5068 49038 5124
rect 13020 5012 13076 5068
rect 13010 4956 13020 5012
rect 13076 4956 13086 5012
rect 20132 4900 20188 5068
rect 21858 4956 21868 5012
rect 21924 4956 24668 5012
rect 24724 4956 24734 5012
rect 33954 4956 33964 5012
rect 34020 4956 34972 5012
rect 35028 4956 35308 5012
rect 35364 4956 35374 5012
rect 41906 4956 41916 5012
rect 41972 4956 42476 5012
rect 42532 4956 42542 5012
rect 43138 4956 43148 5012
rect 43204 4956 44492 5012
rect 44548 4956 44558 5012
rect 18050 4844 18060 4900
rect 18116 4844 18284 4900
rect 18340 4844 18350 4900
rect 20132 4844 24108 4900
rect 24164 4844 25004 4900
rect 25060 4844 27580 4900
rect 27636 4844 28812 4900
rect 28868 4844 28878 4900
rect 30930 4844 30940 4900
rect 30996 4844 31836 4900
rect 31892 4844 31902 4900
rect 39778 4844 39788 4900
rect 39844 4844 40572 4900
rect 40628 4844 41692 4900
rect 41748 4844 42700 4900
rect 42756 4844 42766 4900
rect 28242 4732 28252 4788
rect 28308 4732 30380 4788
rect 30436 4732 34412 4788
rect 34468 4732 34478 4788
rect 42130 4732 42140 4788
rect 42196 4732 44380 4788
rect 44436 4732 45724 4788
rect 45780 4732 45790 4788
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 19618 4508 19628 4564
rect 19684 4508 21756 4564
rect 21812 4508 21822 4564
rect 24658 4508 24668 4564
rect 24724 4508 25788 4564
rect 25844 4508 25854 4564
rect 30370 4508 30380 4564
rect 30436 4508 30828 4564
rect 30884 4508 31500 4564
rect 31556 4508 32844 4564
rect 32900 4508 32910 4564
rect 40114 4508 40124 4564
rect 40180 4508 40684 4564
rect 40740 4508 40750 4564
rect 42018 4508 42028 4564
rect 42084 4508 43148 4564
rect 43204 4508 43214 4564
rect 44482 4508 44492 4564
rect 44548 4508 45724 4564
rect 45780 4508 45790 4564
rect 28466 4396 28476 4452
rect 28532 4396 29820 4452
rect 29876 4396 31948 4452
rect 32004 4396 34076 4452
rect 34132 4396 37604 4452
rect 44818 4396 44828 4452
rect 44884 4396 45612 4452
rect 45668 4396 45678 4452
rect 9090 4284 9100 4340
rect 9156 4284 9772 4340
rect 9828 4284 9838 4340
rect 21298 4284 21308 4340
rect 21364 4284 21532 4340
rect 21588 4284 22204 4340
rect 22260 4284 22270 4340
rect 26450 4284 26460 4340
rect 26516 4284 26796 4340
rect 26852 4284 28196 4340
rect 28354 4284 28364 4340
rect 28420 4284 29036 4340
rect 29092 4284 29708 4340
rect 29764 4284 29774 4340
rect 36530 4284 36540 4340
rect 36596 4284 37212 4340
rect 37268 4284 37278 4340
rect 28140 4228 28196 4284
rect 7634 4172 7644 4228
rect 7700 4172 10220 4228
rect 10276 4172 10286 4228
rect 21634 4172 21644 4228
rect 21700 4172 22652 4228
rect 22708 4172 26908 4228
rect 26964 4172 26974 4228
rect 28130 4172 28140 4228
rect 28196 4172 28206 4228
rect 28364 4116 28420 4284
rect 35410 4172 35420 4228
rect 35476 4172 36988 4228
rect 37044 4172 37324 4228
rect 37380 4172 37390 4228
rect 4274 4060 4284 4116
rect 4340 4060 11228 4116
rect 11284 4060 11294 4116
rect 26338 4060 26348 4116
rect 26404 4060 28420 4116
rect 35298 4060 35308 4116
rect 35364 4060 35532 4116
rect 35588 4060 36204 4116
rect 36260 4060 36270 4116
rect 37548 4004 37604 4396
rect 37874 4060 37884 4116
rect 37940 4060 39004 4116
rect 39060 4060 39070 4116
rect 39330 4060 39340 4116
rect 39396 4060 41020 4116
rect 41076 4060 41916 4116
rect 41972 4060 41982 4116
rect 37548 3948 43708 4004
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 37426 3836 37436 3892
rect 37492 3836 38780 3892
rect 38836 3836 41916 3892
rect 41972 3836 41982 3892
rect 43652 3780 43708 3948
rect 5730 3724 5740 3780
rect 5796 3724 6356 3780
rect 29698 3724 29708 3780
rect 29764 3724 30716 3780
rect 30772 3724 30782 3780
rect 31612 3724 33068 3780
rect 33124 3724 33134 3780
rect 34402 3724 34412 3780
rect 34468 3724 38668 3780
rect 43652 3724 47516 3780
rect 47572 3724 47582 3780
rect 6300 3556 6356 3724
rect 31612 3668 31668 3724
rect 38612 3668 38668 3724
rect 18162 3612 18172 3668
rect 18228 3612 19628 3668
rect 19684 3612 20748 3668
rect 20804 3612 22092 3668
rect 22148 3612 22158 3668
rect 24210 3612 24220 3668
rect 24276 3612 24668 3668
rect 24724 3612 25564 3668
rect 25620 3612 25630 3668
rect 26852 3612 31612 3668
rect 31668 3612 31678 3668
rect 32274 3612 32284 3668
rect 32340 3612 33852 3668
rect 33908 3612 33918 3668
rect 34514 3612 34524 3668
rect 34580 3612 35756 3668
rect 35812 3612 35822 3668
rect 38612 3612 39452 3668
rect 39508 3612 39518 3668
rect 26852 3556 26908 3612
rect 6290 3500 6300 3556
rect 6356 3500 7644 3556
rect 7700 3500 7710 3556
rect 17714 3500 17724 3556
rect 17780 3500 17948 3556
rect 18004 3500 18620 3556
rect 18676 3500 18686 3556
rect 21298 3500 21308 3556
rect 21364 3500 26908 3556
rect 28130 3500 28140 3556
rect 28196 3500 28700 3556
rect 28756 3500 29260 3556
rect 29316 3500 33572 3556
rect 33516 3444 33572 3500
rect 12898 3388 12908 3444
rect 12964 3388 13692 3444
rect 13748 3388 13758 3444
rect 27234 3388 27244 3444
rect 27300 3388 30156 3444
rect 30212 3388 30380 3444
rect 30436 3388 30446 3444
rect 33506 3388 33516 3444
rect 33572 3388 34972 3444
rect 35028 3388 35812 3444
rect 40338 3388 40348 3444
rect 40404 3388 41132 3444
rect 41188 3388 42028 3444
rect 42084 3388 42094 3444
rect 48066 3388 48076 3444
rect 48132 3388 48748 3444
rect 48804 3388 48814 3444
rect 56018 3388 56028 3444
rect 56084 3388 56588 3444
rect 56644 3388 56654 3444
rect 35756 3332 35812 3388
rect 14466 3276 14476 3332
rect 14532 3276 33628 3332
rect 33684 3276 33694 3332
rect 35756 3276 55356 3332
rect 55412 3276 55422 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
<< via3 >>
rect 3724 60844 3780 60900
rect 13692 60732 13748 60788
rect 16492 60620 16548 60676
rect 4476 60340 4532 60396
rect 4580 60340 4636 60396
rect 4684 60340 4740 60396
rect 35196 60340 35252 60396
rect 35300 60340 35356 60396
rect 35404 60340 35460 60396
rect 14924 59948 14980 60004
rect 11788 59724 11844 59780
rect 19836 59556 19892 59612
rect 19940 59556 19996 59612
rect 20044 59556 20100 59612
rect 50556 59556 50612 59612
rect 50660 59556 50716 59612
rect 50764 59556 50820 59612
rect 14700 59388 14756 59444
rect 14924 59388 14980 59444
rect 14700 58940 14756 58996
rect 4476 58772 4532 58828
rect 4580 58772 4636 58828
rect 4684 58772 4740 58828
rect 35196 58772 35252 58828
rect 35300 58772 35356 58828
rect 35404 58772 35460 58828
rect 13468 58716 13524 58772
rect 3388 58156 3444 58212
rect 10780 58044 10836 58100
rect 19836 57988 19892 58044
rect 19940 57988 19996 58044
rect 20044 57988 20100 58044
rect 50556 57988 50612 58044
rect 50660 57988 50716 58044
rect 50764 57988 50820 58044
rect 11900 57932 11956 57988
rect 4172 57820 4228 57876
rect 4956 57708 5012 57764
rect 22540 57708 22596 57764
rect 13468 57596 13524 57652
rect 5068 57484 5124 57540
rect 14364 57484 14420 57540
rect 19404 57260 19460 57316
rect 4476 57204 4532 57260
rect 4580 57204 4636 57260
rect 4684 57204 4740 57260
rect 35196 57204 35252 57260
rect 35300 57204 35356 57260
rect 35404 57204 35460 57260
rect 12124 57148 12180 57204
rect 22540 56924 22596 56980
rect 6748 56700 6804 56756
rect 25676 56700 25732 56756
rect 2604 56588 2660 56644
rect 6524 56588 6580 56644
rect 6860 56588 6916 56644
rect 13580 56588 13636 56644
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 11900 56140 11956 56196
rect 7308 55916 7364 55972
rect 17612 55916 17668 55972
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 4060 55580 4116 55636
rect 18396 55580 18452 55636
rect 4844 55468 4900 55524
rect 16828 55356 16884 55412
rect 3164 55244 3220 55300
rect 7196 55244 7252 55300
rect 16604 55020 16660 55076
rect 3612 54908 3668 54964
rect 17948 54908 18004 54964
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 9100 54684 9156 54740
rect 20188 54460 20244 54516
rect 3276 54348 3332 54404
rect 4172 54348 4228 54404
rect 5740 54348 5796 54404
rect 9996 54348 10052 54404
rect 11340 54348 11396 54404
rect 9772 54236 9828 54292
rect 8540 54124 8596 54180
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 13468 54012 13524 54068
rect 3500 53900 3556 53956
rect 23660 53900 23716 53956
rect 2940 53788 2996 53844
rect 4956 53676 5012 53732
rect 6972 53676 7028 53732
rect 8652 53676 8708 53732
rect 17724 53788 17780 53844
rect 22316 53788 22372 53844
rect 22428 53676 22484 53732
rect 24220 53676 24276 53732
rect 6636 53452 6692 53508
rect 11676 53452 11732 53508
rect 15372 53452 15428 53508
rect 22316 53340 22372 53396
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 16156 53228 16212 53284
rect 24220 53228 24276 53284
rect 4956 53116 5012 53172
rect 9884 53116 9940 53172
rect 26012 53116 26068 53172
rect 11116 53004 11172 53060
rect 13580 53004 13636 53060
rect 7196 52892 7252 52948
rect 22316 52892 22372 52948
rect 23660 52892 23716 52948
rect 24220 52892 24276 52948
rect 3388 52780 3444 52836
rect 18396 52780 18452 52836
rect 18956 52780 19012 52836
rect 2828 52668 2884 52724
rect 4956 52668 5012 52724
rect 16268 52668 16324 52724
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 8540 52220 8596 52276
rect 22316 52220 22372 52276
rect 3052 52108 3108 52164
rect 4956 52108 5012 52164
rect 8428 52108 8484 52164
rect 12460 52108 12516 52164
rect 13020 52108 13076 52164
rect 22428 52108 22484 52164
rect 10444 51996 10500 52052
rect 3164 51884 3220 51940
rect 19404 51772 19460 51828
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 9996 51660 10052 51716
rect 11452 51660 11508 51716
rect 8092 51436 8148 51492
rect 3500 51324 3556 51380
rect 2156 51212 2212 51268
rect 3164 51212 3220 51268
rect 3836 51100 3892 51156
rect 20972 50988 21028 51044
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 15932 50876 15988 50932
rect 5852 50764 5908 50820
rect 12460 50764 12516 50820
rect 13244 50764 13300 50820
rect 16716 50764 16772 50820
rect 2604 50652 2660 50708
rect 3164 50652 3220 50708
rect 5068 50652 5124 50708
rect 5740 50652 5796 50708
rect 2940 50540 2996 50596
rect 3836 50540 3892 50596
rect 9100 50540 9156 50596
rect 11228 50540 11284 50596
rect 11452 50428 11508 50484
rect 15148 50428 15204 50484
rect 15932 50428 15988 50484
rect 20188 50428 20244 50484
rect 3052 50316 3108 50372
rect 4060 50316 4116 50372
rect 7084 50204 7140 50260
rect 11900 50204 11956 50260
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 6972 50092 7028 50148
rect 19404 50092 19460 50148
rect 8540 49756 8596 49812
rect 13804 49756 13860 49812
rect 2940 49644 2996 49700
rect 8092 49644 8148 49700
rect 11228 49644 11284 49700
rect 18956 49644 19012 49700
rect 6748 49532 6804 49588
rect 10780 49532 10836 49588
rect 11004 49532 11060 49588
rect 11788 49420 11844 49476
rect 17836 49420 17892 49476
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 8876 49196 8932 49252
rect 9772 49196 9828 49252
rect 12124 49196 12180 49252
rect 16492 49196 16548 49252
rect 3612 49084 3668 49140
rect 6972 49084 7028 49140
rect 16156 49084 16212 49140
rect 6748 48972 6804 49028
rect 13132 48972 13188 49028
rect 17724 48972 17780 49028
rect 3500 48860 3556 48916
rect 3612 48748 3668 48804
rect 8540 48748 8596 48804
rect 12124 48748 12180 48804
rect 4172 48636 4228 48692
rect 7980 48636 8036 48692
rect 19292 48636 19348 48692
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 7532 48524 7588 48580
rect 2492 48412 2548 48468
rect 3052 48412 3108 48468
rect 10444 48412 10500 48468
rect 11676 48412 11732 48468
rect 21084 48412 21140 48468
rect 34972 48412 35028 48468
rect 17948 48300 18004 48356
rect 3052 48188 3108 48244
rect 8652 48188 8708 48244
rect 14364 48188 14420 48244
rect 16492 48188 16548 48244
rect 5292 48076 5348 48132
rect 13356 48076 13412 48132
rect 14924 48076 14980 48132
rect 17612 48076 17668 48132
rect 18956 48076 19012 48132
rect 16716 47964 16772 48020
rect 4060 47852 4116 47908
rect 7980 47852 8036 47908
rect 28476 47852 28532 47908
rect 34972 47852 35028 47908
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 4172 47740 4228 47796
rect 8988 47740 9044 47796
rect 2828 47628 2884 47684
rect 17724 47516 17780 47572
rect 3276 47404 3332 47460
rect 4060 47404 4116 47460
rect 5516 47404 5572 47460
rect 6524 47404 6580 47460
rect 12124 47404 12180 47460
rect 10556 47180 10612 47236
rect 11116 47180 11172 47236
rect 5068 47068 5124 47124
rect 5292 47068 5348 47124
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 15036 46956 15092 47012
rect 16828 46956 16884 47012
rect 34972 46956 35028 47012
rect 9884 46844 9940 46900
rect 11004 46844 11060 46900
rect 11228 46844 11284 46900
rect 16156 46844 16212 46900
rect 25564 46844 25620 46900
rect 6412 46732 6468 46788
rect 6636 46732 6692 46788
rect 13132 46732 13188 46788
rect 23100 46732 23156 46788
rect 15036 46620 15092 46676
rect 15260 46620 15316 46676
rect 16604 46620 16660 46676
rect 23548 46620 23604 46676
rect 5068 46508 5124 46564
rect 5852 46508 5908 46564
rect 11676 46508 11732 46564
rect 16380 46508 16436 46564
rect 23436 46508 23492 46564
rect 25676 46508 25732 46564
rect 32284 46396 32340 46452
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 3388 46172 3444 46228
rect 8092 46172 8148 46228
rect 8316 46172 8372 46228
rect 8876 46172 8932 46228
rect 9772 46172 9828 46228
rect 15372 46172 15428 46228
rect 25340 46172 25396 46228
rect 3948 45948 4004 46004
rect 7532 45948 7588 46004
rect 4284 45724 4340 45780
rect 6188 45612 6244 45668
rect 6860 45612 6916 45668
rect 7756 45612 7812 45668
rect 11788 45612 11844 45668
rect 22092 45612 22148 45668
rect 6972 45500 7028 45556
rect 13020 45500 13076 45556
rect 13916 45500 13972 45556
rect 20972 45500 21028 45556
rect 23548 45500 23604 45556
rect 24332 45500 24388 45556
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 9660 45388 9716 45444
rect 3164 45276 3220 45332
rect 6972 45276 7028 45332
rect 27580 45276 27636 45332
rect 29260 45276 29316 45332
rect 30940 45276 30996 45332
rect 2156 45164 2212 45220
rect 29596 45164 29652 45220
rect 7308 45052 7364 45108
rect 8204 45052 8260 45108
rect 4844 44940 4900 44996
rect 11564 44940 11620 44996
rect 16380 44940 16436 44996
rect 30940 44940 30996 44996
rect 11900 44828 11956 44884
rect 22204 44828 22260 44884
rect 4844 44716 4900 44772
rect 8540 44716 8596 44772
rect 27580 44716 27636 44772
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 7084 44604 7140 44660
rect 17500 44604 17556 44660
rect 20188 44492 20244 44548
rect 23548 44380 23604 44436
rect 5964 44268 6020 44324
rect 9660 44156 9716 44212
rect 22092 44156 22148 44212
rect 3052 44044 3108 44100
rect 5180 44044 5236 44100
rect 13356 44044 13412 44100
rect 17052 44044 17108 44100
rect 23548 44044 23604 44100
rect 23772 44044 23828 44100
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 25340 43820 25396 43876
rect 7868 43708 7924 43764
rect 10220 43708 10276 43764
rect 9772 43596 9828 43652
rect 10108 43596 10164 43652
rect 11228 43596 11284 43652
rect 11452 43596 11508 43652
rect 15260 43596 15316 43652
rect 18844 43596 18900 43652
rect 13244 43484 13300 43540
rect 16268 43484 16324 43540
rect 17276 43484 17332 43540
rect 3164 43372 3220 43428
rect 8652 43372 8708 43428
rect 14812 43372 14868 43428
rect 25564 43372 25620 43428
rect 27020 43372 27076 43428
rect 3836 43260 3892 43316
rect 13020 43260 13076 43316
rect 15036 43260 15092 43316
rect 26684 43148 26740 43204
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 15372 43036 15428 43092
rect 15708 43036 15764 43092
rect 16156 43036 16212 43092
rect 13468 42924 13524 42980
rect 18956 42924 19012 42980
rect 2940 42812 2996 42868
rect 6636 42812 6692 42868
rect 6972 42812 7028 42868
rect 13916 42812 13972 42868
rect 19516 42812 19572 42868
rect 27020 42812 27076 42868
rect 4060 42700 4116 42756
rect 8988 42700 9044 42756
rect 26796 42700 26852 42756
rect 4284 42588 4340 42644
rect 11564 42588 11620 42644
rect 6300 42476 6356 42532
rect 18284 42476 18340 42532
rect 16604 42364 16660 42420
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 13468 42252 13524 42308
rect 16268 42252 16324 42308
rect 18844 42252 18900 42308
rect 19404 42252 19460 42308
rect 20860 42252 20916 42308
rect 3724 42140 3780 42196
rect 2492 42028 2548 42084
rect 10892 42028 10948 42084
rect 5628 41916 5684 41972
rect 6188 41916 6244 41972
rect 7420 41916 7476 41972
rect 2940 41804 2996 41860
rect 5740 41804 5796 41860
rect 6972 41804 7028 41860
rect 17836 41804 17892 41860
rect 19628 41804 19684 41860
rect 15148 41692 15204 41748
rect 15484 41692 15540 41748
rect 16380 41692 16436 41748
rect 18732 41692 18788 41748
rect 21980 41692 22036 41748
rect 3612 41580 3668 41636
rect 9100 41580 9156 41636
rect 9996 41580 10052 41636
rect 15596 41580 15652 41636
rect 19628 41580 19684 41636
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 12684 41468 12740 41524
rect 13020 41468 13076 41524
rect 19068 41468 19124 41524
rect 19404 41356 19460 41412
rect 3500 41244 3556 41300
rect 5628 41132 5684 41188
rect 13468 41132 13524 41188
rect 15036 41132 15092 41188
rect 21532 41132 21588 41188
rect 6076 41020 6132 41076
rect 7420 41020 7476 41076
rect 15260 41020 15316 41076
rect 17612 41020 17668 41076
rect 4172 40908 4228 40964
rect 16716 40908 16772 40964
rect 19516 40796 19572 40852
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 9100 40684 9156 40740
rect 12684 40684 12740 40740
rect 15596 40684 15652 40740
rect 16604 40684 16660 40740
rect 16940 40684 16996 40740
rect 4844 40572 4900 40628
rect 6412 40572 6468 40628
rect 11676 40572 11732 40628
rect 14700 40572 14756 40628
rect 19180 40572 19236 40628
rect 5964 40460 6020 40516
rect 6636 40460 6692 40516
rect 7980 40460 8036 40516
rect 11228 40460 11284 40516
rect 12012 40460 12068 40516
rect 15036 40460 15092 40516
rect 15260 40460 15316 40516
rect 3388 40348 3444 40404
rect 6748 40348 6804 40404
rect 18508 40348 18564 40404
rect 15372 40236 15428 40292
rect 18844 40236 18900 40292
rect 19292 40236 19348 40292
rect 20188 40236 20244 40292
rect 3388 40012 3444 40068
rect 3948 40012 4004 40068
rect 5068 40012 5124 40068
rect 7308 40012 7364 40068
rect 8540 40012 8596 40068
rect 9996 40012 10052 40068
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 5628 39900 5684 39956
rect 7980 39900 8036 39956
rect 12012 39900 12068 39956
rect 3052 39788 3108 39844
rect 3500 39788 3556 39844
rect 27132 39788 27188 39844
rect 6300 39676 6356 39732
rect 15036 39676 15092 39732
rect 17724 39676 17780 39732
rect 7868 39564 7924 39620
rect 8092 39564 8148 39620
rect 11564 39564 11620 39620
rect 16716 39564 16772 39620
rect 18732 39564 18788 39620
rect 11900 39452 11956 39508
rect 14140 39452 14196 39508
rect 19628 39452 19684 39508
rect 3388 38892 3444 38948
rect 5180 39340 5236 39396
rect 13580 39340 13636 39396
rect 14700 39340 14756 39396
rect 15372 39340 15428 39396
rect 18844 39340 18900 39396
rect 6188 39228 6244 39284
rect 12012 39228 12068 39284
rect 16940 39228 16996 39284
rect 17276 39228 17332 39284
rect 17724 39228 17780 39284
rect 19292 39228 19348 39284
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 13804 39116 13860 39172
rect 14476 39116 14532 39172
rect 23100 39116 23156 39172
rect 3836 39004 3892 39060
rect 9772 39004 9828 39060
rect 12124 39004 12180 39060
rect 13916 39004 13972 39060
rect 15092 39004 15148 39060
rect 18956 39004 19012 39060
rect 4284 38892 4340 38948
rect 8092 38892 8148 38948
rect 14812 38892 14868 38948
rect 20636 38892 20692 38948
rect 2492 38780 2548 38836
rect 7644 38780 7700 38836
rect 7980 38780 8036 38836
rect 11788 38780 11844 38836
rect 13356 38780 13412 38836
rect 17388 38780 17444 38836
rect 21532 38780 21588 38836
rect 5628 38668 5684 38724
rect 6300 38668 6356 38724
rect 15148 38668 15204 38724
rect 15372 38668 15428 38724
rect 38668 38668 38724 38724
rect 6636 38444 6692 38500
rect 11228 38444 11284 38500
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 14252 38220 14308 38276
rect 7420 38108 7476 38164
rect 17052 38108 17108 38164
rect 4284 37996 4340 38052
rect 6524 37996 6580 38052
rect 18284 37996 18340 38052
rect 6188 37884 6244 37940
rect 14588 37884 14644 37940
rect 6412 37772 6468 37828
rect 18620 37772 18676 37828
rect 4956 37660 5012 37716
rect 17612 37660 17668 37716
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 3500 37548 3556 37604
rect 10780 37548 10836 37604
rect 11452 37548 11508 37604
rect 13804 37548 13860 37604
rect 14252 37548 14308 37604
rect 5628 37436 5684 37492
rect 7084 37324 7140 37380
rect 9100 37324 9156 37380
rect 9884 37324 9940 37380
rect 12684 37212 12740 37268
rect 14924 37212 14980 37268
rect 20636 37212 20692 37268
rect 3388 37100 3444 37156
rect 5628 37100 5684 37156
rect 7980 37100 8036 37156
rect 19180 36988 19236 37044
rect 7868 36876 7924 36932
rect 13356 36876 13412 36932
rect 16828 36876 16884 36932
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 13580 36764 13636 36820
rect 10556 36652 10612 36708
rect 10892 36652 10948 36708
rect 14588 36652 14644 36708
rect 16492 36652 16548 36708
rect 9996 36540 10052 36596
rect 15148 36540 15204 36596
rect 18284 36540 18340 36596
rect 38668 36876 38724 36932
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 7644 36316 7700 36372
rect 10556 36316 10612 36372
rect 14140 36316 14196 36372
rect 14476 36316 14532 36372
rect 6412 36204 6468 36260
rect 12012 36092 12068 36148
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 13468 35868 13524 35924
rect 15148 35868 15204 35924
rect 19404 35868 19460 35924
rect 20412 35868 20468 35924
rect 20636 35868 20692 35924
rect 22204 35868 22260 35924
rect 32284 35868 32340 35924
rect 15260 35756 15316 35812
rect 17836 35756 17892 35812
rect 17388 35644 17444 35700
rect 3836 35532 3892 35588
rect 15484 35532 15540 35588
rect 22092 35532 22148 35588
rect 25788 35532 25844 35588
rect 26796 35532 26852 35588
rect 3724 35420 3780 35476
rect 3388 35308 3444 35364
rect 13580 35308 13636 35364
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 13804 35196 13860 35252
rect 26236 35196 26292 35252
rect 8204 35084 8260 35140
rect 12124 34972 12180 35028
rect 3388 34860 3444 34916
rect 5404 34860 5460 34916
rect 7308 34860 7364 34916
rect 10220 34860 10276 34916
rect 8092 34636 8148 34692
rect 15148 34636 15204 34692
rect 16828 34636 16884 34692
rect 21644 34636 21700 34692
rect 6524 34524 6580 34580
rect 16268 34524 16324 34580
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 4284 34412 4340 34468
rect 5404 34412 5460 34468
rect 5740 34412 5796 34468
rect 6412 34412 6468 34468
rect 17612 34412 17668 34468
rect 4172 34300 4228 34356
rect 10780 34076 10836 34132
rect 3612 33964 3668 34020
rect 23100 33964 23156 34020
rect 18508 33852 18564 33908
rect 22652 33852 22708 33908
rect 25564 33852 25620 33908
rect 25676 33740 25732 33796
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 20524 33628 20580 33684
rect 23436 33628 23492 33684
rect 5516 33516 5572 33572
rect 8652 33516 8708 33572
rect 15148 33404 15204 33460
rect 15596 33404 15652 33460
rect 18508 33404 18564 33460
rect 19516 33404 19572 33460
rect 20412 33404 20468 33460
rect 14252 33180 14308 33236
rect 17724 33068 17780 33124
rect 22652 33068 22708 33124
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 14364 32732 14420 32788
rect 15036 32732 15092 32788
rect 17724 32732 17780 32788
rect 26572 32732 26628 32788
rect 3612 32620 3668 32676
rect 10780 32620 10836 32676
rect 5628 32508 5684 32564
rect 13580 32508 13636 32564
rect 15708 32396 15764 32452
rect 13580 32284 13636 32340
rect 27692 32284 27748 32340
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 14476 32060 14532 32116
rect 18508 32060 18564 32116
rect 3612 31836 3668 31892
rect 18508 31836 18564 31892
rect 34972 31836 35028 31892
rect 8204 31724 8260 31780
rect 10220 31724 10276 31780
rect 15036 31724 15092 31780
rect 21980 31724 22036 31780
rect 8652 31612 8708 31668
rect 36876 31612 36932 31668
rect 38780 31612 38836 31668
rect 28364 31500 28420 31556
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 21644 31164 21700 31220
rect 15148 30940 15204 30996
rect 3948 30828 4004 30884
rect 11228 30828 11284 30884
rect 11116 30604 11172 30660
rect 25564 30604 25620 30660
rect 38780 30604 38836 30660
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 30380 30492 30436 30548
rect 19068 30380 19124 30436
rect 7756 30156 7812 30212
rect 25676 30156 25732 30212
rect 31948 30156 32004 30212
rect 19292 30044 19348 30100
rect 10444 29932 10500 29988
rect 33852 29932 33908 29988
rect 6412 29820 6468 29876
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 11676 29708 11732 29764
rect 3500 29596 3556 29652
rect 4060 29596 4116 29652
rect 25676 29596 25732 29652
rect 26012 29596 26068 29652
rect 33404 29596 33460 29652
rect 8316 29484 8372 29540
rect 11004 29484 11060 29540
rect 27132 29484 27188 29540
rect 9884 29372 9940 29428
rect 31948 29372 32004 29428
rect 11116 29260 11172 29316
rect 21084 29260 21140 29316
rect 26236 29148 26292 29204
rect 3948 29036 4004 29092
rect 14028 29036 14084 29092
rect 17612 29036 17668 29092
rect 34524 29036 34580 29092
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 34972 29148 35028 29204
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 57708 28924 57764 28980
rect 7756 28812 7812 28868
rect 17612 28812 17668 28868
rect 39788 28812 39844 28868
rect 3500 28700 3556 28756
rect 6412 28700 6468 28756
rect 17724 28588 17780 28644
rect 25676 28588 25732 28644
rect 27804 28588 27860 28644
rect 34524 28588 34580 28644
rect 8988 28476 9044 28532
rect 13692 28476 13748 28532
rect 57708 28476 57764 28532
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 9996 27916 10052 27972
rect 36540 27916 36596 27972
rect 27804 27804 27860 27860
rect 8988 27692 9044 27748
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 26236 27356 26292 27412
rect 31836 27356 31892 27412
rect 8316 27132 8372 27188
rect 36876 27132 36932 27188
rect 8092 27020 8148 27076
rect 33852 27020 33908 27076
rect 11452 26908 11508 26964
rect 34972 26908 35028 26964
rect 36540 26796 36596 26852
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 11564 26572 11620 26628
rect 6524 26348 6580 26404
rect 28476 26348 28532 26404
rect 30156 26348 30212 26404
rect 26012 26236 26068 26292
rect 39788 26236 39844 26292
rect 11452 26124 11508 26180
rect 20524 26124 20580 26180
rect 25676 26012 25732 26068
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 28476 25788 28532 25844
rect 4284 25676 4340 25732
rect 28364 25340 28420 25396
rect 31836 25340 31892 25396
rect 4284 25228 4340 25284
rect 23548 25228 23604 25284
rect 5628 25116 5684 25172
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 6076 25004 6132 25060
rect 13692 25004 13748 25060
rect 3836 24892 3892 24948
rect 31836 24892 31892 24948
rect 33852 24892 33908 24948
rect 11676 24668 11732 24724
rect 14028 24444 14084 24500
rect 26236 24444 26292 24500
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 8316 24220 8372 24276
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 10444 23996 10500 24052
rect 14252 23884 14308 23940
rect 8204 23772 8260 23828
rect 26572 23772 26628 23828
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 20524 23436 20580 23492
rect 30380 23436 30436 23492
rect 30604 23212 30660 23268
rect 11228 23100 11284 23156
rect 30716 23100 30772 23156
rect 31164 22988 31220 23044
rect 30156 22876 30212 22932
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 28812 22652 28868 22708
rect 33852 22652 33908 22708
rect 3724 22540 3780 22596
rect 23100 22540 23156 22596
rect 10220 22428 10276 22484
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 27692 21756 27748 21812
rect 8540 21644 8596 21700
rect 26796 21644 26852 21700
rect 30604 21644 30660 21700
rect 26348 21532 26404 21588
rect 28700 21420 28756 21476
rect 8204 21196 8260 21252
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 8540 21084 8596 21140
rect 28700 20860 28756 20916
rect 22092 20748 22148 20804
rect 27356 20748 27412 20804
rect 33404 20748 33460 20804
rect 26796 20636 26852 20692
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 7980 20300 8036 20356
rect 27692 20076 27748 20132
rect 27692 19852 27748 19908
rect 23212 19740 23268 19796
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 31164 19404 31220 19460
rect 11004 19292 11060 19348
rect 28812 19292 28868 19348
rect 30156 19068 30212 19124
rect 30716 18956 30772 19012
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 29596 18508 29652 18564
rect 28812 18396 28868 18452
rect 35644 18508 35700 18564
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 35868 17500 35924 17556
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 26348 17052 26404 17108
rect 31164 17052 31220 17108
rect 35756 16828 35812 16884
rect 30604 16716 30660 16772
rect 30380 16492 30436 16548
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 26796 16268 26852 16324
rect 29596 16156 29652 16212
rect 30716 16156 30772 16212
rect 35868 16156 35924 16212
rect 24332 16044 24388 16100
rect 31276 16044 31332 16100
rect 35756 15820 35812 15876
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 31276 15484 31332 15540
rect 29596 15260 29652 15316
rect 6300 15036 6356 15092
rect 18620 15036 18676 15092
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 35644 14700 35700 14756
rect 30716 14588 30772 14644
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 31164 13804 31220 13860
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 17500 13132 17556 13188
rect 23212 12796 23268 12852
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 35644 12348 35700 12404
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 23772 10668 23828 10724
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 25788 9212 25844 9268
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 26012 8316 26068 8372
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 20860 7532 20916 7588
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
<< metal4 >>
rect 3724 60900 3780 60910
rect 3388 58212 3444 58222
rect 2604 56644 2660 56654
rect 2156 51268 2212 51278
rect 2156 45220 2212 51212
rect 2604 50708 2660 56588
rect 3388 55468 3444 58156
rect 3276 55412 3444 55468
rect 3164 55300 3220 55310
rect 2940 53844 2996 53854
rect 2604 50642 2660 50652
rect 2828 52724 2884 52734
rect 2156 45154 2212 45164
rect 2492 48468 2548 48478
rect 2492 42084 2548 48412
rect 2828 47684 2884 52668
rect 2940 50596 2996 53788
rect 2940 50530 2996 50540
rect 3052 52164 3108 52174
rect 3052 50372 3108 52108
rect 3164 51940 3220 55244
rect 3164 51268 3220 51884
rect 3164 51202 3220 51212
rect 3276 54404 3332 55412
rect 2828 47618 2884 47628
rect 2940 49700 2996 49710
rect 2492 38836 2548 42028
rect 2940 42868 2996 49644
rect 3052 48468 3108 50316
rect 3052 48402 3108 48412
rect 3164 50708 3220 50718
rect 2940 41860 2996 42812
rect 2940 41794 2996 41804
rect 3052 48244 3108 48254
rect 3052 44100 3108 48188
rect 3052 39844 3108 44044
rect 3164 45332 3220 50652
rect 3276 47460 3332 54348
rect 3612 54964 3668 54974
rect 3500 53956 3556 53966
rect 3276 47394 3332 47404
rect 3388 52836 3444 52846
rect 3164 43428 3220 45276
rect 3164 43362 3220 43372
rect 3388 46228 3444 52780
rect 3500 51380 3556 53900
rect 3500 51314 3556 51324
rect 3612 49140 3668 54908
rect 3612 49074 3668 49084
rect 3388 40404 3444 46172
rect 3500 48916 3556 48926
rect 3500 41300 3556 48860
rect 3612 48804 3668 48814
rect 3612 41636 3668 48748
rect 3724 42196 3780 60844
rect 13692 60788 13748 60798
rect 4448 60396 4768 60428
rect 4448 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4768 60396
rect 4448 58828 4768 60340
rect 4448 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4768 58828
rect 4172 57876 4228 57886
rect 4060 55636 4116 55646
rect 3836 51156 3892 51166
rect 3836 50596 3892 51100
rect 3836 50530 3892 50540
rect 4060 50372 4116 55580
rect 4172 54404 4228 57820
rect 4172 54338 4228 54348
rect 4448 57260 4768 58772
rect 11788 59780 11844 59790
rect 10780 58100 10836 58110
rect 4448 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4768 57260
rect 4448 55692 4768 57204
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4060 47908 4116 50316
rect 4448 54124 4768 55636
rect 4956 57764 5012 57774
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4060 47842 4116 47852
rect 4172 48692 4228 48702
rect 4172 47796 4228 48636
rect 4172 47730 4228 47740
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4060 47460 4116 47470
rect 3948 46004 4004 46014
rect 3724 42130 3780 42140
rect 3836 43316 3892 43326
rect 3612 41570 3668 41580
rect 3500 41234 3556 41244
rect 3388 40338 3444 40348
rect 3052 39778 3108 39788
rect 3388 40068 3444 40078
rect 3388 38948 3444 40012
rect 3388 38882 3444 38892
rect 3500 39844 3556 39854
rect 2492 38770 2548 38780
rect 3500 37604 3556 39788
rect 3836 39060 3892 43260
rect 3948 40068 4004 45948
rect 3948 40002 4004 40012
rect 4060 42756 4116 47404
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 3836 38994 3892 39004
rect 3388 37156 3444 37166
rect 3388 35364 3444 37100
rect 3388 34916 3444 35308
rect 3388 34850 3444 34860
rect 3500 29652 3556 37548
rect 3836 35588 3892 35598
rect 3724 35476 3780 35486
rect 3612 34020 3668 34030
rect 3612 32676 3668 33964
rect 3612 31892 3668 32620
rect 3612 31826 3668 31836
rect 3500 28756 3556 29596
rect 3500 28690 3556 28700
rect 3724 22596 3780 35420
rect 3836 24948 3892 35532
rect 3948 30884 4004 30894
rect 3948 29092 4004 30828
rect 4060 29652 4116 42700
rect 4284 45780 4340 45790
rect 4284 42644 4340 45724
rect 4172 40964 4228 40974
rect 4172 34356 4228 40908
rect 4284 38948 4340 42588
rect 4284 38882 4340 38892
rect 4448 44716 4768 46228
rect 4844 55524 4900 55534
rect 4844 44996 4900 55468
rect 4956 53732 5012 57708
rect 4956 53172 5012 53676
rect 4956 52724 5012 53116
rect 4956 52658 5012 52668
rect 5068 57540 5124 57550
rect 4844 44930 4900 44940
rect 4956 52164 5012 52174
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4844 44772 4900 44782
rect 4844 40628 4900 44716
rect 4844 40562 4900 40572
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4172 34290 4228 34300
rect 4284 38052 4340 38062
rect 4284 34468 4340 37996
rect 4060 29586 4116 29596
rect 3948 29026 4004 29036
rect 4284 25732 4340 34412
rect 4284 25284 4340 25676
rect 4284 25218 4340 25228
rect 4448 36876 4768 38388
rect 4956 37716 5012 52108
rect 5068 50708 5124 57484
rect 6748 56756 6804 56766
rect 6524 56644 6580 56654
rect 5068 47124 5124 50652
rect 5740 54404 5796 54414
rect 5740 50708 5796 54348
rect 5740 50642 5796 50652
rect 5852 50820 5908 50830
rect 5068 47058 5124 47068
rect 5292 48132 5348 48142
rect 5292 47124 5348 48076
rect 5292 47058 5348 47068
rect 5516 47460 5572 47470
rect 5068 46564 5124 46574
rect 5068 40068 5124 46508
rect 5068 40002 5124 40012
rect 5180 44100 5236 44110
rect 5180 39396 5236 44044
rect 5180 39330 5236 39340
rect 4956 37650 5012 37660
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 5404 34916 5460 34926
rect 5404 34468 5460 34860
rect 5404 34402 5460 34412
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 5516 33572 5572 47404
rect 5852 46564 5908 50764
rect 6524 47460 6580 56588
rect 6524 47394 6580 47404
rect 6636 53508 6692 53518
rect 6636 49028 6692 53452
rect 6748 49588 6804 56700
rect 6748 49522 6804 49532
rect 6860 56644 6916 56654
rect 6748 49028 6804 49038
rect 6636 48972 6748 49028
rect 5852 46498 5908 46508
rect 6412 46788 6468 46798
rect 6188 45668 6244 45678
rect 5964 44324 6020 44334
rect 5628 41972 5684 41982
rect 5628 41188 5684 41916
rect 5628 39956 5684 41132
rect 5628 38724 5684 39900
rect 5628 38658 5684 38668
rect 5740 41860 5796 41870
rect 5516 33506 5572 33516
rect 5628 37492 5684 37502
rect 5628 37156 5684 37436
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 3836 24882 3892 24892
rect 3724 22530 3780 22540
rect 4448 24332 4768 25844
rect 5628 32564 5684 37100
rect 5740 34468 5796 41804
rect 5964 40516 6020 44268
rect 6188 41972 6244 45612
rect 5964 40450 6020 40460
rect 6076 41076 6132 41086
rect 5740 34402 5796 34412
rect 5628 25172 5684 32508
rect 5628 25106 5684 25116
rect 6076 25060 6132 41020
rect 6188 39284 6244 41916
rect 6300 42532 6356 42542
rect 6300 39732 6356 42476
rect 6412 40628 6468 46732
rect 6636 46788 6692 48972
rect 6748 48962 6804 48972
rect 6636 42868 6692 46732
rect 6860 45668 6916 56588
rect 7308 55972 7364 55982
rect 7196 55300 7252 55310
rect 6972 53732 7028 53742
rect 6972 50148 7028 53676
rect 7196 52948 7252 55244
rect 7196 52882 7252 52892
rect 6972 49140 7028 50092
rect 6972 49074 7028 49084
rect 7084 50260 7140 50270
rect 7084 47068 7140 50204
rect 6860 45602 6916 45612
rect 6972 47012 7140 47068
rect 6972 45556 7028 47012
rect 6972 45332 7028 45500
rect 6972 45266 7028 45276
rect 7308 45108 7364 55916
rect 9100 54740 9156 54750
rect 8540 54180 8596 54190
rect 8540 52276 8596 54124
rect 8428 52164 8484 52174
rect 8092 51492 8148 51502
rect 8092 49700 8148 51436
rect 8092 49634 8148 49644
rect 7980 48692 8036 48702
rect 7532 48580 7588 48590
rect 7532 46004 7588 48524
rect 7980 47908 8036 48636
rect 7980 47068 8036 47852
rect 7532 45938 7588 45948
rect 7644 47012 8036 47068
rect 7308 45042 7364 45052
rect 7084 44660 7140 44670
rect 6972 42868 7028 42878
rect 6692 42812 6804 42868
rect 6636 42802 6692 42812
rect 6468 40572 6580 40628
rect 6412 40562 6468 40572
rect 6300 39666 6356 39676
rect 6188 37940 6244 39228
rect 6188 37874 6244 37884
rect 6300 38724 6356 38734
rect 6076 24994 6132 25004
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 6300 15092 6356 38668
rect 6524 38052 6580 40572
rect 6636 40516 6692 40526
rect 6636 38500 6692 40460
rect 6748 40404 6804 42812
rect 6972 41860 7028 42812
rect 6972 41794 7028 41804
rect 6748 40338 6804 40348
rect 6636 38434 6692 38444
rect 6524 37986 6580 37996
rect 6412 37828 6468 37838
rect 6412 36260 6468 37772
rect 7084 37380 7140 44604
rect 7420 41972 7476 41982
rect 7420 41076 7476 41916
rect 7084 37314 7140 37324
rect 7308 40068 7364 40078
rect 6412 36194 6468 36204
rect 7308 34916 7364 40012
rect 7420 38164 7476 41020
rect 7420 38098 7476 38108
rect 7644 38836 7700 47012
rect 8092 46228 8148 46238
rect 7644 36372 7700 38780
rect 7644 36306 7700 36316
rect 7756 45668 7812 45678
rect 7308 34850 7364 34860
rect 6524 34580 6580 34590
rect 6412 34468 6468 34478
rect 6412 29876 6468 34412
rect 6412 28756 6468 29820
rect 6412 28690 6468 28700
rect 6524 26404 6580 34524
rect 7756 30212 7812 45612
rect 7868 43764 7924 43774
rect 7868 39620 7924 43708
rect 7980 40516 8036 40526
rect 7980 39956 8036 40460
rect 7980 39890 8036 39900
rect 7868 39554 7924 39564
rect 8092 39620 8148 46172
rect 8316 46228 8372 46238
rect 8428 46228 8484 52108
rect 8540 49812 8596 52220
rect 8540 49746 8596 49756
rect 8652 53732 8708 53742
rect 8372 46172 8484 46228
rect 8540 48804 8596 48814
rect 8316 46162 8372 46172
rect 8092 38948 8148 39564
rect 7980 38836 8036 38846
rect 7980 38668 8036 38780
rect 7868 38612 8036 38668
rect 7868 36932 7924 38612
rect 7868 36866 7924 36876
rect 7980 37156 8036 37166
rect 7756 28868 7812 30156
rect 7756 28802 7812 28812
rect 6524 26338 6580 26348
rect 7980 20356 8036 37100
rect 8092 34916 8148 38892
rect 8204 45108 8260 45118
rect 8204 35140 8260 45052
rect 8540 44772 8596 48748
rect 8652 48244 8708 53676
rect 9100 50596 9156 54684
rect 9996 54404 10052 54414
rect 9100 50428 9156 50540
rect 8652 48178 8708 48188
rect 8876 50372 9156 50428
rect 9772 54292 9828 54302
rect 8876 49252 8932 50372
rect 8876 46228 8932 49196
rect 9772 49252 9828 54236
rect 9772 49186 9828 49196
rect 9884 53172 9940 53182
rect 8876 46162 8932 46172
rect 8988 47796 9044 47806
rect 8540 40068 8596 44716
rect 8540 40002 8596 40012
rect 8652 43428 8708 43438
rect 8260 35084 8372 35140
rect 8204 35074 8260 35084
rect 8092 34860 8260 34916
rect 8092 34692 8148 34702
rect 8092 27076 8148 34636
rect 8204 31780 8260 34860
rect 8204 31714 8260 31724
rect 8316 29540 8372 35084
rect 8652 33572 8708 43372
rect 8652 31668 8708 33516
rect 8652 31602 8708 31612
rect 8988 42756 9044 47740
rect 9884 46900 9940 53116
rect 9996 51716 10052 54348
rect 9996 51650 10052 51660
rect 10444 52052 10500 52062
rect 10444 48468 10500 51996
rect 10780 49588 10836 58044
rect 11340 54404 11396 54414
rect 11116 53060 11172 53070
rect 10780 49522 10836 49532
rect 11004 49588 11060 49598
rect 10444 48402 10500 48412
rect 9884 46834 9940 46844
rect 10556 47236 10612 47246
rect 9772 46228 9828 46238
rect 9660 45444 9716 45454
rect 9660 44212 9716 45388
rect 9660 44146 9716 44156
rect 8316 29474 8372 29484
rect 8988 28532 9044 42700
rect 9772 43652 9828 46172
rect 10220 43764 10276 43774
rect 9100 41636 9156 41646
rect 9100 40740 9156 41580
rect 9100 37380 9156 40684
rect 9772 39060 9828 43596
rect 10108 43652 10164 43662
rect 9996 41636 10052 41646
rect 10108 41636 10164 43596
rect 10052 41580 10164 41636
rect 9996 41570 10052 41580
rect 9772 38994 9828 39004
rect 9996 40068 10052 40078
rect 9100 37314 9156 37324
rect 9884 37380 9940 37390
rect 9884 29428 9940 37324
rect 9884 29362 9940 29372
rect 9996 36596 10052 40012
rect 8988 27748 9044 28476
rect 9996 27972 10052 36540
rect 10220 34916 10276 43708
rect 10556 36708 10612 47180
rect 11004 46900 11060 49532
rect 11116 47236 11172 53004
rect 11116 47170 11172 47180
rect 11228 50596 11284 50606
rect 11228 49700 11284 50540
rect 11004 46834 11060 46844
rect 11228 46900 11284 49644
rect 11228 46834 11284 46844
rect 11228 43652 11284 43662
rect 11340 43652 11396 54348
rect 11676 53508 11732 53518
rect 11284 43596 11396 43652
rect 11452 51716 11508 51726
rect 11452 50484 11508 51660
rect 11452 43652 11508 50428
rect 11676 48468 11732 53452
rect 11788 49476 11844 59724
rect 13468 58772 13524 58782
rect 11900 57988 11956 57998
rect 11900 56196 11956 57932
rect 13468 57652 13524 58716
rect 11900 50260 11956 56140
rect 11900 50194 11956 50204
rect 12124 57204 12180 57214
rect 11788 49410 11844 49420
rect 11676 48402 11732 48412
rect 12124 49252 12180 57148
rect 13468 54068 13524 57596
rect 13468 54002 13524 54012
rect 13580 56644 13636 56654
rect 13580 53060 13636 56588
rect 13580 52994 13636 53004
rect 12460 52164 12516 52174
rect 12460 50820 12516 52108
rect 12460 50754 12516 50764
rect 13020 52164 13076 52174
rect 12124 48804 12180 49196
rect 12124 47460 12180 48748
rect 12124 47394 12180 47404
rect 11676 46564 11732 46574
rect 11228 43586 11284 43596
rect 10892 42084 10948 42094
rect 10556 36372 10612 36652
rect 10556 36306 10612 36316
rect 10780 37604 10836 37614
rect 10220 34850 10276 34860
rect 10780 34132 10836 37548
rect 10892 36708 10948 42028
rect 11228 40516 11284 40526
rect 11228 38500 11284 40460
rect 11228 38434 11284 38444
rect 11452 37604 11508 43596
rect 11564 44996 11620 45006
rect 11564 42644 11620 44940
rect 11564 39620 11620 42588
rect 11564 39554 11620 39564
rect 11676 40628 11732 46508
rect 11676 38668 11732 40572
rect 11788 45668 11844 45678
rect 11788 38836 11844 45612
rect 13020 45556 13076 52108
rect 13244 50820 13300 50830
rect 13132 49028 13188 49038
rect 13132 46788 13188 48972
rect 13132 46722 13188 46732
rect 13020 45490 13076 45500
rect 11900 44884 11956 44894
rect 11900 39508 11956 44828
rect 13244 43540 13300 50764
rect 13692 50428 13748 60732
rect 16492 60676 16548 60686
rect 14924 60004 14980 60014
rect 14700 59444 14756 59454
rect 14700 58996 14756 59388
rect 14924 59444 14980 59948
rect 14924 59378 14980 59388
rect 14700 58930 14756 58940
rect 13468 50372 13748 50428
rect 14364 57540 14420 57550
rect 13356 48132 13412 48142
rect 13356 44100 13412 48076
rect 13356 44034 13412 44044
rect 13244 43474 13300 43484
rect 13020 43316 13076 43326
rect 12684 41524 12740 41534
rect 12684 40740 12740 41468
rect 13020 41524 13076 43260
rect 13468 42980 13524 50372
rect 13468 42308 13524 42924
rect 13468 42242 13524 42252
rect 13804 49812 13860 49822
rect 13020 41458 13076 41468
rect 12012 40516 12068 40526
rect 12012 39956 12068 40460
rect 12012 39890 12068 39900
rect 11900 39442 11956 39452
rect 11788 38770 11844 38780
rect 12012 39284 12068 39294
rect 11452 37538 11508 37548
rect 11564 38612 11732 38668
rect 10892 36642 10948 36652
rect 10780 32676 10836 34076
rect 10780 32610 10836 32620
rect 9996 27906 10052 27916
rect 10220 31780 10276 31790
rect 8988 27682 9044 27692
rect 8092 27010 8148 27020
rect 8316 27188 8372 27198
rect 8316 24276 8372 27132
rect 8204 24220 8316 24276
rect 8204 23828 8260 24220
rect 8316 24210 8372 24220
rect 8204 21252 8260 23772
rect 10220 22484 10276 31724
rect 11228 30884 11284 30894
rect 11116 30660 11172 30670
rect 10444 29988 10500 29998
rect 10444 24052 10500 29932
rect 10444 23986 10500 23996
rect 11004 29540 11060 29550
rect 10220 22418 10276 22428
rect 8204 21186 8260 21196
rect 8540 21700 8596 21710
rect 8540 21140 8596 21644
rect 8540 21074 8596 21084
rect 7980 20290 8036 20300
rect 11004 19348 11060 29484
rect 11116 29316 11172 30604
rect 11116 29250 11172 29260
rect 11228 23156 11284 30828
rect 11452 26964 11508 26974
rect 11452 26180 11508 26908
rect 11564 26628 11620 38612
rect 12012 36148 12068 39228
rect 12012 36082 12068 36092
rect 12124 39060 12180 39070
rect 12124 35028 12180 39004
rect 12684 37268 12740 40684
rect 13468 41188 13524 41198
rect 12684 37202 12740 37212
rect 13356 38836 13412 38846
rect 13356 36932 13412 38780
rect 13356 36866 13412 36876
rect 13468 35924 13524 41132
rect 13580 39396 13636 39406
rect 13580 36820 13636 39340
rect 13804 39172 13860 49756
rect 14364 48244 14420 57484
rect 15372 53508 15428 53518
rect 13804 39106 13860 39116
rect 13916 45556 13972 45566
rect 13916 42868 13972 45500
rect 13916 39060 13972 42812
rect 13916 38994 13972 39004
rect 14140 39508 14196 39518
rect 13580 36754 13636 36764
rect 13804 37604 13860 37614
rect 13468 35858 13524 35868
rect 12124 34962 12180 34972
rect 13580 35364 13636 35374
rect 13580 32564 13636 35308
rect 13804 35252 13860 37548
rect 14140 36372 14196 39452
rect 14252 38276 14308 38286
rect 14252 37604 14308 38220
rect 14252 37538 14308 37548
rect 14140 36306 14196 36316
rect 13804 35186 13860 35196
rect 13580 32340 13636 32508
rect 13580 32274 13636 32284
rect 14252 33236 14308 33246
rect 11564 26562 11620 26572
rect 11676 29764 11732 29774
rect 11452 26114 11508 26124
rect 11676 24724 11732 29708
rect 14028 29092 14084 29102
rect 13692 28532 13748 28542
rect 13692 25060 13748 28476
rect 13692 24994 13748 25004
rect 11676 24658 11732 24668
rect 14028 24500 14084 29036
rect 14028 24434 14084 24444
rect 14252 23940 14308 33180
rect 14364 32788 14420 48188
rect 15148 50484 15204 50494
rect 14924 48132 14980 48142
rect 14812 43428 14868 43438
rect 14700 40628 14756 40638
rect 14700 39396 14756 40572
rect 14700 39330 14756 39340
rect 14364 32722 14420 32732
rect 14476 39172 14532 39182
rect 14476 36372 14532 39116
rect 14812 38948 14868 43372
rect 14588 38892 14812 38948
rect 14588 37940 14644 38892
rect 14812 38882 14868 38892
rect 14588 36708 14644 37884
rect 14924 37268 14980 48076
rect 15036 47012 15092 47022
rect 15036 46676 15092 46956
rect 15036 43316 15092 46620
rect 15036 41188 15092 43260
rect 15148 41748 15204 50428
rect 15260 46676 15316 46686
rect 15260 43652 15316 46620
rect 15260 43586 15316 43596
rect 15372 46228 15428 53452
rect 16156 53284 16212 53294
rect 15932 50932 15988 50942
rect 15932 50484 15988 50876
rect 15932 50418 15988 50428
rect 16156 49140 16212 53228
rect 16156 49074 16212 49084
rect 16268 52724 16324 52734
rect 16268 47068 16324 52668
rect 16492 49252 16548 60620
rect 19808 59612 20128 60428
rect 19808 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20128 59612
rect 19808 58044 20128 59556
rect 19808 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20128 58044
rect 19404 57316 19460 57326
rect 17612 55972 17668 55982
rect 16828 55412 16884 55422
rect 16492 49186 16548 49196
rect 16604 55076 16660 55086
rect 16492 48244 16548 48254
rect 16268 47012 16436 47068
rect 15148 41682 15204 41692
rect 15372 43092 15428 46172
rect 16156 46900 16212 46910
rect 15036 41122 15092 41132
rect 15260 41076 15316 41086
rect 15148 41020 15260 41076
rect 15036 40516 15092 40526
rect 15148 40516 15204 41020
rect 15260 41010 15316 41020
rect 15092 40460 15204 40516
rect 15260 40516 15316 40526
rect 15036 40450 15092 40460
rect 15036 39732 15092 39742
rect 15036 39070 15092 39676
rect 15036 39060 15148 39070
rect 15036 39004 15092 39060
rect 15092 38994 15148 39004
rect 14924 37202 14980 37212
rect 15148 38724 15204 38734
rect 14588 36642 14644 36652
rect 14476 32116 14532 36316
rect 15148 36596 15204 38668
rect 15148 35924 15204 36540
rect 15148 34692 15204 35868
rect 15260 35812 15316 40460
rect 15372 40292 15428 43036
rect 15708 43092 15764 43102
rect 15372 39396 15428 40236
rect 15372 38724 15428 39340
rect 15372 38658 15428 38668
rect 15484 41748 15540 41758
rect 15260 35746 15316 35756
rect 15484 35588 15540 41692
rect 15484 35522 15540 35532
rect 15596 41636 15652 41646
rect 15596 40740 15652 41580
rect 15148 34626 15204 34636
rect 15148 33460 15204 33470
rect 14476 32050 14532 32060
rect 15036 32788 15092 32798
rect 15036 31780 15092 32732
rect 15036 31714 15092 31724
rect 15148 30996 15204 33404
rect 15596 33460 15652 40684
rect 15596 33394 15652 33404
rect 15708 32452 15764 43036
rect 16156 43092 16212 46844
rect 16380 46564 16436 47012
rect 16380 44996 16436 46508
rect 16156 43026 16212 43036
rect 16268 43540 16324 43550
rect 16268 42308 16324 43484
rect 16268 34580 16324 42252
rect 16380 41748 16436 44940
rect 16380 41682 16436 41692
rect 16492 36708 16548 48188
rect 16604 46676 16660 55020
rect 16716 50820 16772 50830
rect 16716 48020 16772 50764
rect 16716 47954 16772 47964
rect 16828 47012 16884 55356
rect 17612 48132 17668 55916
rect 18396 55636 18452 55646
rect 17948 54964 18004 54974
rect 17612 48066 17668 48076
rect 17724 53844 17780 53854
rect 17724 49028 17780 53788
rect 17724 47572 17780 48972
rect 17724 47506 17780 47516
rect 17836 49476 17892 49486
rect 16828 46946 16884 46956
rect 16604 42420 16660 46620
rect 17500 44660 17556 44670
rect 16604 40740 16660 42364
rect 17052 44100 17108 44110
rect 16604 40674 16660 40684
rect 16716 40964 16772 40974
rect 16716 39620 16772 40908
rect 16716 39554 16772 39564
rect 16940 40740 16996 40750
rect 16940 39284 16996 40684
rect 16940 39218 16996 39228
rect 17052 38164 17108 44044
rect 17276 43540 17332 43550
rect 17276 39284 17332 43484
rect 17276 39218 17332 39228
rect 17052 38098 17108 38108
rect 17388 38836 17444 38846
rect 16492 36642 16548 36652
rect 16828 36932 16884 36942
rect 16828 34692 16884 36876
rect 17388 35700 17444 38780
rect 17388 35634 17444 35644
rect 16828 34626 16884 34636
rect 16268 34514 16324 34524
rect 15708 32386 15764 32396
rect 15148 30930 15204 30940
rect 14252 23874 14308 23884
rect 11228 23090 11284 23100
rect 11004 19282 11060 19292
rect 6300 15026 6356 15036
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 17500 13188 17556 44604
rect 17836 41860 17892 49420
rect 17948 48356 18004 54908
rect 18396 52836 18452 55580
rect 18396 52770 18452 52780
rect 18956 52836 19012 52846
rect 17948 48290 18004 48300
rect 18956 49700 19012 52780
rect 19404 51828 19460 57260
rect 19404 50148 19460 51772
rect 19404 50082 19460 50092
rect 19808 56476 20128 57988
rect 35168 60396 35488 60428
rect 35168 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35488 60396
rect 35168 58828 35488 60340
rect 35168 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35488 58828
rect 22540 57764 22596 57774
rect 22540 56980 22596 57708
rect 22540 56914 22596 56924
rect 35168 57260 35488 58772
rect 35168 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35488 57260
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 25676 56756 25732 56766
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 20188 54516 20244 54526
rect 20188 50484 20244 54460
rect 23660 53956 23716 53966
rect 22316 53844 22372 53854
rect 22316 53396 22372 53788
rect 22316 52948 22372 53340
rect 22316 52276 22372 52892
rect 22316 52210 22372 52220
rect 22428 53732 22484 53742
rect 22428 52164 22484 53676
rect 23660 52948 23716 53900
rect 23660 52882 23716 52892
rect 24220 53732 24276 53742
rect 24220 53284 24276 53676
rect 24220 52948 24276 53228
rect 24220 52882 24276 52892
rect 22428 52098 22484 52108
rect 20188 50418 20244 50428
rect 20972 51044 21028 51054
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 18956 48132 19012 49644
rect 18956 48066 19012 48076
rect 19292 48692 19348 48702
rect 18844 43652 18900 43662
rect 17612 41076 17668 41086
rect 17612 37716 17668 41020
rect 17724 39732 17780 39742
rect 17724 39284 17780 39676
rect 17724 39218 17780 39228
rect 17612 37650 17668 37660
rect 17836 35812 17892 41804
rect 18284 42532 18340 42542
rect 18284 38052 18340 42476
rect 18844 42308 18900 43596
rect 18844 42242 18900 42252
rect 18956 42980 19012 42990
rect 18732 41748 18788 41758
rect 18284 36596 18340 37996
rect 18284 36530 18340 36540
rect 18508 40404 18564 40414
rect 17836 35746 17892 35756
rect 17612 34468 17668 34478
rect 17612 29092 17668 34412
rect 18508 33908 18564 40348
rect 18732 39620 18788 41692
rect 18732 39554 18788 39564
rect 18844 40292 18900 40302
rect 18844 39396 18900 40236
rect 18844 39330 18900 39340
rect 18956 39060 19012 42924
rect 18956 38994 19012 39004
rect 19068 41524 19124 41534
rect 18508 33842 18564 33852
rect 18620 37828 18676 37838
rect 18508 33460 18564 33470
rect 17612 28868 17668 29036
rect 17612 28802 17668 28812
rect 17724 33124 17780 33134
rect 17724 32788 17780 33068
rect 17724 28644 17780 32732
rect 18508 32116 18564 33404
rect 18508 31892 18564 32060
rect 18508 31826 18564 31836
rect 17724 28578 17780 28588
rect 18620 15092 18676 37772
rect 19068 30436 19124 41468
rect 19292 41188 19348 48636
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 20972 45556 21028 50988
rect 20972 45490 21028 45500
rect 21084 48468 21140 48478
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19516 42868 19572 42878
rect 19404 42308 19460 42318
rect 19404 41412 19460 42252
rect 19404 41346 19460 41356
rect 19292 41132 19460 41188
rect 19180 40628 19236 40638
rect 19180 37044 19236 40572
rect 19180 36978 19236 36988
rect 19292 40292 19348 40302
rect 19292 39284 19348 40236
rect 19068 30370 19124 30380
rect 19292 30100 19348 39228
rect 19404 35924 19460 41132
rect 19404 35858 19460 35868
rect 19516 40852 19572 42812
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19516 33460 19572 40796
rect 19628 41860 19684 41870
rect 19628 41636 19684 41804
rect 19628 39508 19684 41580
rect 19628 39442 19684 39452
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19516 33394 19572 33404
rect 19808 39228 20128 40740
rect 20188 44548 20244 44558
rect 20188 40292 20244 44492
rect 20188 40226 20244 40236
rect 20860 42308 20916 42318
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 20636 38948 20692 38958
rect 20636 37268 20692 38892
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19292 30034 19348 30044
rect 19808 32956 20128 34468
rect 20412 35924 20468 35934
rect 20412 33460 20468 35868
rect 20636 35924 20692 37212
rect 20636 35858 20692 35868
rect 20412 33394 20468 33404
rect 20524 33684 20580 33694
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 18620 15026 18676 15036
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 20524 26180 20580 33628
rect 20524 23492 20580 26124
rect 20524 23426 20580 23436
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 17500 13122 17556 13132
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 20860 7588 20916 42252
rect 21084 29316 21140 48412
rect 25564 46900 25620 46910
rect 23100 46788 23156 46798
rect 22092 45668 22148 45678
rect 22092 44212 22148 45612
rect 22092 44146 22148 44156
rect 22204 44884 22260 44894
rect 21980 41748 22036 41758
rect 21532 41188 21588 41198
rect 21532 38836 21588 41132
rect 21532 38770 21588 38780
rect 21644 34692 21700 34702
rect 21644 31220 21700 34636
rect 21980 31780 22036 41692
rect 22204 35924 22260 44828
rect 23100 39172 23156 46732
rect 23548 46676 23604 46686
rect 23100 39106 23156 39116
rect 23436 46564 23492 46574
rect 22204 35858 22260 35868
rect 21980 31714 22036 31724
rect 22092 35588 22148 35598
rect 21644 31154 21700 31164
rect 21084 29250 21140 29260
rect 22092 20804 22148 35532
rect 23100 34020 23156 34030
rect 22652 33908 22708 33918
rect 22652 33124 22708 33852
rect 22652 33058 22708 33068
rect 23100 22596 23156 33964
rect 23436 33684 23492 46508
rect 23548 45556 23604 46620
rect 25340 46228 25396 46238
rect 23548 45490 23604 45500
rect 24332 45556 24388 45566
rect 23436 33618 23492 33628
rect 23548 44436 23604 44446
rect 23548 44100 23604 44380
rect 23548 25284 23604 44044
rect 23548 25218 23604 25228
rect 23772 44100 23828 44110
rect 23100 22530 23156 22540
rect 22092 20738 22148 20748
rect 23212 19796 23268 19806
rect 23212 12852 23268 19740
rect 23212 12786 23268 12796
rect 23772 10724 23828 44044
rect 24332 16100 24388 45500
rect 25340 43876 25396 46172
rect 25340 43810 25396 43820
rect 25564 43428 25620 46844
rect 25676 46564 25732 56700
rect 35168 55692 35488 57204
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 25676 46498 25732 46508
rect 26012 53172 26068 53182
rect 25564 43362 25620 43372
rect 25788 35588 25844 35598
rect 25564 33908 25620 33918
rect 25564 30660 25620 33852
rect 25564 30594 25620 30604
rect 25676 33796 25732 33806
rect 25676 30212 25732 33740
rect 25676 30146 25732 30156
rect 25676 29652 25732 29662
rect 25676 28644 25732 29596
rect 25676 26068 25732 28588
rect 25676 26002 25732 26012
rect 24332 16034 24388 16044
rect 23772 10658 23828 10668
rect 25788 9268 25844 35532
rect 26012 29652 26068 53116
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 34972 48468 35028 48478
rect 28476 47908 28532 47918
rect 27580 45332 27636 45342
rect 27580 44772 27636 45276
rect 27580 44706 27636 44716
rect 27020 43428 27076 43438
rect 26684 43204 26740 43214
rect 26684 42756 26740 43148
rect 27020 42868 27076 43372
rect 27020 42802 27076 42812
rect 26796 42756 26852 42766
rect 26684 42700 26796 42756
rect 26796 35588 26852 42700
rect 26796 35522 26852 35532
rect 27132 39844 27188 39854
rect 26012 26292 26068 29596
rect 26236 35252 26292 35262
rect 26236 29204 26292 35196
rect 26236 29138 26292 29148
rect 26572 32788 26628 32798
rect 26012 26226 26068 26236
rect 26236 27412 26292 27422
rect 26236 24500 26292 27356
rect 26236 24434 26292 24444
rect 26572 23828 26628 32732
rect 27132 29540 27188 39788
rect 27132 26908 27188 29484
rect 27692 32340 27748 32350
rect 27132 26852 27412 26908
rect 26572 23762 26628 23772
rect 26796 21700 26852 21710
rect 26348 21588 26404 21598
rect 26348 17108 26404 21532
rect 26348 17042 26404 17052
rect 26796 20692 26852 21644
rect 27356 20804 27412 26852
rect 27356 20738 27412 20748
rect 27692 21812 27748 32284
rect 28364 31556 28420 31566
rect 27804 28644 27860 28654
rect 27804 27860 27860 28588
rect 27804 27794 27860 27804
rect 28364 25396 28420 31500
rect 28476 26404 28532 47852
rect 34972 47908 35028 48412
rect 34972 47842 35028 47852
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 34972 47012 35028 47022
rect 32284 46452 32340 46462
rect 29260 45332 29316 45342
rect 29260 45220 29316 45276
rect 30940 45332 30996 45342
rect 29596 45220 29652 45230
rect 29260 45164 29596 45220
rect 29596 45154 29652 45164
rect 30940 44996 30996 45276
rect 30940 44930 30996 44940
rect 32284 35924 32340 46396
rect 32284 35858 32340 35868
rect 34972 31892 35028 46956
rect 34972 31826 35028 31836
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 50528 59612 50848 60428
rect 50528 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50848 59612
rect 50528 58044 50848 59556
rect 50528 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50848 58044
rect 50528 56476 50848 57988
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 38668 38724 38724 38734
rect 38668 36932 38724 38668
rect 38668 36866 38724 36876
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 30380 30548 30436 30558
rect 28476 25844 28532 26348
rect 28476 25778 28532 25788
rect 30156 26404 30212 26414
rect 28364 25330 28420 25340
rect 30156 22932 30212 26348
rect 30380 23492 30436 30492
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 31948 30212 32004 30222
rect 31948 29428 32004 30156
rect 33852 29988 33908 29998
rect 31948 29362 32004 29372
rect 33404 29652 33460 29662
rect 31836 27412 31892 27422
rect 31836 25396 31892 27356
rect 31836 24948 31892 25340
rect 31836 24882 31892 24892
rect 30380 23426 30436 23436
rect 26796 16324 26852 20636
rect 27692 20132 27748 21756
rect 28812 22708 28868 22718
rect 28700 21476 28756 21486
rect 28700 20916 28756 21420
rect 28700 20850 28756 20860
rect 27692 19908 27748 20076
rect 27692 19842 27748 19852
rect 28812 19348 28868 22652
rect 28812 18452 28868 19292
rect 30156 19124 30212 22876
rect 30604 23268 30660 23278
rect 30604 21700 30660 23212
rect 30604 21634 30660 21644
rect 30716 23156 30772 23166
rect 30156 19058 30212 19068
rect 30716 19012 30772 23100
rect 30716 18946 30772 18956
rect 31164 23044 31220 23054
rect 31164 19460 31220 22988
rect 33404 20804 33460 29596
rect 33852 27076 33908 29932
rect 34972 29204 35028 29214
rect 34524 29092 34580 29102
rect 34524 28644 34580 29036
rect 34524 28578 34580 28588
rect 33852 27010 33908 27020
rect 34972 26964 35028 29148
rect 34972 26898 35028 26908
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 36876 31668 36932 31678
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 36540 27972 36596 27982
rect 36540 26852 36596 27916
rect 36876 27188 36932 31612
rect 38780 31668 38836 31678
rect 38780 30660 38836 31612
rect 38780 30594 38836 30604
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 36876 27122 36932 27132
rect 39788 28868 39844 28878
rect 36540 26786 36596 26796
rect 39788 26292 39844 28812
rect 39788 26226 39844 26236
rect 50528 28252 50848 29764
rect 57708 28980 57764 28990
rect 57708 28532 57764 28924
rect 57708 28466 57764 28476
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 33852 24948 33908 24958
rect 33852 22708 33908 24892
rect 33852 22642 33908 22652
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 33404 20738 33460 20748
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 28812 18386 28868 18396
rect 29596 18564 29652 18574
rect 26796 16258 26852 16268
rect 29596 16212 29652 18508
rect 31164 17108 31220 19404
rect 30604 16772 30660 16782
rect 30380 16548 30436 16558
rect 30604 16548 30660 16716
rect 30436 16492 30660 16548
rect 30380 16482 30436 16492
rect 29596 15316 29652 16156
rect 29596 15250 29652 15260
rect 30716 16212 30772 16222
rect 30716 14644 30772 16156
rect 30716 14578 30772 14588
rect 31164 13860 31220 17052
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 31276 16100 31332 16110
rect 31276 15540 31332 16044
rect 31276 15474 31332 15484
rect 31164 13794 31220 13804
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 25788 8428 25844 9212
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35644 18564 35700 18574
rect 35644 14756 35700 18508
rect 35868 17556 35924 17566
rect 35756 16884 35812 16894
rect 35756 15876 35812 16828
rect 35868 16212 35924 17500
rect 35868 16146 35924 16156
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 35756 15810 35812 15820
rect 35644 12404 35700 14700
rect 35644 12338 35700 12348
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 25788 8372 26068 8428
rect 26012 8306 26068 8316
rect 20860 7522 20916 7532
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1601__I Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 2688 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1602__A1
timestamp 1669390400
transform 1 0 16016 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1602__A2
timestamp 1669390400
transform 1 0 15568 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1603__I
timestamp 1669390400
transform 1 0 20832 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1604__I
timestamp 1669390400
transform 1 0 26432 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1605__A1
timestamp 1669390400
transform 1 0 14672 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1605__A2
timestamp 1669390400
transform 1 0 12208 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1606__I
timestamp 1669390400
transform -1 0 14672 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1608__A1
timestamp 1669390400
transform 1 0 3696 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1608__A2
timestamp 1669390400
transform 1 0 4144 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1610__A1
timestamp 1669390400
transform -1 0 2800 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1610__A2
timestamp 1669390400
transform 1 0 7840 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1611__A1
timestamp 1669390400
transform 1 0 2128 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1613__A1
timestamp 1669390400
transform -1 0 2800 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1613__A2
timestamp 1669390400
transform 1 0 4592 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1614__A1
timestamp 1669390400
transform 1 0 3136 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1614__A2
timestamp 1669390400
transform 1 0 7168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1615__A1
timestamp 1669390400
transform 1 0 6832 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1615__A2
timestamp 1669390400
transform 1 0 8960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1615__B
timestamp 1669390400
transform 1 0 7280 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1616__A1
timestamp 1669390400
transform 1 0 3360 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1616__A2
timestamp 1669390400
transform -1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1617__I
timestamp 1669390400
transform -1 0 5824 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1618__I
timestamp 1669390400
transform 1 0 2800 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1619__A1
timestamp 1669390400
transform -1 0 7168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1619__A2
timestamp 1669390400
transform -1 0 1904 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1621__I
timestamp 1669390400
transform 1 0 1904 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1622__A1
timestamp 1669390400
transform 1 0 3584 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1622__A2
timestamp 1669390400
transform 1 0 8400 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1624__I
timestamp 1669390400
transform -1 0 4032 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1625__A1
timestamp 1669390400
transform 1 0 3584 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1625__A2
timestamp 1669390400
transform 1 0 4480 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1627__I
timestamp 1669390400
transform 1 0 3248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1628__A1
timestamp 1669390400
transform -1 0 12096 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1628__A2
timestamp 1669390400
transform -1 0 10752 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1628__B
timestamp 1669390400
transform -1 0 11648 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1629__A1
timestamp 1669390400
transform 1 0 14560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1629__A2
timestamp 1669390400
transform 1 0 15008 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1630__I
timestamp 1669390400
transform 1 0 12096 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1631__A1
timestamp 1669390400
transform 1 0 8064 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1631__B
timestamp 1669390400
transform 1 0 10416 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1632__A1
timestamp 1669390400
transform 1 0 4928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1632__A2
timestamp 1669390400
transform 1 0 7392 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1633__I
timestamp 1669390400
transform 1 0 3472 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1635__I
timestamp 1669390400
transform 1 0 3024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1636__A1
timestamp 1669390400
transform 1 0 1904 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1636__A2
timestamp 1669390400
transform -1 0 2688 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1636__B
timestamp 1669390400
transform -1 0 1904 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1637__I
timestamp 1669390400
transform -1 0 2800 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1638__I
timestamp 1669390400
transform 1 0 9184 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1639__A1
timestamp 1669390400
transform -1 0 10976 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1639__A2
timestamp 1669390400
transform -1 0 10304 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1639__A3
timestamp 1669390400
transform -1 0 9856 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1640__A1
timestamp 1669390400
transform 1 0 2352 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1640__A2
timestamp 1669390400
transform 1 0 4368 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1640__B
timestamp 1669390400
transform -1 0 3024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1641__A1
timestamp 1669390400
transform -1 0 11424 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1641__A2
timestamp 1669390400
transform 1 0 10752 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1641__B2
timestamp 1669390400
transform -1 0 10528 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1642__I
timestamp 1669390400
transform 1 0 3920 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1643__A1
timestamp 1669390400
transform -1 0 13776 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1643__B2
timestamp 1669390400
transform 1 0 11872 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1644__I
timestamp 1669390400
transform 1 0 2128 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1645__A1
timestamp 1669390400
transform -1 0 8288 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1645__A2
timestamp 1669390400
transform 1 0 11088 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1646__A1
timestamp 1669390400
transform 1 0 12880 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1647__I
timestamp 1669390400
transform -1 0 4256 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1648__A1
timestamp 1669390400
transform 1 0 14896 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1648__A2
timestamp 1669390400
transform -1 0 12096 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1648__A3
timestamp 1669390400
transform -1 0 14224 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1648__A4
timestamp 1669390400
transform 1 0 12768 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1649__A1
timestamp 1669390400
transform 1 0 15344 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1650__A1
timestamp 1669390400
transform 1 0 22624 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1650__A2
timestamp 1669390400
transform 1 0 23072 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1651__A1
timestamp 1669390400
transform 1 0 13552 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1651__A2
timestamp 1669390400
transform 1 0 14000 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1652__A1
timestamp 1669390400
transform 1 0 4928 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1652__A2
timestamp 1669390400
transform -1 0 12432 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1652__B
timestamp 1669390400
transform -1 0 13328 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1653__A1
timestamp 1669390400
transform -1 0 11200 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1653__A2
timestamp 1669390400
transform 1 0 12320 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1654__A1
timestamp 1669390400
transform 1 0 17584 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1654__A2
timestamp 1669390400
transform -1 0 18256 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1654__B1
timestamp 1669390400
transform 1 0 16912 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1655__A1
timestamp 1669390400
transform -1 0 20720 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1656__A1
timestamp 1669390400
transform 1 0 21840 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1656__A2
timestamp 1669390400
transform -1 0 21728 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1656__B1
timestamp 1669390400
transform 1 0 22736 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1656__B2
timestamp 1669390400
transform 1 0 21616 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1657__I
timestamp 1669390400
transform -1 0 14336 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1658__A1
timestamp 1669390400
transform -1 0 18928 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1658__A2
timestamp 1669390400
transform 1 0 16464 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1659__I
timestamp 1669390400
transform -1 0 18368 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1660__A1
timestamp 1669390400
transform 1 0 12880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1660__A2
timestamp 1669390400
transform 1 0 14112 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1661__I
timestamp 1669390400
transform 1 0 6496 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1662__I
timestamp 1669390400
transform -1 0 4704 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1663__A1
timestamp 1669390400
transform 1 0 21056 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1663__A2
timestamp 1669390400
transform 1 0 19824 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1664__A1
timestamp 1669390400
transform -1 0 19600 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1665__A1
timestamp 1669390400
transform 1 0 19824 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1665__A2
timestamp 1669390400
transform -1 0 19376 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1665__B1
timestamp 1669390400
transform 1 0 22064 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1665__B2
timestamp 1669390400
transform 1 0 21168 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__A1
timestamp 1669390400
transform 1 0 21952 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__A2
timestamp 1669390400
transform 1 0 23744 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__B1
timestamp 1669390400
transform 1 0 22848 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__B2
timestamp 1669390400
transform 1 0 22400 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1668__A1
timestamp 1669390400
transform 1 0 22288 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1668__A2
timestamp 1669390400
transform -1 0 23408 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1669__A1
timestamp 1669390400
transform 1 0 22064 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1669__A2
timestamp 1669390400
transform 1 0 26768 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1670__A1
timestamp 1669390400
transform 1 0 23632 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1670__A2
timestamp 1669390400
transform 1 0 22512 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1673__I
timestamp 1669390400
transform 1 0 15232 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1674__I
timestamp 1669390400
transform 1 0 2576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1675__I0
timestamp 1669390400
transform 1 0 8960 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1675__I1
timestamp 1669390400
transform 1 0 9632 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1675__S
timestamp 1669390400
transform 1 0 12208 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1676__I
timestamp 1669390400
transform 1 0 3136 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1677__A1
timestamp 1669390400
transform 1 0 21504 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1677__A2
timestamp 1669390400
transform 1 0 20832 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1677__B
timestamp 1669390400
transform 1 0 18592 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1678__A1
timestamp 1669390400
transform 1 0 2688 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1679__A1
timestamp 1669390400
transform 1 0 6720 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1679__A2
timestamp 1669390400
transform -1 0 2352 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1680__A2
timestamp 1669390400
transform -1 0 4144 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1680__B
timestamp 1669390400
transform 1 0 4368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1681__I
timestamp 1669390400
transform 1 0 6720 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1682__A1
timestamp 1669390400
transform -1 0 4816 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1682__A2
timestamp 1669390400
transform 1 0 2016 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1682__B
timestamp 1669390400
transform 1 0 4928 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1682__C
timestamp 1669390400
transform -1 0 2464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1683__I
timestamp 1669390400
transform 1 0 18144 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1684__A2
timestamp 1669390400
transform -1 0 20048 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1684__B
timestamp 1669390400
transform 1 0 19376 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1685__A1
timestamp 1669390400
transform 1 0 6496 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1685__A2
timestamp 1669390400
transform 1 0 6048 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1686__I
timestamp 1669390400
transform 1 0 13552 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1687__A1
timestamp 1669390400
transform 1 0 9968 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1687__A2
timestamp 1669390400
transform 1 0 9968 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1687__B
timestamp 1669390400
transform 1 0 10864 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1688__A1
timestamp 1669390400
transform 1 0 2576 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1688__A2
timestamp 1669390400
transform 1 0 4816 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1688__B
timestamp 1669390400
transform 1 0 4368 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1689__A1
timestamp 1669390400
transform 1 0 18816 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1689__A2
timestamp 1669390400
transform 1 0 17248 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1689__B
timestamp 1669390400
transform 1 0 12880 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1690__A1
timestamp 1669390400
transform 1 0 7616 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1690__A2
timestamp 1669390400
transform 1 0 6720 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1690__A3
timestamp 1669390400
transform 1 0 11312 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1691__A1
timestamp 1669390400
transform -1 0 6384 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1692__A1
timestamp 1669390400
transform 1 0 9632 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1692__A2
timestamp 1669390400
transform 1 0 7168 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1693__A1
timestamp 1669390400
transform 1 0 13552 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1693__A2
timestamp 1669390400
transform 1 0 12320 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1694__A1
timestamp 1669390400
transform 1 0 16912 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1694__A2
timestamp 1669390400
transform 1 0 16912 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1694__A3
timestamp 1669390400
transform 1 0 15568 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1694__B1
timestamp 1669390400
transform -1 0 10304 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1694__B2
timestamp 1669390400
transform 1 0 7616 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1695__A1
timestamp 1669390400
transform 1 0 14896 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1695__A2
timestamp 1669390400
transform 1 0 9632 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1696__A1
timestamp 1669390400
transform 1 0 16800 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1696__B2
timestamp 1669390400
transform 1 0 16464 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1697__A1
timestamp 1669390400
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1697__A2
timestamp 1669390400
transform 1 0 26320 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1697__A3
timestamp 1669390400
transform 1 0 25872 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1698__A1
timestamp 1669390400
transform -1 0 28784 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1698__A2
timestamp 1669390400
transform 1 0 25648 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1698__B
timestamp 1669390400
transform 1 0 30688 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1700__I
timestamp 1669390400
transform -1 0 17136 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1701__A1
timestamp 1669390400
transform 1 0 8624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1701__A2
timestamp 1669390400
transform 1 0 14224 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1701__B
timestamp 1669390400
transform 1 0 7616 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1701__C
timestamp 1669390400
transform 1 0 11312 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1702__A1
timestamp 1669390400
transform 1 0 14336 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1702__A2
timestamp 1669390400
transform 1 0 11984 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1702__C
timestamp 1669390400
transform 1 0 8512 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1703__A1
timestamp 1669390400
transform 1 0 6048 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1703__A2
timestamp 1669390400
transform 1 0 11312 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1703__A3
timestamp 1669390400
transform 1 0 5600 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1704__B
timestamp 1669390400
transform 1 0 4928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1705__A1
timestamp 1669390400
transform -1 0 18928 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1705__A2
timestamp 1669390400
transform 1 0 16352 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1705__B
timestamp 1669390400
transform 1 0 19488 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1706__A1
timestamp 1669390400
transform 1 0 21504 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1708__A1
timestamp 1669390400
transform 1 0 17360 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1708__A2
timestamp 1669390400
transform 1 0 15120 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1708__B
timestamp 1669390400
transform 1 0 16464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1708__C
timestamp 1669390400
transform 1 0 13776 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1709__A1
timestamp 1669390400
transform 1 0 8512 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1709__A2
timestamp 1669390400
transform 1 0 8960 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1709__B
timestamp 1669390400
transform 1 0 10416 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1710__A1
timestamp 1669390400
transform 1 0 13776 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1710__B
timestamp 1669390400
transform 1 0 13888 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1711__A1
timestamp 1669390400
transform 1 0 3920 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1711__A2
timestamp 1669390400
transform 1 0 3472 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1712__A1
timestamp 1669390400
transform 1 0 11984 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1712__A2
timestamp 1669390400
transform 1 0 13888 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1713__I
timestamp 1669390400
transform -1 0 2352 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1714__I
timestamp 1669390400
transform 1 0 2128 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1715__A1
timestamp 1669390400
transform 1 0 13888 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1715__A2
timestamp 1669390400
transform 1 0 7392 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1715__B
timestamp 1669390400
transform 1 0 7840 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1716__A1
timestamp 1669390400
transform -1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1716__A2
timestamp 1669390400
transform 1 0 16464 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1717__C
timestamp 1669390400
transform -1 0 16240 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1718__B
timestamp 1669390400
transform 1 0 20384 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1719__A1
timestamp 1669390400
transform 1 0 22288 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1721__A1
timestamp 1669390400
transform 1 0 23968 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1721__A2
timestamp 1669390400
transform -1 0 24640 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1721__B1
timestamp 1669390400
transform -1 0 23744 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1721__B2
timestamp 1669390400
transform 1 0 23072 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1722__A1
timestamp 1669390400
transform 1 0 27888 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1722__A2
timestamp 1669390400
transform 1 0 26544 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1723__A1
timestamp 1669390400
transform 1 0 4592 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1723__A2
timestamp 1669390400
transform 1 0 4032 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1724__A1
timestamp 1669390400
transform 1 0 4032 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1724__A2
timestamp 1669390400
transform 1 0 3024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1725__A1
timestamp 1669390400
transform 1 0 6608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1725__A2
timestamp 1669390400
transform -1 0 5488 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1726__A1
timestamp 1669390400
transform 1 0 2800 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1726__A2
timestamp 1669390400
transform 1 0 3248 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1726__B
timestamp 1669390400
transform 1 0 2352 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1727__A1
timestamp 1669390400
transform -1 0 1904 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1727__A2
timestamp 1669390400
transform 1 0 4144 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1727__A3
timestamp 1669390400
transform -1 0 4256 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1728__I
timestamp 1669390400
transform 1 0 2688 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1729__I
timestamp 1669390400
transform -1 0 3360 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1730__I0
timestamp 1669390400
transform -1 0 5936 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1730__I1
timestamp 1669390400
transform -1 0 2016 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1731__A1
timestamp 1669390400
transform 1 0 3472 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1731__A2
timestamp 1669390400
transform 1 0 3920 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1731__A3
timestamp 1669390400
transform 1 0 4368 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1732__B
timestamp 1669390400
transform 1 0 3696 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1733__I
timestamp 1669390400
transform -1 0 11984 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1734__A1
timestamp 1669390400
transform 1 0 8064 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1734__A2
timestamp 1669390400
transform 1 0 7168 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1734__A3
timestamp 1669390400
transform 1 0 7616 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1734__B
timestamp 1669390400
transform 1 0 6384 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1735__A1
timestamp 1669390400
transform 1 0 3584 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1735__A2
timestamp 1669390400
transform -1 0 5152 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1736__A1
timestamp 1669390400
transform -1 0 2464 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1737__A1
timestamp 1669390400
transform 1 0 4480 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1737__A2
timestamp 1669390400
transform 1 0 4032 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1738__A1
timestamp 1669390400
transform 1 0 4032 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1738__A2
timestamp 1669390400
transform -1 0 5152 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1739__A1
timestamp 1669390400
transform 1 0 2688 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1739__A2
timestamp 1669390400
transform 1 0 4032 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1740__A1
timestamp 1669390400
transform -1 0 4928 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1740__A2
timestamp 1669390400
transform -1 0 2352 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1741__C
timestamp 1669390400
transform 1 0 5824 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1742__A1
timestamp 1669390400
transform -1 0 26096 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1742__A2
timestamp 1669390400
transform 1 0 25760 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1742__B
timestamp 1669390400
transform -1 0 25088 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1743__A1
timestamp 1669390400
transform 1 0 23184 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1743__A2
timestamp 1669390400
transform -1 0 26544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1743__A3
timestamp 1669390400
transform -1 0 23856 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1745__A1
timestamp 1669390400
transform 1 0 9744 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1745__A2
timestamp 1669390400
transform 1 0 8960 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1745__B1
timestamp 1669390400
transform 1 0 9744 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1745__B2
timestamp 1669390400
transform 1 0 7168 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1745__C
timestamp 1669390400
transform 1 0 14000 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1746__A1
timestamp 1669390400
transform 1 0 7952 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1746__A2
timestamp 1669390400
transform 1 0 12432 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1747__A1
timestamp 1669390400
transform 1 0 10640 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1747__A2
timestamp 1669390400
transform -1 0 10416 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1748__A1
timestamp 1669390400
transform -1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1748__A2
timestamp 1669390400
transform -1 0 12656 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1748__B
timestamp 1669390400
transform 1 0 8288 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1749__B
timestamp 1669390400
transform 1 0 15904 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1750__B
timestamp 1669390400
transform -1 0 5152 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1751__A1
timestamp 1669390400
transform 1 0 4928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1751__A2
timestamp 1669390400
transform -1 0 2016 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1752__A1
timestamp 1669390400
transform 1 0 9632 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1752__A2
timestamp 1669390400
transform 1 0 8960 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1753__A1
timestamp 1669390400
transform 1 0 8064 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1753__A2
timestamp 1669390400
transform 1 0 4928 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1753__A3
timestamp 1669390400
transform -1 0 4704 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1753__B1
timestamp 1669390400
transform -1 0 4704 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1753__B2
timestamp 1669390400
transform 1 0 4928 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1754__A1
timestamp 1669390400
transform 1 0 9632 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1754__A2
timestamp 1669390400
transform 1 0 7616 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1755__A1
timestamp 1669390400
transform 1 0 5936 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1755__A2
timestamp 1669390400
transform -1 0 4704 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1755__B
timestamp 1669390400
transform 1 0 8064 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1756__A1
timestamp 1669390400
transform 1 0 2240 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1756__B
timestamp 1669390400
transform 1 0 3920 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1757__A1
timestamp 1669390400
transform 1 0 6048 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1757__A2
timestamp 1669390400
transform 1 0 5600 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1758__B1
timestamp 1669390400
transform 1 0 6384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1758__B2
timestamp 1669390400
transform -1 0 2576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1758__C
timestamp 1669390400
transform 1 0 8960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1759__A1
timestamp 1669390400
transform -1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1759__C
timestamp 1669390400
transform 1 0 5600 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1760__A1
timestamp 1669390400
transform 1 0 23072 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1760__A2
timestamp 1669390400
transform -1 0 23744 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1760__A3
timestamp 1669390400
transform 1 0 23520 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1761__A1
timestamp 1669390400
transform 1 0 24416 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1761__A2
timestamp 1669390400
transform 1 0 23968 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1761__B
timestamp 1669390400
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1763__A1
timestamp 1669390400
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1763__A2
timestamp 1669390400
transform 1 0 32592 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1763__B1
timestamp 1669390400
transform -1 0 25088 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1763__B2
timestamp 1669390400
transform 1 0 28336 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1764__I
timestamp 1669390400
transform 1 0 31808 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1766__A1
timestamp 1669390400
transform 1 0 23856 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1766__A2
timestamp 1669390400
transform 1 0 28336 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1767__A1
timestamp 1669390400
transform 1 0 36176 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1767__A2
timestamp 1669390400
transform -1 0 28112 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1770__A1
timestamp 1669390400
transform -1 0 6944 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1770__A2
timestamp 1669390400
transform -1 0 7392 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1770__B
timestamp 1669390400
transform -1 0 7840 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1771__A1
timestamp 1669390400
transform -1 0 3696 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1771__A2
timestamp 1669390400
transform 1 0 3920 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1772__A1
timestamp 1669390400
transform -1 0 4256 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1772__A2
timestamp 1669390400
transform -1 0 2576 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1772__B
timestamp 1669390400
transform -1 0 4704 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1773__A1
timestamp 1669390400
transform -1 0 2464 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1774__A1
timestamp 1669390400
transform -1 0 7616 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1774__A2
timestamp 1669390400
transform 1 0 8064 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1774__A3
timestamp 1669390400
transform 1 0 7168 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1775__A1
timestamp 1669390400
transform -1 0 8288 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1775__A2
timestamp 1669390400
transform -1 0 6944 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1775__B1
timestamp 1669390400
transform -1 0 6496 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1775__B2
timestamp 1669390400
transform -1 0 6048 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1775__C
timestamp 1669390400
transform 1 0 4928 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1776__A1
timestamp 1669390400
transform 1 0 4928 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1776__A2
timestamp 1669390400
transform -1 0 2464 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1776__B
timestamp 1669390400
transform 1 0 4480 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1777__I
timestamp 1669390400
transform 1 0 10864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1778__A1
timestamp 1669390400
transform 1 0 13440 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1778__A2
timestamp 1669390400
transform 1 0 9632 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1779__A1
timestamp 1669390400
transform 1 0 9856 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1779__A2
timestamp 1669390400
transform -1 0 12432 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1780__A1
timestamp 1669390400
transform -1 0 9184 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1780__A2
timestamp 1669390400
transform -1 0 5040 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1781__A1
timestamp 1669390400
transform -1 0 6496 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1781__C
timestamp 1669390400
transform -1 0 6832 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1782__A1
timestamp 1669390400
transform 1 0 9184 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1782__A2
timestamp 1669390400
transform 1 0 8960 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1782__B
timestamp 1669390400
transform 1 0 11200 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1783__A1
timestamp 1669390400
transform 1 0 9408 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1783__A2
timestamp 1669390400
transform -1 0 7392 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1783__B1
timestamp 1669390400
transform -1 0 6944 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1783__C
timestamp 1669390400
transform -1 0 9856 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1784__A1
timestamp 1669390400
transform -1 0 7728 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1785__A1
timestamp 1669390400
transform 1 0 9632 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1786__A1
timestamp 1669390400
transform 1 0 28336 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1786__A2
timestamp 1669390400
transform 1 0 22848 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1787__A1
timestamp 1669390400
transform 1 0 8736 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1787__A2
timestamp 1669390400
transform -1 0 10080 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1787__B1
timestamp 1669390400
transform -1 0 10640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1787__B2
timestamp 1669390400
transform 1 0 2352 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1787__C
timestamp 1669390400
transform 1 0 11536 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1788__A1
timestamp 1669390400
transform 1 0 3136 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1788__A2
timestamp 1669390400
transform -1 0 11088 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1788__A3
timestamp 1669390400
transform -1 0 10640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1789__A1
timestamp 1669390400
transform 1 0 3472 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1789__A2
timestamp 1669390400
transform 1 0 7056 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1789__B1
timestamp 1669390400
transform -1 0 6832 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1789__B2
timestamp 1669390400
transform 1 0 4480 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1789__C
timestamp 1669390400
transform 1 0 1792 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1790__B
timestamp 1669390400
transform -1 0 12656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1791__A1
timestamp 1669390400
transform 1 0 3248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1791__A2
timestamp 1669390400
transform 1 0 3696 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1792__A1
timestamp 1669390400
transform 1 0 4144 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1792__A2
timestamp 1669390400
transform 1 0 5936 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1792__A3
timestamp 1669390400
transform 1 0 6384 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1793__A1
timestamp 1669390400
transform -1 0 2912 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1793__A2
timestamp 1669390400
transform -1 0 5936 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1793__C
timestamp 1669390400
transform -1 0 2464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1794__A1
timestamp 1669390400
transform 1 0 7504 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1794__A2
timestamp 1669390400
transform -1 0 10752 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1794__B
timestamp 1669390400
transform -1 0 12656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1795__I0
timestamp 1669390400
transform -1 0 9856 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1795__I1
timestamp 1669390400
transform 1 0 2688 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1796__B
timestamp 1669390400
transform -1 0 10304 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1797__B1
timestamp 1669390400
transform -1 0 9072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1798__A1
timestamp 1669390400
transform -1 0 19152 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1799__I
timestamp 1669390400
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1800__A1
timestamp 1669390400
transform 1 0 16464 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1800__A2
timestamp 1669390400
transform 1 0 15456 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1800__B
timestamp 1669390400
transform 1 0 12880 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1801__A1
timestamp 1669390400
transform 1 0 18144 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1801__B
timestamp 1669390400
transform 1 0 16016 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1802__A1
timestamp 1669390400
transform 1 0 4480 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1802__A2
timestamp 1669390400
transform -1 0 3920 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1802__B
timestamp 1669390400
transform 1 0 8176 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1803__A1
timestamp 1669390400
transform -1 0 17136 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1803__A2
timestamp 1669390400
transform -1 0 16688 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1804__A1
timestamp 1669390400
transform 1 0 8736 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1804__A2
timestamp 1669390400
transform 1 0 7168 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1804__B
timestamp 1669390400
transform 1 0 14336 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1805__A1
timestamp 1669390400
transform 1 0 16912 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1805__A2
timestamp 1669390400
transform 1 0 16912 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1806__A1
timestamp 1669390400
transform 1 0 17584 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1806__A2
timestamp 1669390400
transform 1 0 18032 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1806__B1
timestamp 1669390400
transform 1 0 17136 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1806__C
timestamp 1669390400
transform 1 0 17584 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1807__I
timestamp 1669390400
transform 1 0 17920 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1808__A1
timestamp 1669390400
transform -1 0 16688 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1808__B
timestamp 1669390400
transform -1 0 16240 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1808__C
timestamp 1669390400
transform 1 0 12096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1809__A1
timestamp 1669390400
transform 1 0 19712 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1809__A3
timestamp 1669390400
transform 1 0 18368 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1810__A1
timestamp 1669390400
transform 1 0 19936 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1810__B
timestamp 1669390400
transform 1 0 20384 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1811__A1
timestamp 1669390400
transform 1 0 19376 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1811__A2
timestamp 1669390400
transform 1 0 21504 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1811__B
timestamp 1669390400
transform 1 0 19152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1813__A1
timestamp 1669390400
transform 1 0 19600 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1813__A2
timestamp 1669390400
transform -1 0 20608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1813__A3
timestamp 1669390400
transform 1 0 23632 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1814__A1
timestamp 1669390400
transform 1 0 23184 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1814__A2
timestamp 1669390400
transform -1 0 17808 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1814__B
timestamp 1669390400
transform 1 0 18256 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1815__A2
timestamp 1669390400
transform -1 0 28560 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1816__A1
timestamp 1669390400
transform 1 0 4928 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1816__A2
timestamp 1669390400
transform -1 0 2128 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1816__B
timestamp 1669390400
transform -1 0 2240 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1817__A1
timestamp 1669390400
transform -1 0 2128 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1817__B
timestamp 1669390400
transform -1 0 2464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1818__A1
timestamp 1669390400
transform 1 0 5824 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1818__A2
timestamp 1669390400
transform 1 0 5264 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1819__A1
timestamp 1669390400
transform 1 0 3136 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1819__A2
timestamp 1669390400
transform 1 0 2688 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1819__B
timestamp 1669390400
transform 1 0 5600 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1820__A1
timestamp 1669390400
transform -1 0 8512 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1820__B1
timestamp 1669390400
transform 1 0 4480 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1820__C
timestamp 1669390400
transform 1 0 7840 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1821__B
timestamp 1669390400
transform 1 0 5824 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1822__A1
timestamp 1669390400
transform 1 0 12992 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1822__A2
timestamp 1669390400
transform 1 0 14224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1823__A1
timestamp 1669390400
transform -1 0 9072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1824__A1
timestamp 1669390400
transform 1 0 9632 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1824__A2
timestamp 1669390400
transform -1 0 2016 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1824__B
timestamp 1669390400
transform 1 0 10080 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1825__A1
timestamp 1669390400
transform -1 0 13216 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1825__A2
timestamp 1669390400
transform -1 0 12768 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1825__B1
timestamp 1669390400
transform 1 0 12880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1825__B2
timestamp 1669390400
transform -1 0 12656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1826__A1
timestamp 1669390400
transform 1 0 8960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1826__A2
timestamp 1669390400
transform 1 0 5936 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1826__B
timestamp 1669390400
transform 1 0 8400 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1827__A1
timestamp 1669390400
transform 1 0 13216 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1827__A2
timestamp 1669390400
transform -1 0 13888 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1827__B
timestamp 1669390400
transform -1 0 18816 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1827__C
timestamp 1669390400
transform 1 0 10416 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1828__A1
timestamp 1669390400
transform 1 0 12096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1828__C
timestamp 1669390400
transform -1 0 13776 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1829__A1
timestamp 1669390400
transform -1 0 21056 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1829__A2
timestamp 1669390400
transform -1 0 22848 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1829__A3
timestamp 1669390400
transform -1 0 22400 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1830__A1
timestamp 1669390400
transform -1 0 24640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1830__A2
timestamp 1669390400
transform 1 0 22400 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1830__B
timestamp 1669390400
transform -1 0 23744 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1832__I
timestamp 1669390400
transform 1 0 24304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1833__I
timestamp 1669390400
transform 1 0 28336 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1834__A2
timestamp 1669390400
transform -1 0 29456 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1835__I
timestamp 1669390400
transform 1 0 31024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1836__A1
timestamp 1669390400
transform 1 0 15568 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1837__A1
timestamp 1669390400
transform 1 0 19376 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1837__A2
timestamp 1669390400
transform 1 0 20160 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1837__B
timestamp 1669390400
transform 1 0 18704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1837__C
timestamp 1669390400
transform 1 0 20384 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1838__A1
timestamp 1669390400
transform -1 0 18816 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1838__B
timestamp 1669390400
transform 1 0 19040 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1839__A1
timestamp 1669390400
transform -1 0 16016 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1839__A2
timestamp 1669390400
transform 1 0 8960 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1840__A1
timestamp 1669390400
transform 1 0 13216 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1840__A2
timestamp 1669390400
transform 1 0 13664 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1840__A3
timestamp 1669390400
transform -1 0 11984 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1840__B
timestamp 1669390400
transform 1 0 12208 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1841__A1
timestamp 1669390400
transform 1 0 17136 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1841__A2
timestamp 1669390400
transform 1 0 16912 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1842__A1
timestamp 1669390400
transform 1 0 11984 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1842__A2
timestamp 1669390400
transform 1 0 11536 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1842__A3
timestamp 1669390400
transform 1 0 13552 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1843__A1
timestamp 1669390400
transform 1 0 6496 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1843__A2
timestamp 1669390400
transform -1 0 8288 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1844__A1
timestamp 1669390400
transform -1 0 2016 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1844__A2
timestamp 1669390400
transform -1 0 2912 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1845__A2
timestamp 1669390400
transform 1 0 7616 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1845__B1
timestamp 1669390400
transform -1 0 7168 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1846__A1
timestamp 1669390400
transform 1 0 5824 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1846__A2
timestamp 1669390400
transform 1 0 15568 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1847__A1
timestamp 1669390400
transform -1 0 15232 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1847__B1
timestamp 1669390400
transform 1 0 12880 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1847__B2
timestamp 1669390400
transform 1 0 12096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1848__A1
timestamp 1669390400
transform 1 0 22624 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1848__A3
timestamp 1669390400
transform 1 0 22848 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1849__A2
timestamp 1669390400
transform 1 0 23968 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1849__B
timestamp 1669390400
transform 1 0 24416 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1851__A2
timestamp 1669390400
transform 1 0 31808 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1852__A1
timestamp 1669390400
transform 1 0 9856 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1852__A2
timestamp 1669390400
transform 1 0 8512 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1853__A1
timestamp 1669390400
transform 1 0 11536 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1853__A2
timestamp 1669390400
transform 1 0 9184 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1853__B2
timestamp 1669390400
transform 1 0 11984 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1853__C
timestamp 1669390400
transform 1 0 12432 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1854__A1
timestamp 1669390400
transform 1 0 12432 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1854__A2
timestamp 1669390400
transform 1 0 11984 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1854__C
timestamp 1669390400
transform 1 0 15792 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1855__B
timestamp 1669390400
transform -1 0 18368 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1856__A1
timestamp 1669390400
transform 1 0 10304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1856__A2
timestamp 1669390400
transform -1 0 6160 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1856__A3
timestamp 1669390400
transform 1 0 9744 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1857__B
timestamp 1669390400
transform 1 0 5488 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1858__A2
timestamp 1669390400
transform 1 0 17472 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1858__B
timestamp 1669390400
transform 1 0 17920 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1859__A1
timestamp 1669390400
transform -1 0 18928 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1859__A2
timestamp 1669390400
transform 1 0 17696 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1860__A1
timestamp 1669390400
transform 1 0 16800 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1860__C
timestamp 1669390400
transform 1 0 17808 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1861__A1
timestamp 1669390400
transform -1 0 25088 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1862__B
timestamp 1669390400
transform 1 0 24976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1863__A1
timestamp 1669390400
transform 1 0 27888 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1863__A2
timestamp 1669390400
transform -1 0 27664 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1864__A1
timestamp 1669390400
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1864__A2
timestamp 1669390400
transform 1 0 30016 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1866__A1
timestamp 1669390400
transform 1 0 12656 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1866__A2
timestamp 1669390400
transform 1 0 11424 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1866__B1
timestamp 1669390400
transform -1 0 11200 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1866__B2
timestamp 1669390400
transform 1 0 11760 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1866__C
timestamp 1669390400
transform 1 0 10864 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1867__A1
timestamp 1669390400
transform -1 0 2016 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1867__A2
timestamp 1669390400
transform 1 0 2688 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1867__B
timestamp 1669390400
transform -1 0 2016 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1868__A1
timestamp 1669390400
transform -1 0 8288 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1868__A2
timestamp 1669390400
transform 1 0 12208 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1868__C
timestamp 1669390400
transform 1 0 11760 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1870__A1
timestamp 1669390400
transform 1 0 1904 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1870__A2
timestamp 1669390400
transform 1 0 3584 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1871__A1
timestamp 1669390400
transform -1 0 17472 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1871__A2
timestamp 1669390400
transform -1 0 17024 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1871__B
timestamp 1669390400
transform -1 0 12656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1871__C
timestamp 1669390400
transform 1 0 16128 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1872__A1
timestamp 1669390400
transform 1 0 18928 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1872__A2
timestamp 1669390400
transform 1 0 18480 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1872__B
timestamp 1669390400
transform 1 0 18032 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1872__C
timestamp 1669390400
transform -1 0 18704 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1873__A1
timestamp 1669390400
transform 1 0 17696 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1873__A3
timestamp 1669390400
transform 1 0 20160 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1874__A1
timestamp 1669390400
transform 1 0 20048 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1874__A2
timestamp 1669390400
transform 1 0 16688 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1874__A3
timestamp 1669390400
transform 1 0 19600 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1874__B
timestamp 1669390400
transform 1 0 17584 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1875__A1
timestamp 1669390400
transform 1 0 18480 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1875__A2
timestamp 1669390400
transform -1 0 18256 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1876__A1
timestamp 1669390400
transform -1 0 24528 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1876__A2
timestamp 1669390400
transform -1 0 25088 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1877__A1
timestamp 1669390400
transform 1 0 27552 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1877__A2
timestamp 1669390400
transform -1 0 29008 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1877__B
timestamp 1669390400
transform 1 0 28000 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1877__C
timestamp 1669390400
transform 1 0 28336 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1878__A2
timestamp 1669390400
transform -1 0 28112 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1880__A2
timestamp 1669390400
transform -1 0 31136 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1881__A1
timestamp 1669390400
transform 1 0 28336 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1881__B1
timestamp 1669390400
transform 1 0 32704 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1881__B2
timestamp 1669390400
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1882__A1
timestamp 1669390400
transform 1 0 10304 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1882__A2
timestamp 1669390400
transform 1 0 8064 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1882__B
timestamp 1669390400
transform 1 0 7616 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1883__A1
timestamp 1669390400
transform 1 0 7616 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1883__A2
timestamp 1669390400
transform 1 0 4816 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1883__B2
timestamp 1669390400
transform 1 0 10080 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1883__C
timestamp 1669390400
transform 1 0 8512 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1884__A1
timestamp 1669390400
transform 1 0 5040 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1884__A2
timestamp 1669390400
transform 1 0 6048 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1884__B
timestamp 1669390400
transform -1 0 2016 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1885__A2
timestamp 1669390400
transform -1 0 8960 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1885__B1
timestamp 1669390400
transform -1 0 9184 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1885__B2
timestamp 1669390400
transform 1 0 9408 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1885__C
timestamp 1669390400
transform 1 0 4928 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1886__B
timestamp 1669390400
transform -1 0 2688 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1887__I0
timestamp 1669390400
transform -1 0 2240 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1887__I1
timestamp 1669390400
transform -1 0 2016 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1887__S
timestamp 1669390400
transform -1 0 1904 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1888__A1
timestamp 1669390400
transform 1 0 10080 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1888__A2
timestamp 1669390400
transform 1 0 10304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1888__B
timestamp 1669390400
transform 1 0 10640 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1889__A1
timestamp 1669390400
transform 1 0 9744 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1889__A2
timestamp 1669390400
transform 1 0 12432 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1889__B1
timestamp 1669390400
transform 1 0 16016 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1889__B2
timestamp 1669390400
transform 1 0 17808 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1889__C
timestamp 1669390400
transform 1 0 19936 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1890__A1
timestamp 1669390400
transform -1 0 17808 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1890__C
timestamp 1669390400
transform 1 0 19152 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1891__A1
timestamp 1669390400
transform 1 0 25984 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1891__A2
timestamp 1669390400
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1891__A3
timestamp 1669390400
transform 1 0 24416 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1892__A1
timestamp 1669390400
transform -1 0 25648 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1892__A2
timestamp 1669390400
transform -1 0 26880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1892__B
timestamp 1669390400
transform 1 0 23968 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1894__A1
timestamp 1669390400
transform 1 0 28560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1894__A2
timestamp 1669390400
transform -1 0 28224 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1894__B1
timestamp 1669390400
transform -1 0 23184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1894__B2
timestamp 1669390400
transform 1 0 23744 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1895__A1
timestamp 1669390400
transform 1 0 26320 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1895__A2
timestamp 1669390400
transform -1 0 26880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1896__I
timestamp 1669390400
transform 1 0 19936 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1897__A1
timestamp 1669390400
transform 1 0 27440 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1897__A2
timestamp 1669390400
transform -1 0 28112 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1898__B1
timestamp 1669390400
transform -1 0 28336 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1898__B2
timestamp 1669390400
transform 1 0 25648 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1899__A1
timestamp 1669390400
transform 1 0 24416 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1899__A2
timestamp 1669390400
transform -1 0 24976 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1899__B1
timestamp 1669390400
transform -1 0 26320 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1899__B2
timestamp 1669390400
transform 1 0 25648 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1900__A1
timestamp 1669390400
transform 1 0 22736 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1900__A2
timestamp 1669390400
transform -1 0 25088 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1900__B1
timestamp 1669390400
transform 1 0 26096 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1900__B2
timestamp 1669390400
transform 1 0 26320 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1901__A1
timestamp 1669390400
transform 1 0 25760 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1901__A2
timestamp 1669390400
transform 1 0 23184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1902__A2
timestamp 1669390400
transform -1 0 23632 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1905__I
timestamp 1669390400
transform -1 0 3808 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1906__I
timestamp 1669390400
transform -1 0 16688 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1907__A1
timestamp 1669390400
transform -1 0 16688 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1907__A2
timestamp 1669390400
transform -1 0 16688 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1909__A1
timestamp 1669390400
transform -1 0 16240 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1910__A1
timestamp 1669390400
transform 1 0 8512 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1910__A2
timestamp 1669390400
transform 1 0 8960 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1911__A1
timestamp 1669390400
transform -1 0 6496 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1912__A1
timestamp 1669390400
transform 1 0 12096 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1913__A1
timestamp 1669390400
transform -1 0 17696 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1914__A1
timestamp 1669390400
transform -1 0 14112 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1915__A1
timestamp 1669390400
transform -1 0 13664 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1915__B2
timestamp 1669390400
transform -1 0 7392 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1916__A1
timestamp 1669390400
transform -1 0 12880 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1917__A1
timestamp 1669390400
transform 1 0 24080 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1917__A2
timestamp 1669390400
transform 1 0 20160 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1917__B1
timestamp 1669390400
transform 1 0 25536 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1917__B2
timestamp 1669390400
transform 1 0 24528 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1918__A1
timestamp 1669390400
transform 1 0 16016 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1919__A1
timestamp 1669390400
transform -1 0 19264 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1920__A1
timestamp 1669390400
transform -1 0 20832 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1921__A1
timestamp 1669390400
transform 1 0 20944 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1921__A2
timestamp 1669390400
transform 1 0 21728 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1921__B1
timestamp 1669390400
transform 1 0 22176 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1921__B2
timestamp 1669390400
transform 1 0 21392 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1922__A1
timestamp 1669390400
transform -1 0 15792 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1923__A1
timestamp 1669390400
transform -1 0 18144 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1924__A1
timestamp 1669390400
transform -1 0 21056 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1924__A2
timestamp 1669390400
transform 1 0 20944 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1924__B1
timestamp 1669390400
transform 1 0 21392 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1924__B2
timestamp 1669390400
transform -1 0 19936 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1926__A1
timestamp 1669390400
transform 1 0 21840 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1926__A2
timestamp 1669390400
transform 1 0 22288 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1927__A1
timestamp 1669390400
transform 1 0 5040 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1928__A1
timestamp 1669390400
transform 1 0 6048 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1928__A2
timestamp 1669390400
transform 1 0 6496 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1929__A1
timestamp 1669390400
transform 1 0 8960 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1930__A1
timestamp 1669390400
transform 1 0 2240 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1930__A2
timestamp 1669390400
transform 1 0 2352 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1930__B
timestamp 1669390400
transform 1 0 4816 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1931__A1
timestamp 1669390400
transform -1 0 2240 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1931__A2
timestamp 1669390400
transform -1 0 5152 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1931__A3
timestamp 1669390400
transform -1 0 2016 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1931__B1
timestamp 1669390400
transform -1 0 9856 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1931__B2
timestamp 1669390400
transform -1 0 1904 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1932__A1
timestamp 1669390400
transform 1 0 2912 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1932__A2
timestamp 1669390400
transform -1 0 4368 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1932__B
timestamp 1669390400
transform 1 0 4480 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1933__A1
timestamp 1669390400
transform 1 0 5712 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1933__A2
timestamp 1669390400
transform 1 0 2800 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1933__B
timestamp 1669390400
transform -1 0 3360 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1934__A1
timestamp 1669390400
transform -1 0 2128 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1934__C
timestamp 1669390400
transform -1 0 2352 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1935__A1
timestamp 1669390400
transform -1 0 11312 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1936__A1
timestamp 1669390400
transform -1 0 21056 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1937__A1
timestamp 1669390400
transform -1 0 11424 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1937__A2
timestamp 1669390400
transform 1 0 11648 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1937__B
timestamp 1669390400
transform 1 0 12096 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1938__A2
timestamp 1669390400
transform -1 0 10976 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1938__B
timestamp 1669390400
transform -1 0 14560 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1939__A1
timestamp 1669390400
transform 1 0 3584 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1939__A2
timestamp 1669390400
transform 1 0 3136 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1940__A1
timestamp 1669390400
transform 1 0 6384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1940__A2
timestamp 1669390400
transform 1 0 2352 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1940__B1
timestamp 1669390400
transform 1 0 4032 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1940__B2
timestamp 1669390400
transform 1 0 9856 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1940__C
timestamp 1669390400
transform 1 0 5600 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1941__A1
timestamp 1669390400
transform -1 0 16128 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1941__A3
timestamp 1669390400
transform 1 0 15456 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1942__A1
timestamp 1669390400
transform 1 0 8512 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1942__A2
timestamp 1669390400
transform 1 0 7616 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1943__A1
timestamp 1669390400
transform 1 0 12544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1943__A2
timestamp 1669390400
transform 1 0 12992 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1943__B
timestamp 1669390400
transform 1 0 15456 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1944__A2
timestamp 1669390400
transform 1 0 15120 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1945__A1
timestamp 1669390400
transform 1 0 16016 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1945__B2
timestamp 1669390400
transform 1 0 12432 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1946__A1
timestamp 1669390400
transform 1 0 16912 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1947__A1
timestamp 1669390400
transform 1 0 22848 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1948__A1
timestamp 1669390400
transform 1 0 21504 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1948__A2
timestamp 1669390400
transform 1 0 25648 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1948__B1
timestamp 1669390400
transform -1 0 26096 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1948__B2
timestamp 1669390400
transform 1 0 24416 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1949__A1
timestamp 1669390400
transform 1 0 9184 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1949__A2
timestamp 1669390400
transform 1 0 8288 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1950__A1
timestamp 1669390400
transform 1 0 12432 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1950__A2
timestamp 1669390400
transform 1 0 12880 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1950__B
timestamp 1669390400
transform 1 0 12432 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1951__A1
timestamp 1669390400
transform 1 0 6720 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1951__A2
timestamp 1669390400
transform 1 0 6272 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1952__A1
timestamp 1669390400
transform -1 0 5152 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1953__A1
timestamp 1669390400
transform -1 0 5600 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1953__B2
timestamp 1669390400
transform -1 0 6048 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1954__A1
timestamp 1669390400
transform 1 0 19264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1954__A2
timestamp 1669390400
transform 1 0 15568 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1954__C
timestamp 1669390400
transform 1 0 16912 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1955__A1
timestamp 1669390400
transform 1 0 4144 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1955__B1
timestamp 1669390400
transform -1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1955__B2
timestamp 1669390400
transform 1 0 13104 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1956__A1
timestamp 1669390400
transform 1 0 11424 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1957__A1
timestamp 1669390400
transform 1 0 19264 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1958__A1
timestamp 1669390400
transform 1 0 19936 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1959__A1
timestamp 1669390400
transform 1 0 3584 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1959__A2
timestamp 1669390400
transform -1 0 2016 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1959__B
timestamp 1669390400
transform -1 0 4928 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1960__A1
timestamp 1669390400
transform -1 0 2016 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1960__B
timestamp 1669390400
transform 1 0 3024 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1961__A1
timestamp 1669390400
transform 1 0 2240 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1961__A2
timestamp 1669390400
transform -1 0 2688 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1962__A1
timestamp 1669390400
transform 1 0 2688 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1962__A2
timestamp 1669390400
transform -1 0 5712 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1962__B1
timestamp 1669390400
transform 1 0 3136 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1962__B2
timestamp 1669390400
transform -1 0 2128 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1962__C
timestamp 1669390400
transform 1 0 4144 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1963__A1
timestamp 1669390400
transform -1 0 3808 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1964__A1
timestamp 1669390400
transform -1 0 2912 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1964__A2
timestamp 1669390400
transform -1 0 2128 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1965__A1
timestamp 1669390400
transform -1 0 3808 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1965__B1
timestamp 1669390400
transform -1 0 1904 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1965__B2
timestamp 1669390400
transform -1 0 4704 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1965__C
timestamp 1669390400
transform 1 0 2352 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1966__A1
timestamp 1669390400
transform -1 0 2240 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1966__A2
timestamp 1669390400
transform 1 0 4032 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1966__A3
timestamp 1669390400
transform -1 0 3024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1966__B
timestamp 1669390400
transform -1 0 2464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1968__A1
timestamp 1669390400
transform 1 0 23520 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1968__A2
timestamp 1669390400
transform 1 0 23072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1969__A1
timestamp 1669390400
transform 1 0 2576 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1969__A2
timestamp 1669390400
transform 1 0 3472 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1970__A1
timestamp 1669390400
transform -1 0 4032 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1970__A2
timestamp 1669390400
transform 1 0 4256 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1971__A1
timestamp 1669390400
transform 1 0 5600 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1971__A2
timestamp 1669390400
transform 1 0 4816 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1972__A1
timestamp 1669390400
transform 1 0 6048 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1972__A2
timestamp 1669390400
transform -1 0 2352 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1972__B
timestamp 1669390400
transform 1 0 5712 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1973__A1
timestamp 1669390400
transform 1 0 5712 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1973__A2
timestamp 1669390400
transform -1 0 2016 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1973__B1
timestamp 1669390400
transform -1 0 2464 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1973__B2
timestamp 1669390400
transform -1 0 2016 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1973__C
timestamp 1669390400
transform 1 0 6944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1974__C
timestamp 1669390400
transform 1 0 9184 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1975__A1
timestamp 1669390400
transform -1 0 5152 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1976__A1
timestamp 1669390400
transform 1 0 22176 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1976__A2
timestamp 1669390400
transform -1 0 19152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1977__A1
timestamp 1669390400
transform -1 0 3024 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1977__A2
timestamp 1669390400
transform -1 0 3472 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1978__A1
timestamp 1669390400
transform -1 0 2016 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1978__A2
timestamp 1669390400
transform -1 0 2912 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1979__B
timestamp 1669390400
transform -1 0 3808 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1979__C
timestamp 1669390400
transform -1 0 4592 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1980__A1
timestamp 1669390400
transform -1 0 8736 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1980__A2
timestamp 1669390400
transform -1 0 6160 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1980__B
timestamp 1669390400
transform -1 0 7952 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1981__A1
timestamp 1669390400
transform -1 0 8736 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1981__A2
timestamp 1669390400
transform 1 0 5264 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1981__C
timestamp 1669390400
transform -1 0 7056 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1982__A1
timestamp 1669390400
transform 1 0 10528 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1982__A2
timestamp 1669390400
transform 1 0 8512 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1982__B1
timestamp 1669390400
transform -1 0 10304 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1982__C
timestamp 1669390400
transform -1 0 9632 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1983__A1
timestamp 1669390400
transform -1 0 10080 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1983__B
timestamp 1669390400
transform -1 0 5152 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1983__C
timestamp 1669390400
transform 1 0 5376 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1984__A1
timestamp 1669390400
transform 1 0 8736 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1986__A1
timestamp 1669390400
transform 1 0 22624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1986__A2
timestamp 1669390400
transform 1 0 22176 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1987__A1
timestamp 1669390400
transform -1 0 2016 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1987__A2
timestamp 1669390400
transform -1 0 2128 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1987__B1
timestamp 1669390400
transform -1 0 3024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1988__A1
timestamp 1669390400
transform -1 0 10752 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1988__A2
timestamp 1669390400
transform -1 0 10304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1988__B
timestamp 1669390400
transform -1 0 1904 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1989__A1
timestamp 1669390400
transform 1 0 3024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1989__B
timestamp 1669390400
transform 1 0 7952 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1990__A1
timestamp 1669390400
transform -1 0 10192 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1990__A2
timestamp 1669390400
transform -1 0 11536 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1990__B2
timestamp 1669390400
transform -1 0 10640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1991__A1
timestamp 1669390400
transform -1 0 11088 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1991__B2
timestamp 1669390400
transform -1 0 11536 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1991__C
timestamp 1669390400
transform 1 0 11760 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1992__A1
timestamp 1669390400
transform -1 0 5152 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1992__A2
timestamp 1669390400
transform 1 0 5152 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1992__B1
timestamp 1669390400
transform 1 0 8288 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1992__B2
timestamp 1669390400
transform 1 0 8736 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1993__A1
timestamp 1669390400
transform 1 0 8624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1994__A1
timestamp 1669390400
transform -1 0 5936 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1994__A2
timestamp 1669390400
transform -1 0 10416 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1994__A3
timestamp 1669390400
transform -1 0 5152 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1994__A4
timestamp 1669390400
transform -1 0 14560 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1996__A1
timestamp 1669390400
transform 1 0 18256 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1997__A1
timestamp 1669390400
transform 1 0 5376 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1998__A1
timestamp 1669390400
transform 1 0 8176 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1998__A2
timestamp 1669390400
transform 1 0 3024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1999__I0
timestamp 1669390400
transform 1 0 4032 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1999__I1
timestamp 1669390400
transform -1 0 4592 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2000__A2
timestamp 1669390400
transform -1 0 4704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2000__B1
timestamp 1669390400
transform -1 0 7504 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2000__B2
timestamp 1669390400
transform 1 0 5824 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2001__B2
timestamp 1669390400
transform -1 0 4704 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2002__A1
timestamp 1669390400
transform -1 0 5600 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2002__A2
timestamp 1669390400
transform -1 0 1904 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2002__B
timestamp 1669390400
transform 1 0 3024 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2003__A1
timestamp 1669390400
transform 1 0 5376 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2003__A2
timestamp 1669390400
transform -1 0 6496 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2003__A3
timestamp 1669390400
transform -1 0 3248 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2003__A4
timestamp 1669390400
transform -1 0 5152 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2004__A2
timestamp 1669390400
transform -1 0 1904 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2004__B
timestamp 1669390400
transform 1 0 6272 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2005__A1
timestamp 1669390400
transform -1 0 7392 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2005__C
timestamp 1669390400
transform 1 0 7616 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2006__A1
timestamp 1669390400
transform -1 0 6384 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2007__A1
timestamp 1669390400
transform 1 0 22736 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2007__A2
timestamp 1669390400
transform -1 0 23408 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2008__A1
timestamp 1669390400
transform -1 0 15792 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2008__A2
timestamp 1669390400
transform -1 0 13888 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2008__B1
timestamp 1669390400
transform -1 0 12656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2008__B2
timestamp 1669390400
transform 1 0 11760 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2009__A1
timestamp 1669390400
transform -1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2010__A1
timestamp 1669390400
transform -1 0 12208 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2010__B
timestamp 1669390400
transform 1 0 11088 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2011__A1
timestamp 1669390400
transform -1 0 6496 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2011__A2
timestamp 1669390400
transform -1 0 11872 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2011__B
timestamp 1669390400
transform 1 0 11200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2011__C
timestamp 1669390400
transform 1 0 13440 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2012__C
timestamp 1669390400
transform 1 0 8400 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2013__A1
timestamp 1669390400
transform 1 0 15120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2013__A2
timestamp 1669390400
transform -1 0 14112 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2013__A3
timestamp 1669390400
transform -1 0 14896 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2014__A1
timestamp 1669390400
transform 1 0 8400 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2014__A2
timestamp 1669390400
transform 1 0 12544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2014__A3
timestamp 1669390400
transform 1 0 13552 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2014__B
timestamp 1669390400
transform -1 0 14448 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2015__A1
timestamp 1669390400
transform 1 0 14112 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2015__A3
timestamp 1669390400
transform -1 0 15904 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2015__A4
timestamp 1669390400
transform -1 0 14560 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2016__A1
timestamp 1669390400
transform 1 0 18928 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2017__B
timestamp 1669390400
transform 1 0 18480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2018__A1
timestamp 1669390400
transform 1 0 41440 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2018__A2
timestamp 1669390400
transform -1 0 38528 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2019__A1
timestamp 1669390400
transform 1 0 17248 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2020__A1
timestamp 1669390400
transform -1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2020__A2
timestamp 1669390400
transform 1 0 9184 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2020__A3
timestamp 1669390400
transform 1 0 8512 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2021__A1
timestamp 1669390400
transform 1 0 8512 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2021__A2
timestamp 1669390400
transform 1 0 12880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2021__B2
timestamp 1669390400
transform -1 0 9744 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2022__B2
timestamp 1669390400
transform 1 0 12432 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2023__A1
timestamp 1669390400
transform 1 0 20832 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2024__A1
timestamp 1669390400
transform -1 0 17136 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2024__A2
timestamp 1669390400
transform 1 0 21952 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2024__A3
timestamp 1669390400
transform 1 0 16464 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2025__A1
timestamp 1669390400
transform 1 0 14560 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2025__A2
timestamp 1669390400
transform 1 0 12880 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2025__B
timestamp 1669390400
transform 1 0 15344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2026__B
timestamp 1669390400
transform 1 0 20608 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2027__A1
timestamp 1669390400
transform 1 0 20832 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2028__A1
timestamp 1669390400
transform 1 0 19488 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2029__I
timestamp 1669390400
transform 1 0 39312 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2030__I
timestamp 1669390400
transform 1 0 42112 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2031__A1
timestamp 1669390400
transform 1 0 14560 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2031__A2
timestamp 1669390400
transform -1 0 15456 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2031__B1
timestamp 1669390400
transform 1 0 11312 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2031__B2
timestamp 1669390400
transform 1 0 11312 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2032__A1
timestamp 1669390400
transform 1 0 2352 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2032__B
timestamp 1669390400
transform -1 0 15120 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2032__C
timestamp 1669390400
transform -1 0 8064 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2033__A1
timestamp 1669390400
transform -1 0 15008 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2034__A1
timestamp 1669390400
transform -1 0 16240 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2034__A2
timestamp 1669390400
transform -1 0 15792 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2035__A1
timestamp 1669390400
transform 1 0 16464 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2035__A2
timestamp 1669390400
transform 1 0 15120 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2035__B2
timestamp 1669390400
transform 1 0 17360 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2036__A1
timestamp 1669390400
transform 1 0 17808 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2036__A2
timestamp 1669390400
transform 1 0 17584 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2037__A2
timestamp 1669390400
transform 1 0 16016 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2037__B1
timestamp 1669390400
transform 1 0 14784 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2037__C
timestamp 1669390400
transform -1 0 15456 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2038__A1
timestamp 1669390400
transform 1 0 16912 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2038__B2
timestamp 1669390400
transform 1 0 16464 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2039__A1
timestamp 1669390400
transform 1 0 16912 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2039__A2
timestamp 1669390400
transform -1 0 15456 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2040__A1
timestamp 1669390400
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2040__A2
timestamp 1669390400
transform 1 0 31584 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2040__B
timestamp 1669390400
transform -1 0 30464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2040__C
timestamp 1669390400
transform 1 0 30688 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2041__A1
timestamp 1669390400
transform 1 0 4256 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2041__A2
timestamp 1669390400
transform -1 0 3584 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2042__B
timestamp 1669390400
transform 1 0 5824 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2043__A1
timestamp 1669390400
transform -1 0 2128 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2043__A2
timestamp 1669390400
transform 1 0 6272 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2043__A3
timestamp 1669390400
transform 1 0 8064 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2044__A1
timestamp 1669390400
transform 1 0 4480 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2044__C
timestamp 1669390400
transform 1 0 5600 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2045__A1
timestamp 1669390400
transform 1 0 8960 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2045__A2
timestamp 1669390400
transform -1 0 2688 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2045__B1
timestamp 1669390400
transform 1 0 6048 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2045__B2
timestamp 1669390400
transform -1 0 2912 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2045__C
timestamp 1669390400
transform -1 0 9856 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2046__A1
timestamp 1669390400
transform 1 0 2912 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2047__A1
timestamp 1669390400
transform 1 0 6720 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2048__A1
timestamp 1669390400
transform 1 0 16464 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2048__A2
timestamp 1669390400
transform 1 0 16912 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2049__A1
timestamp 1669390400
transform 1 0 28336 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2049__A2
timestamp 1669390400
transform 1 0 32032 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2049__B1
timestamp 1669390400
transform -1 0 31136 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2049__B2
timestamp 1669390400
transform 1 0 29344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2050__A1
timestamp 1669390400
transform 1 0 31136 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2050__A2
timestamp 1669390400
transform 1 0 35616 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2050__B1
timestamp 1669390400
transform 1 0 35168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2050__B2
timestamp 1669390400
transform 1 0 31584 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2052__A1
timestamp 1669390400
transform 1 0 22960 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2052__A2
timestamp 1669390400
transform -1 0 23632 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2052__B1
timestamp 1669390400
transform -1 0 26992 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2052__B2
timestamp 1669390400
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2053__A1
timestamp 1669390400
transform 1 0 25648 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2053__A2
timestamp 1669390400
transform -1 0 28560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2053__B1
timestamp 1669390400
transform -1 0 23072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2053__B2
timestamp 1669390400
transform 1 0 27216 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2054__B1
timestamp 1669390400
transform 1 0 24976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2054__B2
timestamp 1669390400
transform 1 0 25424 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2055__A1
timestamp 1669390400
transform 1 0 26432 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2055__A2
timestamp 1669390400
transform 1 0 25872 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2056__A1
timestamp 1669390400
transform 1 0 21504 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2056__A2
timestamp 1669390400
transform -1 0 23296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2057__A1
timestamp 1669390400
transform -1 0 22176 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2057__A2
timestamp 1669390400
transform -1 0 20608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2058__A1
timestamp 1669390400
transform 1 0 20384 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2058__A2
timestamp 1669390400
transform -1 0 23296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2058__B1
timestamp 1669390400
transform -1 0 23744 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2058__B2
timestamp 1669390400
transform 1 0 20832 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2059__A1
timestamp 1669390400
transform 1 0 24416 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2059__A2
timestamp 1669390400
transform 1 0 25536 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2059__B1
timestamp 1669390400
transform 1 0 23968 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2059__B2
timestamp 1669390400
transform 1 0 22624 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2061__A1
timestamp 1669390400
transform 1 0 20832 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2061__A2
timestamp 1669390400
transform -1 0 23184 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2061__B1
timestamp 1669390400
transform -1 0 22848 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2061__B2
timestamp 1669390400
transform 1 0 22960 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2062__A1
timestamp 1669390400
transform 1 0 24640 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2062__A2
timestamp 1669390400
transform 1 0 23744 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2064__A1
timestamp 1669390400
transform 1 0 23968 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2064__A2
timestamp 1669390400
transform -1 0 25760 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2069__I
timestamp 1669390400
transform 1 0 19376 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2071__A1
timestamp 1669390400
transform -1 0 16464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2071__A2
timestamp 1669390400
transform 1 0 23744 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2071__A3
timestamp 1669390400
transform -1 0 16240 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2072__A1
timestamp 1669390400
transform 1 0 40432 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2072__A2
timestamp 1669390400
transform -1 0 41888 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2073__A1
timestamp 1669390400
transform 1 0 46704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2073__A2
timestamp 1669390400
transform 1 0 46480 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2074__A2
timestamp 1669390400
transform -1 0 21504 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2074__A3
timestamp 1669390400
transform 1 0 17136 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2074__B
timestamp 1669390400
transform -1 0 21056 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2075__I
timestamp 1669390400
transform -1 0 20608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2076__A2
timestamp 1669390400
transform -1 0 18928 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2076__A3
timestamp 1669390400
transform -1 0 19936 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2078__A2
timestamp 1669390400
transform -1 0 19600 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2079__A1
timestamp 1669390400
transform 1 0 47376 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2079__A2
timestamp 1669390400
transform 1 0 45808 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2079__B1
timestamp 1669390400
transform 1 0 46480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2079__B2
timestamp 1669390400
transform 1 0 46928 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2080__A1
timestamp 1669390400
transform 1 0 49280 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2081__A1
timestamp 1669390400
transform -1 0 45584 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2081__A2
timestamp 1669390400
transform 1 0 44912 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2082__A1
timestamp 1669390400
transform 1 0 19936 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2082__A2
timestamp 1669390400
transform 1 0 18704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2084__A1
timestamp 1669390400
transform -1 0 40320 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2084__A2
timestamp 1669390400
transform -1 0 40992 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2085__A1
timestamp 1669390400
transform 1 0 45136 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2085__A2
timestamp 1669390400
transform -1 0 45808 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2086__A1
timestamp 1669390400
transform 1 0 47712 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2087__A1
timestamp 1669390400
transform 1 0 49168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2090__A1
timestamp 1669390400
transform 1 0 52640 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2091__A1
timestamp 1669390400
transform 1 0 23520 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2091__A2
timestamp 1669390400
transform 1 0 23968 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2092__I
timestamp 1669390400
transform -1 0 17136 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2093__A2
timestamp 1669390400
transform 1 0 17808 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2094__I
timestamp 1669390400
transform -1 0 27216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2095__A2
timestamp 1669390400
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2097__A1
timestamp 1669390400
transform -1 0 18928 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2097__A2
timestamp 1669390400
transform -1 0 17136 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2098__A1
timestamp 1669390400
transform -1 0 43120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2098__A2
timestamp 1669390400
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2099__A1
timestamp 1669390400
transform 1 0 19152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2099__A2
timestamp 1669390400
transform 1 0 18032 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2100__A1
timestamp 1669390400
transform -1 0 17136 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2101__A1
timestamp 1669390400
transform 1 0 18480 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2103__I
timestamp 1669390400
transform 1 0 42448 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2104__A1
timestamp 1669390400
transform -1 0 42336 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2104__B
timestamp 1669390400
transform 1 0 42560 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2104__C
timestamp 1669390400
transform 1 0 44240 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2107__A2
timestamp 1669390400
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2108__A3
timestamp 1669390400
transform 1 0 22736 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2110__A1
timestamp 1669390400
transform -1 0 24080 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2110__A2
timestamp 1669390400
transform -1 0 23632 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2110__A3
timestamp 1669390400
transform 1 0 20384 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2111__B
timestamp 1669390400
transform 1 0 28336 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2112__I0
timestamp 1669390400
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2112__I1
timestamp 1669390400
transform 1 0 37408 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2112__S
timestamp 1669390400
transform 1 0 36960 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2113__A1
timestamp 1669390400
transform 1 0 35168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2113__A2
timestamp 1669390400
transform 1 0 34720 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2114__A1
timestamp 1669390400
transform 1 0 38080 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2114__A2
timestamp 1669390400
transform 1 0 35840 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2115__A1
timestamp 1669390400
transform 1 0 43792 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2115__A2
timestamp 1669390400
transform 1 0 43344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2116__A1
timestamp 1669390400
transform 1 0 24416 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2116__A2
timestamp 1669390400
transform 1 0 19488 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2117__A1
timestamp 1669390400
transform 1 0 33488 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2117__A2
timestamp 1669390400
transform 1 0 31696 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2118__A1
timestamp 1669390400
transform -1 0 39648 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2118__A2
timestamp 1669390400
transform 1 0 37072 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2118__B
timestamp 1669390400
transform 1 0 37408 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2123__I
timestamp 1669390400
transform 1 0 48160 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2124__A1
timestamp 1669390400
transform 1 0 45696 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2124__A2
timestamp 1669390400
transform 1 0 48272 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2125__A1
timestamp 1669390400
transform 1 0 45248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2125__A2
timestamp 1669390400
transform -1 0 45584 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2126__A1
timestamp 1669390400
transform -1 0 46144 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2126__B
timestamp 1669390400
transform 1 0 46368 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2127__A1
timestamp 1669390400
transform 1 0 23520 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2127__A2
timestamp 1669390400
transform 1 0 23072 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2128__A2
timestamp 1669390400
transform -1 0 26320 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2129__A1
timestamp 1669390400
transform 1 0 40768 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2129__A2
timestamp 1669390400
transform 1 0 40992 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2129__B1
timestamp 1669390400
transform -1 0 39424 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2129__B2
timestamp 1669390400
transform 1 0 41440 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2130__A1
timestamp 1669390400
transform 1 0 47040 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2130__A2
timestamp 1669390400
transform 1 0 47488 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2132__A1
timestamp 1669390400
transform 1 0 51184 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2133__A1
timestamp 1669390400
transform -1 0 51632 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2134__A1
timestamp 1669390400
transform 1 0 53088 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2136__B
timestamp 1669390400
transform -1 0 29792 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2137__A1
timestamp 1669390400
transform -1 0 36960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2138__A2
timestamp 1669390400
transform 1 0 20832 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2139__A1
timestamp 1669390400
transform 1 0 19824 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2140__A2
timestamp 1669390400
transform 1 0 20048 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2142__A1
timestamp 1669390400
transform 1 0 28336 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2142__A2
timestamp 1669390400
transform 1 0 20832 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2143__A2
timestamp 1669390400
transform -1 0 21056 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2144__A1
timestamp 1669390400
transform 1 0 19152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2147__A1
timestamp 1669390400
transform 1 0 31248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2147__A2
timestamp 1669390400
transform 1 0 31696 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2147__B1
timestamp 1669390400
transform 1 0 32144 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2147__C1
timestamp 1669390400
transform 1 0 29904 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2147__C2
timestamp 1669390400
transform 1 0 30352 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2149__I
timestamp 1669390400
transform -1 0 25872 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2150__A1
timestamp 1669390400
transform -1 0 29904 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2150__A2
timestamp 1669390400
transform 1 0 32928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2151__A1
timestamp 1669390400
transform 1 0 33376 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2151__A2
timestamp 1669390400
transform 1 0 33488 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2152__A1
timestamp 1669390400
transform 1 0 30240 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2152__A2
timestamp 1669390400
transform -1 0 29344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2152__B
timestamp 1669390400
transform 1 0 30800 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2153__A2
timestamp 1669390400
transform -1 0 32480 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2154__A1
timestamp 1669390400
transform 1 0 41216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2154__A2
timestamp 1669390400
transform 1 0 29456 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2154__B1
timestamp 1669390400
transform 1 0 29904 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2154__B2
timestamp 1669390400
transform 1 0 29344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2154__C1
timestamp 1669390400
transform -1 0 25872 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2156__A1
timestamp 1669390400
transform 1 0 44688 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2156__A2
timestamp 1669390400
transform -1 0 44128 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2158__A1
timestamp 1669390400
transform 1 0 45472 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2158__A2
timestamp 1669390400
transform -1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2160__A3
timestamp 1669390400
transform 1 0 32480 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2161__A2
timestamp 1669390400
transform 1 0 29792 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2163__A1
timestamp 1669390400
transform 1 0 34496 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2163__A2
timestamp 1669390400
transform 1 0 33488 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2165__B
timestamp 1669390400
transform 1 0 26768 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2166__A1
timestamp 1669390400
transform 1 0 33376 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2166__A2
timestamp 1669390400
transform 1 0 32032 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2167__I0
timestamp 1669390400
transform 1 0 34272 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2167__I1
timestamp 1669390400
transform 1 0 33824 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2167__S
timestamp 1669390400
transform -1 0 36848 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2169__A1
timestamp 1669390400
transform -1 0 25088 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2169__A2
timestamp 1669390400
transform 1 0 26432 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2169__B1
timestamp 1669390400
transform 1 0 29456 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2169__B2
timestamp 1669390400
transform 1 0 29792 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2169__C1
timestamp 1669390400
transform 1 0 25200 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2169__C2
timestamp 1669390400
transform 1 0 30800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2170__A1
timestamp 1669390400
transform 1 0 46144 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2170__A2
timestamp 1669390400
transform -1 0 44576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2171__A1
timestamp 1669390400
transform 1 0 45472 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2173__A1
timestamp 1669390400
transform -1 0 31136 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2173__A2
timestamp 1669390400
transform 1 0 32928 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2173__B
timestamp 1669390400
transform -1 0 30800 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2174__A1
timestamp 1669390400
transform -1 0 32704 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2175__A1
timestamp 1669390400
transform -1 0 40880 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2175__A2
timestamp 1669390400
transform 1 0 43008 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2176__A1
timestamp 1669390400
transform 1 0 31136 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2176__A2
timestamp 1669390400
transform -1 0 32592 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2177__A1
timestamp 1669390400
transform 1 0 30128 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2177__A2
timestamp 1669390400
transform 1 0 32816 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2177__B
timestamp 1669390400
transform 1 0 32592 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2178__A2
timestamp 1669390400
transform 1 0 43456 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2179__A2
timestamp 1669390400
transform 1 0 44912 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2181__A1
timestamp 1669390400
transform -1 0 54880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2181__A2
timestamp 1669390400
transform 1 0 54432 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2183__A1
timestamp 1669390400
transform -1 0 55328 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2183__A2
timestamp 1669390400
transform -1 0 54880 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2185__A1
timestamp 1669390400
transform 1 0 47040 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2187__A1
timestamp 1669390400
transform -1 0 45584 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2187__A2
timestamp 1669390400
transform -1 0 45024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2188__A2
timestamp 1669390400
transform -1 0 41328 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2189__A1
timestamp 1669390400
transform 1 0 35840 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2189__A2
timestamp 1669390400
transform 1 0 34720 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2190__A1
timestamp 1669390400
transform 1 0 36176 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2190__A2
timestamp 1669390400
transform 1 0 35728 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2191__A1
timestamp 1669390400
transform 1 0 36176 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2191__A2
timestamp 1669390400
transform 1 0 35728 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2192__A1
timestamp 1669390400
transform -1 0 42336 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2192__A2
timestamp 1669390400
transform -1 0 40544 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2193__A1
timestamp 1669390400
transform -1 0 25984 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2193__A2
timestamp 1669390400
transform 1 0 22624 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2194__A1
timestamp 1669390400
transform -1 0 30128 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2194__A2
timestamp 1669390400
transform -1 0 29680 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2194__B
timestamp 1669390400
transform 1 0 28560 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2195__A2
timestamp 1669390400
transform -1 0 39424 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2196__A1
timestamp 1669390400
transform -1 0 42224 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2198__A3
timestamp 1669390400
transform 1 0 32592 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2199__A2
timestamp 1669390400
transform -1 0 36400 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2200__I
timestamp 1669390400
transform 1 0 30800 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2201__A1
timestamp 1669390400
transform 1 0 37520 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2201__A2
timestamp 1669390400
transform 1 0 37072 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2201__B
timestamp 1669390400
transform 1 0 33488 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2205__A1
timestamp 1669390400
transform 1 0 31136 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2205__A2
timestamp 1669390400
transform 1 0 30688 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2206__A2
timestamp 1669390400
transform -1 0 33712 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2206__B1
timestamp 1669390400
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2206__B2
timestamp 1669390400
transform 1 0 31808 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2207__A1
timestamp 1669390400
transform 1 0 38752 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2207__A3
timestamp 1669390400
transform 1 0 37408 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2208__A3
timestamp 1669390400
transform -1 0 45808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2211__A1
timestamp 1669390400
transform 1 0 49840 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2212__A1
timestamp 1669390400
transform 1 0 44352 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2213__A1
timestamp 1669390400
transform -1 0 44128 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2215__A1
timestamp 1669390400
transform 1 0 53760 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2215__A2
timestamp 1669390400
transform 1 0 53536 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2216__A1
timestamp 1669390400
transform 1 0 47152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2216__A2
timestamp 1669390400
transform 1 0 46256 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2217__A1
timestamp 1669390400
transform -1 0 42672 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2217__A2
timestamp 1669390400
transform 1 0 42000 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2218__A1
timestamp 1669390400
transform 1 0 47600 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2218__A2
timestamp 1669390400
transform 1 0 47152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2219__A1
timestamp 1669390400
transform 1 0 48944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2219__A2
timestamp 1669390400
transform 1 0 47824 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2220__A1
timestamp 1669390400
transform 1 0 46928 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2220__A2
timestamp 1669390400
transform 1 0 46256 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2220__B
timestamp 1669390400
transform 1 0 48608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2221__A1
timestamp 1669390400
transform 1 0 48160 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2221__A3
timestamp 1669390400
transform 1 0 47712 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2222__A1
timestamp 1669390400
transform 1 0 51968 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2223__A1
timestamp 1669390400
transform -1 0 51296 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2229__A1
timestamp 1669390400
transform 1 0 52640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2233__A1
timestamp 1669390400
transform 1 0 49392 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2233__A2
timestamp 1669390400
transform 1 0 48944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2235__A1
timestamp 1669390400
transform 1 0 51184 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2237__A1
timestamp 1669390400
transform 1 0 44352 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2239__A1
timestamp 1669390400
transform 1 0 50736 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2239__A2
timestamp 1669390400
transform 1 0 49504 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2240__A1
timestamp 1669390400
transform 1 0 18592 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2241__I
timestamp 1669390400
transform -1 0 40096 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2242__A1
timestamp 1669390400
transform -1 0 39760 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2242__A2
timestamp 1669390400
transform -1 0 41664 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2243__A1
timestamp 1669390400
transform 1 0 46032 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2243__A2
timestamp 1669390400
transform 1 0 46480 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2243__A3
timestamp 1669390400
transform 1 0 47376 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2244__A1
timestamp 1669390400
transform 1 0 49952 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2244__A2
timestamp 1669390400
transform 1 0 51184 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2245__A2
timestamp 1669390400
transform 1 0 49728 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2248__A2
timestamp 1669390400
transform -1 0 46816 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2249__A2
timestamp 1669390400
transform 1 0 47824 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2251__A2
timestamp 1669390400
transform 1 0 41440 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2253__A2
timestamp 1669390400
transform 1 0 35280 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2253__B
timestamp 1669390400
transform 1 0 36400 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2254__A1
timestamp 1669390400
transform 1 0 36624 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2256__I
timestamp 1669390400
transform -1 0 26432 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2257__I
timestamp 1669390400
transform -1 0 44128 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2258__A1
timestamp 1669390400
transform 1 0 36624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2258__A2
timestamp 1669390400
transform 1 0 38080 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2258__B1
timestamp 1669390400
transform 1 0 39872 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2258__B2
timestamp 1669390400
transform 1 0 38528 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2259__A1
timestamp 1669390400
transform -1 0 39200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2259__A2
timestamp 1669390400
transform 1 0 37520 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2262__A1
timestamp 1669390400
transform 1 0 32144 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2262__A2
timestamp 1669390400
transform -1 0 33040 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2265__A3
timestamp 1669390400
transform -1 0 35728 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2266__A1
timestamp 1669390400
transform 1 0 35952 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2266__A2
timestamp 1669390400
transform -1 0 33712 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2267__I0
timestamp 1669390400
transform 1 0 35952 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2267__S
timestamp 1669390400
transform -1 0 35280 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2271__A1
timestamp 1669390400
transform 1 0 26096 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2271__A2
timestamp 1669390400
transform 1 0 25536 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2271__B1
timestamp 1669390400
transform 1 0 27888 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2271__B2
timestamp 1669390400
transform -1 0 26208 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2271__C1
timestamp 1669390400
transform 1 0 36400 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2271__C2
timestamp 1669390400
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2273__A1
timestamp 1669390400
transform -1 0 43232 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2284__A1
timestamp 1669390400
transform 1 0 47824 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2285__A1
timestamp 1669390400
transform -1 0 48944 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2285__A2
timestamp 1669390400
transform -1 0 48496 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2289__A1
timestamp 1669390400
transform 1 0 46928 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2290__A1
timestamp 1669390400
transform 1 0 25648 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2290__A2
timestamp 1669390400
transform -1 0 28112 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2291__A1
timestamp 1669390400
transform -1 0 46704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2291__A2
timestamp 1669390400
transform 1 0 44688 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2292__A1
timestamp 1669390400
transform 1 0 44464 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2292__A2
timestamp 1669390400
transform 1 0 44912 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2293__A1
timestamp 1669390400
transform -1 0 45584 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2295__A1
timestamp 1669390400
transform 1 0 47040 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2297__A1
timestamp 1669390400
transform -1 0 42784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2300__A1
timestamp 1669390400
transform -1 0 37968 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2301__A1
timestamp 1669390400
transform 1 0 40768 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2301__A2
timestamp 1669390400
transform 1 0 42000 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2302__A1
timestamp 1669390400
transform -1 0 40544 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2302__A2
timestamp 1669390400
transform 1 0 40768 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2302__B1
timestamp 1669390400
transform 1 0 41440 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2302__B2
timestamp 1669390400
transform 1 0 41552 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2303__A2
timestamp 1669390400
transform -1 0 42112 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2305__A1
timestamp 1669390400
transform 1 0 29008 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2305__A2
timestamp 1669390400
transform -1 0 32928 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2306__I1
timestamp 1669390400
transform 1 0 37296 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2306__S
timestamp 1669390400
transform 1 0 36848 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2307__A1
timestamp 1669390400
transform 1 0 40320 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2308__A1
timestamp 1669390400
transform 1 0 29456 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2308__A2
timestamp 1669390400
transform 1 0 27216 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2308__B1
timestamp 1669390400
transform 1 0 26768 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2308__B2
timestamp 1669390400
transform 1 0 27440 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2308__C1
timestamp 1669390400
transform 1 0 30800 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2308__C2
timestamp 1669390400
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2321__A2
timestamp 1669390400
transform 1 0 54880 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2322__A1
timestamp 1669390400
transform 1 0 56672 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2324__A1
timestamp 1669390400
transform 1 0 45360 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2324__A2
timestamp 1669390400
transform 1 0 48608 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2325__A1
timestamp 1669390400
transform 1 0 41776 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2325__A2
timestamp 1669390400
transform 1 0 41328 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2325__A3
timestamp 1669390400
transform 1 0 43568 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2326__A1
timestamp 1669390400
transform 1 0 46032 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2326__A2
timestamp 1669390400
transform 1 0 44688 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2326__B
timestamp 1669390400
transform 1 0 44240 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2328__A1
timestamp 1669390400
transform 1 0 49840 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2329__A1
timestamp 1669390400
transform 1 0 49392 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2330__B2
timestamp 1669390400
transform -1 0 50512 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2331__B
timestamp 1669390400
transform 1 0 32480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2332__I0
timestamp 1669390400
transform 1 0 37856 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2332__I1
timestamp 1669390400
transform 1 0 33936 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2332__S
timestamp 1669390400
transform 1 0 31584 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2333__A1
timestamp 1669390400
transform -1 0 33040 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2333__A2
timestamp 1669390400
transform 1 0 37408 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2334__A1
timestamp 1669390400
transform -1 0 33712 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2334__A2
timestamp 1669390400
transform 1 0 33824 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2335__A1
timestamp 1669390400
transform 1 0 43008 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2335__A2
timestamp 1669390400
transform 1 0 40432 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2336__A1
timestamp 1669390400
transform 1 0 44016 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2338__A3
timestamp 1669390400
transform 1 0 43456 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2339__A1
timestamp 1669390400
transform 1 0 38528 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2339__A2
timestamp 1669390400
transform 1 0 37408 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2339__B
timestamp 1669390400
transform 1 0 36624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2340__A1
timestamp 1669390400
transform -1 0 44688 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2340__A2
timestamp 1669390400
transform 1 0 42224 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2341__A2
timestamp 1669390400
transform 1 0 41888 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2342__A1
timestamp 1669390400
transform 1 0 53312 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2343__A1
timestamp 1669390400
transform 1 0 56112 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2344__A1
timestamp 1669390400
transform 1 0 54880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2346__A1
timestamp 1669390400
transform 1 0 32256 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2346__A2
timestamp 1669390400
transform 1 0 31808 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2347__A1
timestamp 1669390400
transform -1 0 24192 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2347__A2
timestamp 1669390400
transform -1 0 18144 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2348__A1
timestamp 1669390400
transform 1 0 32592 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2348__A2
timestamp 1669390400
transform -1 0 34944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2348__B1
timestamp 1669390400
transform -1 0 32368 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2348__B2
timestamp 1669390400
transform 1 0 34832 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2349__A2
timestamp 1669390400
transform 1 0 31248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2349__B1
timestamp 1669390400
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2349__B2
timestamp 1669390400
transform -1 0 24640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2349__C1
timestamp 1669390400
transform -1 0 29792 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2349__C2
timestamp 1669390400
transform 1 0 30800 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2350__A1
timestamp 1669390400
transform 1 0 39200 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2352__A1
timestamp 1669390400
transform 1 0 37856 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2355__A1
timestamp 1669390400
transform 1 0 42672 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2357__A1
timestamp 1669390400
transform 1 0 44352 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2360__A1
timestamp 1669390400
transform 1 0 56672 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2360__A2
timestamp 1669390400
transform -1 0 56672 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2361__A2
timestamp 1669390400
transform -1 0 54432 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2362__A1
timestamp 1669390400
transform -1 0 56448 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2362__A2
timestamp 1669390400
transform -1 0 56896 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2371__A1
timestamp 1669390400
transform 1 0 58464 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2374__A1
timestamp 1669390400
transform 1 0 41328 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2374__A2
timestamp 1669390400
transform 1 0 44464 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2375__A1
timestamp 1669390400
transform 1 0 22512 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2375__A2
timestamp 1669390400
transform -1 0 25088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2376__A1
timestamp 1669390400
transform -1 0 15904 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2376__A2
timestamp 1669390400
transform -1 0 13776 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2377__A1
timestamp 1669390400
transform 1 0 39984 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2377__A2
timestamp 1669390400
transform -1 0 39648 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2377__B1
timestamp 1669390400
transform 1 0 40432 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2377__B2
timestamp 1669390400
transform 1 0 38976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2378__I0
timestamp 1669390400
transform 1 0 38752 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2378__I1
timestamp 1669390400
transform 1 0 38304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2378__S
timestamp 1669390400
transform -1 0 37856 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2379__A1
timestamp 1669390400
transform 1 0 37856 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2379__A2
timestamp 1669390400
transform 1 0 38864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2379__B2
timestamp 1669390400
transform -1 0 36512 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2380__A1
timestamp 1669390400
transform 1 0 44016 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2380__A2
timestamp 1669390400
transform 1 0 43120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2382__A1
timestamp 1669390400
transform -1 0 40544 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2383__A1
timestamp 1669390400
transform 1 0 44576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2383__B2
timestamp 1669390400
transform 1 0 41440 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2384__A1
timestamp 1669390400
transform 1 0 51968 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2385__A1
timestamp 1669390400
transform -1 0 45136 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2385__A2
timestamp 1669390400
transform 1 0 48272 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2386__I0
timestamp 1669390400
transform 1 0 47712 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2386__S
timestamp 1669390400
transform 1 0 47488 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2387__A1
timestamp 1669390400
transform 1 0 45360 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2387__B2
timestamp 1669390400
transform 1 0 46928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2388__A1
timestamp 1669390400
transform 1 0 48720 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2391__A1
timestamp 1669390400
transform 1 0 51296 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2392__A1
timestamp 1669390400
transform 1 0 52080 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2394__A1
timestamp 1669390400
transform -1 0 52864 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2395__A1
timestamp 1669390400
transform 1 0 37744 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2396__A1
timestamp 1669390400
transform -1 0 27664 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2396__A2
timestamp 1669390400
transform -1 0 19264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2397__A1
timestamp 1669390400
transform 1 0 29456 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2397__B
timestamp 1669390400
transform 1 0 28784 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2397__C
timestamp 1669390400
transform 1 0 28336 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2398__A1
timestamp 1669390400
transform 1 0 38304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2399__A1
timestamp 1669390400
transform 1 0 35280 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2399__A3
timestamp 1669390400
transform 1 0 36064 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2401__A2
timestamp 1669390400
transform 1 0 39872 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2404__A1
timestamp 1669390400
transform 1 0 44352 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2408__A1
timestamp 1669390400
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2418__A1
timestamp 1669390400
transform 1 0 56560 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2419__A1
timestamp 1669390400
transform 1 0 58240 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2420__A1
timestamp 1669390400
transform 1 0 56560 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2421__A1
timestamp 1669390400
transform 1 0 57680 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2423__A1
timestamp 1669390400
transform 1 0 57568 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2424__A1
timestamp 1669390400
transform 1 0 41888 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2424__A2
timestamp 1669390400
transform 1 0 42336 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2424__A3
timestamp 1669390400
transform 1 0 42784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2425__A1
timestamp 1669390400
transform 1 0 41440 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2425__A2
timestamp 1669390400
transform 1 0 40320 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2426__A1
timestamp 1669390400
transform 1 0 43232 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2426__A2
timestamp 1669390400
transform 1 0 42560 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2428__A1
timestamp 1669390400
transform 1 0 38080 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2428__A2
timestamp 1669390400
transform 1 0 40768 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2429__A1
timestamp 1669390400
transform 1 0 42336 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2430__A1
timestamp 1669390400
transform 1 0 44352 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2432__A1
timestamp 1669390400
transform 1 0 43904 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2434__A1
timestamp 1669390400
transform 1 0 48272 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2437__A1
timestamp 1669390400
transform 1 0 40320 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2437__A2
timestamp 1669390400
transform 1 0 41664 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2438__A1
timestamp 1669390400
transform -1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2438__A2
timestamp 1669390400
transform -1 0 37408 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2439__A1
timestamp 1669390400
transform 1 0 39648 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2439__A2
timestamp 1669390400
transform 1 0 38752 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2440__A1
timestamp 1669390400
transform 1 0 36512 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2440__A2
timestamp 1669390400
transform 1 0 36064 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2440__B1
timestamp 1669390400
transform -1 0 35840 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2440__B2
timestamp 1669390400
transform 1 0 37408 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2441__A3
timestamp 1669390400
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2442__A1
timestamp 1669390400
transform 1 0 34272 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2442__A2
timestamp 1669390400
transform 1 0 38976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2442__B1
timestamp 1669390400
transform 1 0 32928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2442__B2
timestamp 1669390400
transform 1 0 33824 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2442__C
timestamp 1669390400
transform 1 0 31472 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2443__A1
timestamp 1669390400
transform 1 0 39424 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2443__B2
timestamp 1669390400
transform -1 0 37184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2444__A1
timestamp 1669390400
transform 1 0 38528 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2444__A2
timestamp 1669390400
transform 1 0 38192 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2445__A1
timestamp 1669390400
transform 1 0 39872 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2447__A1
timestamp 1669390400
transform 1 0 48608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2447__A2
timestamp 1669390400
transform 1 0 48160 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2449__A1
timestamp 1669390400
transform -1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2449__A2
timestamp 1669390400
transform -1 0 47936 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2452__A2
timestamp 1669390400
transform -1 0 49392 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2453__A2
timestamp 1669390400
transform 1 0 52080 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2462__A1
timestamp 1669390400
transform -1 0 54992 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2462__A2
timestamp 1669390400
transform 1 0 54320 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2462__A3
timestamp 1669390400
transform 1 0 56672 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2462__B
timestamp 1669390400
transform -1 0 56448 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2466__A1
timestamp 1669390400
transform 1 0 42112 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2466__A2
timestamp 1669390400
transform -1 0 44464 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2467__I
timestamp 1669390400
transform 1 0 43904 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2468__A1
timestamp 1669390400
transform 1 0 40880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2468__A2
timestamp 1669390400
transform 1 0 41888 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2469__A1
timestamp 1669390400
transform -1 0 44688 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2470__A1
timestamp 1669390400
transform 1 0 44688 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2470__A2
timestamp 1669390400
transform 1 0 45136 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2470__B1
timestamp 1669390400
transform 1 0 43792 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2471__A1
timestamp 1669390400
transform 1 0 31360 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2471__A2
timestamp 1669390400
transform 1 0 31808 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2472__A1
timestamp 1669390400
transform -1 0 35392 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2473__A1
timestamp 1669390400
transform -1 0 40992 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2473__A2
timestamp 1669390400
transform 1 0 40880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2474__A1
timestamp 1669390400
transform 1 0 43008 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2474__A2
timestamp 1669390400
transform 1 0 41888 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2476__A1
timestamp 1669390400
transform -1 0 43008 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2477__A1
timestamp 1669390400
transform 1 0 44688 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2479__A1
timestamp 1669390400
transform -1 0 46480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2483__A1
timestamp 1669390400
transform 1 0 33376 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2483__A2
timestamp 1669390400
transform 1 0 33488 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2484__A2
timestamp 1669390400
transform -1 0 32704 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2485__A1
timestamp 1669390400
transform 1 0 37408 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2485__A2
timestamp 1669390400
transform -1 0 36848 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2485__B1
timestamp 1669390400
transform 1 0 36512 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2486__A1
timestamp 1669390400
transform 1 0 36736 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2486__A2
timestamp 1669390400
transform -1 0 35056 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2487__A1
timestamp 1669390400
transform 1 0 37408 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2487__A2
timestamp 1669390400
transform 1 0 34720 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2487__B
timestamp 1669390400
transform 1 0 34720 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2488__A1
timestamp 1669390400
transform -1 0 35280 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2488__B2
timestamp 1669390400
transform 1 0 37856 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2489__A1
timestamp 1669390400
transform 1 0 37856 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2492__A1
timestamp 1669390400
transform 1 0 38752 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2493__A1
timestamp 1669390400
transform 1 0 36736 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2494__A1
timestamp 1669390400
transform 1 0 38752 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2495__A3
timestamp 1669390400
transform -1 0 38528 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2500__A1
timestamp 1669390400
transform -1 0 46144 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2500__A2
timestamp 1669390400
transform 1 0 45696 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2511__A1
timestamp 1669390400
transform 1 0 55664 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2512__A1
timestamp 1669390400
transform 1 0 55440 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2515__A1
timestamp 1669390400
transform 1 0 58464 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2516__A1
timestamp 1669390400
transform 1 0 39536 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2516__A2
timestamp 1669390400
transform 1 0 41440 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2516__A3
timestamp 1669390400
transform 1 0 41664 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2517__A1
timestamp 1669390400
transform 1 0 38416 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2517__A2
timestamp 1669390400
transform 1 0 41216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2518__A1
timestamp 1669390400
transform -1 0 38976 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2519__A1
timestamp 1669390400
transform 1 0 41776 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2520__I1
timestamp 1669390400
transform 1 0 42000 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2520__S
timestamp 1669390400
transform 1 0 44128 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2521__A1
timestamp 1669390400
transform 1 0 43008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2523__A1
timestamp 1669390400
transform 1 0 45584 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2525__A1
timestamp 1669390400
transform 1 0 43120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2528__B
timestamp 1669390400
transform 1 0 49168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2530__A1
timestamp 1669390400
transform -1 0 48944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2531__A1
timestamp 1669390400
transform -1 0 33712 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2531__A2
timestamp 1669390400
transform 1 0 33936 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2532__A1
timestamp 1669390400
transform 1 0 37408 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2533__B
timestamp 1669390400
transform 1 0 37856 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2534__A2
timestamp 1669390400
transform -1 0 29008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2534__B
timestamp 1669390400
transform -1 0 31136 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2535__I0
timestamp 1669390400
transform 1 0 31360 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2535__I1
timestamp 1669390400
transform -1 0 32368 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2535__S
timestamp 1669390400
transform 1 0 32592 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2536__A1
timestamp 1669390400
transform -1 0 34608 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2536__A2
timestamp 1669390400
transform 1 0 36512 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2538__A1
timestamp 1669390400
transform 1 0 39200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2541__A1
timestamp 1669390400
transform -1 0 38976 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2542__A1
timestamp 1669390400
transform 1 0 47824 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2542__A2
timestamp 1669390400
transform 1 0 48160 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2544__A1
timestamp 1669390400
transform 1 0 45584 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2544__A2
timestamp 1669390400
transform 1 0 46032 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2557__A1
timestamp 1669390400
transform 1 0 53760 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2558__A1
timestamp 1669390400
transform 1 0 52192 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2561__A1
timestamp 1669390400
transform -1 0 57344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2562__A1
timestamp 1669390400
transform 1 0 42672 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2562__A2
timestamp 1669390400
transform -1 0 42448 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2563__A1
timestamp 1669390400
transform 1 0 43904 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2563__A2
timestamp 1669390400
transform 1 0 44688 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2564__A1
timestamp 1669390400
transform 1 0 45136 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2565__A1
timestamp 1669390400
transform 1 0 45024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2567__A1
timestamp 1669390400
transform 1 0 48720 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2568__A1
timestamp 1669390400
transform 1 0 48272 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2571__I1
timestamp 1669390400
transform 1 0 33152 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2571__S
timestamp 1669390400
transform 1 0 29568 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2572__A1
timestamp 1669390400
transform 1 0 31696 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2572__A2
timestamp 1669390400
transform -1 0 32816 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2572__B1
timestamp 1669390400
transform 1 0 32144 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2572__B2
timestamp 1669390400
transform 1 0 31472 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2574__A1
timestamp 1669390400
transform 1 0 45136 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2574__A2
timestamp 1669390400
transform 1 0 43120 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2575__A1
timestamp 1669390400
transform 1 0 43456 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2576__A1
timestamp 1669390400
transform 1 0 47040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2576__A2
timestamp 1669390400
transform 1 0 45584 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2580__A2
timestamp 1669390400
transform 1 0 45360 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2581__A2
timestamp 1669390400
transform 1 0 45920 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2583__A1
timestamp 1669390400
transform -1 0 46032 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2583__A2
timestamp 1669390400
transform -1 0 45808 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2593__A1
timestamp 1669390400
transform -1 0 33712 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2593__A2
timestamp 1669390400
transform 1 0 33712 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2594__A1
timestamp 1669390400
transform 1 0 35392 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2594__A2
timestamp 1669390400
transform 1 0 36288 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2595__I0
timestamp 1669390400
transform 1 0 33936 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2595__S
timestamp 1669390400
transform 1 0 33488 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2596__A1
timestamp 1669390400
transform -1 0 32480 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2596__B2
timestamp 1669390400
transform -1 0 32032 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2597__A1
timestamp 1669390400
transform 1 0 34944 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2597__A2
timestamp 1669390400
transform 1 0 35952 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2598__A1
timestamp 1669390400
transform -1 0 40768 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2598__A2
timestamp 1669390400
transform -1 0 41664 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2599__A1
timestamp 1669390400
transform 1 0 45472 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2600__A1
timestamp 1669390400
transform -1 0 42112 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2601__A1
timestamp 1669390400
transform -1 0 43904 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2603__A1
timestamp 1669390400
transform 1 0 35952 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2604__A2
timestamp 1669390400
transform -1 0 34272 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2606__A1
timestamp 1669390400
transform 1 0 45360 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2607__A1
timestamp 1669390400
transform -1 0 41664 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2607__B2
timestamp 1669390400
transform -1 0 44576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2608__A1
timestamp 1669390400
transform 1 0 43232 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2616__A2
timestamp 1669390400
transform 1 0 53760 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2623__A1
timestamp 1669390400
transform 1 0 36400 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2623__A2
timestamp 1669390400
transform -1 0 36064 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2625__A1
timestamp 1669390400
transform -1 0 33712 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2625__B2
timestamp 1669390400
transform 1 0 32928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2626__I
timestamp 1669390400
transform 1 0 36176 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2627__A1
timestamp 1669390400
transform -1 0 33040 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2628__A2
timestamp 1669390400
transform 1 0 35728 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2629__A1
timestamp 1669390400
transform 1 0 41888 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2629__A2
timestamp 1669390400
transform 1 0 39760 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2629__B
timestamp 1669390400
transform 1 0 41440 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2630__A1
timestamp 1669390400
transform 1 0 38304 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2630__A2
timestamp 1669390400
transform -1 0 40320 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2631__A1
timestamp 1669390400
transform -1 0 39424 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2632__A1
timestamp 1669390400
transform -1 0 35504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2632__A2
timestamp 1669390400
transform -1 0 34608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2636__A1
timestamp 1669390400
transform -1 0 41888 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2636__B2
timestamp 1669390400
transform -1 0 39872 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2639__A1
timestamp 1669390400
transform -1 0 40432 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2642__A1
timestamp 1669390400
transform 1 0 43120 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2644__A1
timestamp 1669390400
transform -1 0 34160 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2644__A2
timestamp 1669390400
transform 1 0 33488 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2645__A1
timestamp 1669390400
transform -1 0 34720 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2647__I1
timestamp 1669390400
transform 1 0 35392 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2648__A1
timestamp 1669390400
transform -1 0 36624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2651__A1
timestamp 1669390400
transform 1 0 42560 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2652__A1
timestamp 1669390400
transform -1 0 41664 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2659__A1
timestamp 1669390400
transform 1 0 45360 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2660__A1
timestamp 1669390400
transform 1 0 39984 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2661__A1
timestamp 1669390400
transform 1 0 37856 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2662__A1
timestamp 1669390400
transform 1 0 38416 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2662__A2
timestamp 1669390400
transform 1 0 38864 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2681__B
timestamp 1669390400
transform 1 0 57680 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2682__A1
timestamp 1669390400
transform 1 0 56112 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2683__A1
timestamp 1669390400
transform 1 0 53760 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2688__A3
timestamp 1669390400
transform -1 0 56336 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2689__A1
timestamp 1669390400
transform -1 0 58128 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2693__A1
timestamp 1669390400
transform 1 0 58352 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2694__A2
timestamp 1669390400
transform 1 0 43344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2695__A1
timestamp 1669390400
transform 1 0 43568 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2695__A2
timestamp 1669390400
transform -1 0 44800 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2696__A1
timestamp 1669390400
transform 1 0 45696 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2697__A1
timestamp 1669390400
transform 1 0 44128 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2704__A1
timestamp 1669390400
transform 1 0 38752 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2704__B1
timestamp 1669390400
transform 1 0 37520 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2705__A1
timestamp 1669390400
transform -1 0 38528 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2705__A2
timestamp 1669390400
transform 1 0 41216 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2705__B1
timestamp 1669390400
transform 1 0 42112 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2705__B2
timestamp 1669390400
transform 1 0 38528 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2706__A1
timestamp 1669390400
transform 1 0 42896 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2707__A1
timestamp 1669390400
transform 1 0 41440 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2709__A1
timestamp 1669390400
transform -1 0 25088 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2709__A2
timestamp 1669390400
transform -1 0 24640 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2710__A1
timestamp 1669390400
transform -1 0 36624 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2710__A2
timestamp 1669390400
transform 1 0 37296 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2710__B1
timestamp 1669390400
transform 1 0 36848 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2710__B2
timestamp 1669390400
transform 1 0 37744 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2711__A1
timestamp 1669390400
transform 1 0 39088 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2711__A2
timestamp 1669390400
transform 1 0 29680 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2711__B1
timestamp 1669390400
transform 1 0 28784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2711__B2
timestamp 1669390400
transform -1 0 29008 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2711__C1
timestamp 1669390400
transform 1 0 28336 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2711__C2
timestamp 1669390400
transform 1 0 31584 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2720__A1
timestamp 1669390400
transform -1 0 42672 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2724__A1
timestamp 1669390400
transform 1 0 41440 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2725__A1
timestamp 1669390400
transform 1 0 41776 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2725__A2
timestamp 1669390400
transform 1 0 42672 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2726__A1
timestamp 1669390400
transform 1 0 43792 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2727__A1
timestamp 1669390400
transform 1 0 38640 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2727__A2
timestamp 1669390400
transform 1 0 38192 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2731__A1
timestamp 1669390400
transform -1 0 40320 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2731__A2
timestamp 1669390400
transform 1 0 36512 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2732__A1
timestamp 1669390400
transform 1 0 38304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2732__A2
timestamp 1669390400
transform 1 0 37408 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2732__B
timestamp 1669390400
transform 1 0 37856 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2733__A2
timestamp 1669390400
transform -1 0 37632 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2734__A1
timestamp 1669390400
transform 1 0 27888 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2734__A2
timestamp 1669390400
transform 1 0 36400 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2734__B1
timestamp 1669390400
transform 1 0 29792 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2734__B2
timestamp 1669390400
transform -1 0 29680 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2734__C1
timestamp 1669390400
transform 1 0 36736 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2734__C2
timestamp 1669390400
transform 1 0 38080 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2735__A2
timestamp 1669390400
transform -1 0 37184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2741__A1
timestamp 1669390400
transform 1 0 48832 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2759__A1
timestamp 1669390400
transform -1 0 41440 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2763__A2
timestamp 1669390400
transform 1 0 39424 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2764__A1
timestamp 1669390400
transform 1 0 39872 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2764__A2
timestamp 1669390400
transform 1 0 40992 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2765__A1
timestamp 1669390400
transform 1 0 40320 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2767__A2
timestamp 1669390400
transform 1 0 37856 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2768__A1
timestamp 1669390400
transform -1 0 32256 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2768__A2
timestamp 1669390400
transform 1 0 35168 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2769__A1
timestamp 1669390400
transform 1 0 37072 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2769__A2
timestamp 1669390400
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2769__B
timestamp 1669390400
transform -1 0 37072 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2771__A1
timestamp 1669390400
transform -1 0 37632 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2771__A2
timestamp 1669390400
transform 1 0 26544 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2771__B1
timestamp 1669390400
transform 1 0 25648 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2771__B2
timestamp 1669390400
transform -1 0 27664 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2771__C1
timestamp 1669390400
transform 1 0 28336 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2771__C2
timestamp 1669390400
transform 1 0 28784 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2776__A1
timestamp 1669390400
transform 1 0 41104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2785__A1
timestamp 1669390400
transform 1 0 38416 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2785__A2
timestamp 1669390400
transform 1 0 40544 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2785__B
timestamp 1669390400
transform -1 0 38080 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2787__A1
timestamp 1669390400
transform 1 0 29008 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2787__A2
timestamp 1669390400
transform 1 0 28672 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2788__A1
timestamp 1669390400
transform -1 0 29008 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2788__A2
timestamp 1669390400
transform 1 0 25648 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2788__B
timestamp 1669390400
transform -1 0 31248 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2790__A1
timestamp 1669390400
transform 1 0 26096 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2790__A2
timestamp 1669390400
transform 1 0 27888 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2790__B1
timestamp 1669390400
transform 1 0 28336 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2790__B2
timestamp 1669390400
transform 1 0 38304 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2790__C1
timestamp 1669390400
transform 1 0 28784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2790__C2
timestamp 1669390400
transform -1 0 28560 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2796__A1
timestamp 1669390400
transform 1 0 40320 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2805__A2
timestamp 1669390400
transform -1 0 54096 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2815__A1
timestamp 1669390400
transform 1 0 53088 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2815__A2
timestamp 1669390400
transform 1 0 52864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2829__A1
timestamp 1669390400
transform 1 0 26096 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2829__A2
timestamp 1669390400
transform 1 0 26208 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2829__B
timestamp 1669390400
transform -1 0 26880 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2832__A1
timestamp 1669390400
transform -1 0 32144 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2832__A2
timestamp 1669390400
transform 1 0 22624 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2832__B1
timestamp 1669390400
transform 1 0 26320 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2832__B2
timestamp 1669390400
transform 1 0 34272 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2832__C1
timestamp 1669390400
transform 1 0 34720 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2832__C2
timestamp 1669390400
transform 1 0 25760 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2833__A1
timestamp 1669390400
transform 1 0 27440 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2833__A2
timestamp 1669390400
transform 1 0 27888 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2834__A1
timestamp 1669390400
transform 1 0 24416 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2834__A2
timestamp 1669390400
transform 1 0 27888 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2834__B
timestamp 1669390400
transform -1 0 26096 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2853__A1
timestamp 1669390400
transform -1 0 20272 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2853__A2
timestamp 1669390400
transform -1 0 20608 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2854__A1
timestamp 1669390400
transform 1 0 28448 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2854__A2
timestamp 1669390400
transform -1 0 19824 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2854__B1
timestamp 1669390400
transform -1 0 20720 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2854__B2
timestamp 1669390400
transform -1 0 18816 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2856__A1
timestamp 1669390400
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2856__A2
timestamp 1669390400
transform 1 0 22960 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2856__B1
timestamp 1669390400
transform 1 0 23296 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2856__B2
timestamp 1669390400
transform -1 0 32592 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2856__C1
timestamp 1669390400
transform 1 0 33824 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2856__C2
timestamp 1669390400
transform 1 0 37408 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2857__A2
timestamp 1669390400
transform -1 0 21504 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2860__A2
timestamp 1669390400
transform -1 0 21952 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2868__A1
timestamp 1669390400
transform 1 0 36960 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2869__A1
timestamp 1669390400
transform -1 0 35616 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2872__A1
timestamp 1669390400
transform 1 0 45920 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2875__A2
timestamp 1669390400
transform 1 0 36960 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2881__A1
timestamp 1669390400
transform -1 0 7840 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2881__A2
timestamp 1669390400
transform -1 0 2800 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2882__A1
timestamp 1669390400
transform -1 0 8176 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2882__A2
timestamp 1669390400
transform -1 0 8624 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2883__A1
timestamp 1669390400
transform -1 0 22064 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2883__A2
timestamp 1669390400
transform -1 0 25088 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2883__B1
timestamp 1669390400
transform -1 0 25424 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2883__B2
timestamp 1669390400
transform -1 0 21616 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2884__A2
timestamp 1669390400
transform -1 0 7280 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2886__I
timestamp 1669390400
transform 1 0 26992 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2888__A2
timestamp 1669390400
transform 1 0 27776 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2893__A1
timestamp 1669390400
transform 1 0 31248 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2893__A2
timestamp 1669390400
transform -1 0 29456 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2896__A1
timestamp 1669390400
transform 1 0 30128 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2896__A2
timestamp 1669390400
transform -1 0 30800 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2899__A1
timestamp 1669390400
transform -1 0 35728 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2900__I
timestamp 1669390400
transform 1 0 54432 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2901__A1
timestamp 1669390400
transform 1 0 52640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2903__A1
timestamp 1669390400
transform -1 0 55440 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2904__A1
timestamp 1669390400
transform -1 0 53536 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2906__A1
timestamp 1669390400
transform -1 0 55888 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2912__A1
timestamp 1669390400
transform 1 0 55440 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2912__B
timestamp 1669390400
transform 1 0 54992 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2913__B2
timestamp 1669390400
transform 1 0 58464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2915__A3
timestamp 1669390400
transform 1 0 56672 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2916__A1
timestamp 1669390400
transform 1 0 58240 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2918__A2
timestamp 1669390400
transform 1 0 55216 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2920__A1
timestamp 1669390400
transform -1 0 43008 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2923__A1
timestamp 1669390400
transform -1 0 45024 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2925__B
timestamp 1669390400
transform 1 0 41216 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2926__A1
timestamp 1669390400
transform 1 0 35056 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2926__B1
timestamp 1669390400
transform 1 0 35504 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2928__A1
timestamp 1669390400
transform 1 0 45472 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2930__A1
timestamp 1669390400
transform 1 0 37408 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2930__B2
timestamp 1669390400
transform 1 0 37632 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2931__I
timestamp 1669390400
transform 1 0 28560 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2932__A2
timestamp 1669390400
transform 1 0 54432 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2936__A1
timestamp 1669390400
transform 1 0 53984 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2936__A2
timestamp 1669390400
transform 1 0 53536 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2939__A1
timestamp 1669390400
transform 1 0 47712 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2939__A2
timestamp 1669390400
transform -1 0 49168 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2939__B2
timestamp 1669390400
transform 1 0 48384 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2940__A2
timestamp 1669390400
transform 1 0 56560 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2940__A3
timestamp 1669390400
transform 1 0 56448 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2943__A1
timestamp 1669390400
transform 1 0 54432 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2943__A2
timestamp 1669390400
transform -1 0 54208 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2944__A1
timestamp 1669390400
transform 1 0 55776 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2944__A2
timestamp 1669390400
transform 1 0 55328 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2945__A1
timestamp 1669390400
transform 1 0 52640 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2945__A2
timestamp 1669390400
transform 1 0 53536 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2947__A1
timestamp 1669390400
transform 1 0 57120 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2947__A2
timestamp 1669390400
transform 1 0 56672 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2949__A1
timestamp 1669390400
transform -1 0 52304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2949__B
timestamp 1669390400
transform 1 0 51856 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2952__A1
timestamp 1669390400
transform -1 0 50288 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2953__A1
timestamp 1669390400
transform 1 0 51072 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2954__A1
timestamp 1669390400
transform 1 0 53088 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2956__A1
timestamp 1669390400
transform 1 0 50848 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2956__B2
timestamp 1669390400
transform -1 0 51520 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2957__A1
timestamp 1669390400
transform 1 0 54096 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2958__A1
timestamp 1669390400
transform 1 0 51072 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2958__A2
timestamp 1669390400
transform 1 0 53088 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2964__A1
timestamp 1669390400
transform 1 0 47264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2965__A2
timestamp 1669390400
transform -1 0 48384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2965__B2
timestamp 1669390400
transform 1 0 46480 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2966__I
timestamp 1669390400
transform 1 0 35616 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2967__A1
timestamp 1669390400
transform 1 0 45024 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2971__B
timestamp 1669390400
transform 1 0 42560 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2972__A1
timestamp 1669390400
transform 1 0 40992 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2973__A1
timestamp 1669390400
transform -1 0 43456 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2973__B2
timestamp 1669390400
transform 1 0 42784 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2978__A1
timestamp 1669390400
transform 1 0 6720 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2978__A2
timestamp 1669390400
transform 1 0 8064 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2979__A2
timestamp 1669390400
transform -1 0 5152 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2980__A1
timestamp 1669390400
transform -1 0 2128 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2980__A2
timestamp 1669390400
transform 1 0 8960 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2981__A1
timestamp 1669390400
transform -1 0 24976 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2981__A2
timestamp 1669390400
transform -1 0 22176 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2981__B1
timestamp 1669390400
transform -1 0 20608 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2981__B2
timestamp 1669390400
transform 1 0 20832 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2982__A2
timestamp 1669390400
transform -1 0 9072 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2996__A1
timestamp 1669390400
transform -1 0 34832 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2997__B
timestamp 1669390400
transform 1 0 32592 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2998__A1
timestamp 1669390400
transform 1 0 32144 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2999__B1
timestamp 1669390400
transform 1 0 40320 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3003__A2
timestamp 1669390400
transform -1 0 33264 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3004__A1
timestamp 1669390400
transform 1 0 45360 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3004__C
timestamp 1669390400
transform 1 0 41440 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3005__A2
timestamp 1669390400
transform -1 0 5936 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3006__A1
timestamp 1669390400
transform -1 0 6048 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3006__A2
timestamp 1669390400
transform 1 0 6272 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3007__A2
timestamp 1669390400
transform 1 0 10080 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3008__A1
timestamp 1669390400
transform 1 0 22624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3008__A2
timestamp 1669390400
transform -1 0 22400 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3009__A1
timestamp 1669390400
transform 1 0 28224 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3009__A2
timestamp 1669390400
transform 1 0 25984 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3010__A2
timestamp 1669390400
transform -1 0 12992 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3016__A2
timestamp 1669390400
transform 1 0 25200 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3016__A3
timestamp 1669390400
transform 1 0 24528 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3018__A1
timestamp 1669390400
transform 1 0 11648 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3018__A2
timestamp 1669390400
transform 1 0 8512 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3018__A3
timestamp 1669390400
transform -1 0 10528 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3020__A1
timestamp 1669390400
transform 1 0 26544 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3021__A1
timestamp 1669390400
transform 1 0 24192 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3021__A2
timestamp 1669390400
transform 1 0 24640 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3022__A1
timestamp 1669390400
transform -1 0 25872 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3023__A2
timestamp 1669390400
transform -1 0 25760 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3023__A3
timestamp 1669390400
transform 1 0 24864 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3025__A1
timestamp 1669390400
transform -1 0 24304 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3028__I
timestamp 1669390400
transform 1 0 21616 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3029__A1
timestamp 1669390400
transform -1 0 22400 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3029__B2
timestamp 1669390400
transform 1 0 27328 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3031__A1
timestamp 1669390400
transform 1 0 26096 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3032__A1
timestamp 1669390400
transform 1 0 25536 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3034__A2
timestamp 1669390400
transform -1 0 38304 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3034__B
timestamp 1669390400
transform 1 0 38528 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3035__I
timestamp 1669390400
transform -1 0 29344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3036__A1
timestamp 1669390400
transform -1 0 26880 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3036__A2
timestamp 1669390400
transform -1 0 26432 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3036__A3
timestamp 1669390400
transform -1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3037__A1
timestamp 1669390400
transform -1 0 24640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3039__I
timestamp 1669390400
transform -1 0 29792 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3040__A1
timestamp 1669390400
transform 1 0 34384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3040__A2
timestamp 1669390400
transform -1 0 28672 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3040__A3
timestamp 1669390400
transform -1 0 34160 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3040__A4
timestamp 1669390400
transform -1 0 35056 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3041__A1
timestamp 1669390400
transform 1 0 32816 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3042__A1
timestamp 1669390400
transform 1 0 33040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3044__I
timestamp 1669390400
transform -1 0 28224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3045__A1
timestamp 1669390400
transform 1 0 32816 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3045__A2
timestamp 1669390400
transform 1 0 30688 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3046__A1
timestamp 1669390400
transform 1 0 29792 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3046__A2
timestamp 1669390400
transform 1 0 27552 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3047__A1
timestamp 1669390400
transform 1 0 32592 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3048__A1
timestamp 1669390400
transform 1 0 30352 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3049__A1
timestamp 1669390400
transform 1 0 33712 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3052__A1
timestamp 1669390400
transform 1 0 30240 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3052__A2
timestamp 1669390400
transform 1 0 33264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3053__A1
timestamp 1669390400
transform 1 0 31136 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3053__A2
timestamp 1669390400
transform 1 0 27552 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3054__A1
timestamp 1669390400
transform -1 0 30352 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3058__A1
timestamp 1669390400
transform 1 0 28784 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3058__A2
timestamp 1669390400
transform -1 0 28560 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3059__A1
timestamp 1669390400
transform -1 0 30800 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3060__A1
timestamp 1669390400
transform 1 0 29680 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3061__A1
timestamp 1669390400
transform 1 0 30128 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3062__A1
timestamp 1669390400
transform 1 0 29120 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3063__A1
timestamp 1669390400
transform 1 0 32144 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3067__I
timestamp 1669390400
transform -1 0 26880 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3068__A1
timestamp 1669390400
transform 1 0 27440 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3068__A2
timestamp 1669390400
transform 1 0 26656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3069__A2
timestamp 1669390400
transform 1 0 27776 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3070__A2
timestamp 1669390400
transform 1 0 29232 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3072__A1
timestamp 1669390400
transform 1 0 25424 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3074__A1
timestamp 1669390400
transform 1 0 25760 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3074__A2
timestamp 1669390400
transform 1 0 26208 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3076__A1
timestamp 1669390400
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3077__A1
timestamp 1669390400
transform 1 0 24192 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3078__A1
timestamp 1669390400
transform -1 0 26096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3079__A1
timestamp 1669390400
transform -1 0 27328 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3083__A1
timestamp 1669390400
transform 1 0 27888 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3083__A2
timestamp 1669390400
transform 1 0 27104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3084__A1
timestamp 1669390400
transform -1 0 24528 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3084__A2
timestamp 1669390400
transform 1 0 26544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3085__A1
timestamp 1669390400
transform -1 0 29232 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3085__A2
timestamp 1669390400
transform 1 0 26992 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3087__A1
timestamp 1669390400
transform -1 0 24976 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3089__A1
timestamp 1669390400
transform 1 0 26320 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3089__B
timestamp 1669390400
transform -1 0 25088 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3090__A1
timestamp 1669390400
transform -1 0 24192 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3090__A2
timestamp 1669390400
transform -1 0 25536 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3092__A1
timestamp 1669390400
transform -1 0 23968 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3093__A1
timestamp 1669390400
transform 1 0 22960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3095__A2
timestamp 1669390400
transform -1 0 24752 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3097__I
timestamp 1669390400
transform -1 0 25984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3098__A1
timestamp 1669390400
transform -1 0 25536 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3098__A2
timestamp 1669390400
transform -1 0 26096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3099__A1
timestamp 1669390400
transform -1 0 23408 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3100__A2
timestamp 1669390400
transform -1 0 24304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3101__A1
timestamp 1669390400
transform -1 0 19936 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3104__A1
timestamp 1669390400
transform 1 0 25424 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3104__B
timestamp 1669390400
transform 1 0 25648 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3105__A1
timestamp 1669390400
transform -1 0 28672 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3105__A3
timestamp 1669390400
transform 1 0 28000 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3107__A1
timestamp 1669390400
transform 1 0 23408 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3107__B
timestamp 1669390400
transform 1 0 22512 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3108__A1
timestamp 1669390400
transform -1 0 22960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3108__A2
timestamp 1669390400
transform -1 0 23856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3113__A1
timestamp 1669390400
transform -1 0 21392 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3115__A1
timestamp 1669390400
transform 1 0 19600 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3117__I
timestamp 1669390400
transform -1 0 23632 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3118__A2
timestamp 1669390400
transform 1 0 25088 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3120__A1
timestamp 1669390400
transform 1 0 23520 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3120__B
timestamp 1669390400
transform 1 0 20832 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3121__A1
timestamp 1669390400
transform 1 0 23968 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3121__A2
timestamp 1669390400
transform 1 0 22960 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3125__A2
timestamp 1669390400
transform 1 0 24192 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3129__A1
timestamp 1669390400
transform 1 0 24752 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3131__I
timestamp 1669390400
transform 1 0 23408 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3132__A2
timestamp 1669390400
transform -1 0 26544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3134__A1
timestamp 1669390400
transform 1 0 21616 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3135__A1
timestamp 1669390400
transform 1 0 23184 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3139__A1
timestamp 1669390400
transform -1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3139__A2
timestamp 1669390400
transform 1 0 25872 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3142__A1
timestamp 1669390400
transform 1 0 20384 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3145__A1
timestamp 1669390400
transform 1 0 20832 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3146__A1
timestamp 1669390400
transform -1 0 18480 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3148__A1
timestamp 1669390400
transform 1 0 11088 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3148__A2
timestamp 1669390400
transform -1 0 11760 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3150__A1
timestamp 1669390400
transform 1 0 11312 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3150__A2
timestamp 1669390400
transform 1 0 10640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3154__A1
timestamp 1669390400
transform 1 0 4928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3156__I
timestamp 1669390400
transform 1 0 4816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3157__A1
timestamp 1669390400
transform -1 0 5152 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3161__A1
timestamp 1669390400
transform 1 0 7616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3161__A2
timestamp 1669390400
transform -1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3163__A1
timestamp 1669390400
transform 1 0 5600 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3163__A2
timestamp 1669390400
transform 1 0 5152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3164__A1
timestamp 1669390400
transform -1 0 7392 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3166__A1
timestamp 1669390400
transform 1 0 8624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3166__A2
timestamp 1669390400
transform 1 0 7168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3166__A3
timestamp 1669390400
transform 1 0 6720 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3167__A1
timestamp 1669390400
transform -1 0 8624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3169__A1
timestamp 1669390400
transform 1 0 8176 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3169__A2
timestamp 1669390400
transform 1 0 5824 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3169__A3
timestamp 1669390400
transform -1 0 6496 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3169__A4
timestamp 1669390400
transform -1 0 4704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3170__A1
timestamp 1669390400
transform -1 0 2464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3172__A1
timestamp 1669390400
transform 1 0 8736 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3173__A1
timestamp 1669390400
transform -1 0 1904 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3175__A1
timestamp 1669390400
transform -1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3176__A1
timestamp 1669390400
transform -1 0 1904 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3177__A1
timestamp 1669390400
transform -1 0 14672 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3177__A2
timestamp 1669390400
transform -1 0 13776 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3189__A1
timestamp 1669390400
transform -1 0 15792 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3189__A2
timestamp 1669390400
transform -1 0 15120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3191__A1
timestamp 1669390400
transform -1 0 16240 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3191__A2
timestamp 1669390400
transform 1 0 18032 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3192__A1
timestamp 1669390400
transform -1 0 17808 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3194__A1
timestamp 1669390400
transform -1 0 15344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3195__A1
timestamp 1669390400
transform 1 0 17808 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3197__A2
timestamp 1669390400
transform 1 0 19152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3197__B
timestamp 1669390400
transform -1 0 19712 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3198__A1
timestamp 1669390400
transform -1 0 19600 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3201__CLK
timestamp 1669390400
transform -1 0 16912 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3201__RN
timestamp 1669390400
transform 1 0 22064 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3202__CLK
timestamp 1669390400
transform 1 0 13552 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3202__D
timestamp 1669390400
transform 1 0 14448 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3202__RN
timestamp 1669390400
transform 1 0 14000 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3203__CLK
timestamp 1669390400
transform 1 0 9632 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3203__D
timestamp 1669390400
transform -1 0 14336 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3203__RN
timestamp 1669390400
transform 1 0 14336 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3204__CLK
timestamp 1669390400
transform 1 0 17584 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3204__D
timestamp 1669390400
transform -1 0 18704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3204__RN
timestamp 1669390400
transform 1 0 18032 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3205__CLK
timestamp 1669390400
transform 1 0 13552 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3205__D
timestamp 1669390400
transform -1 0 13104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3205__RN
timestamp 1669390400
transform 1 0 14000 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3206__CLK
timestamp 1669390400
transform 1 0 17584 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3206__D
timestamp 1669390400
transform 1 0 18480 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3206__RN
timestamp 1669390400
transform 1 0 18032 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3207__CLK
timestamp 1669390400
transform 1 0 10864 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3207__D
timestamp 1669390400
transform 1 0 16240 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3207__RN
timestamp 1669390400
transform 1 0 14560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3208__CLK
timestamp 1669390400
transform 1 0 14448 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3208__RN
timestamp 1669390400
transform 1 0 19264 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3209__CLK
timestamp 1669390400
transform 1 0 14896 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3209__RN
timestamp 1669390400
transform -1 0 18256 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3210__CLK
timestamp 1669390400
transform 1 0 15120 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3210__RN
timestamp 1669390400
transform -1 0 15792 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3211__CLK
timestamp 1669390400
transform 1 0 19040 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3211__RN
timestamp 1669390400
transform 1 0 19488 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3212__CLK
timestamp 1669390400
transform 1 0 19152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3212__RN
timestamp 1669390400
transform 1 0 18704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3213__CLK
timestamp 1669390400
transform 1 0 14784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3213__RN
timestamp 1669390400
transform 1 0 19264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3214__CLK
timestamp 1669390400
transform 1 0 14896 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3214__RN
timestamp 1669390400
transform 1 0 19600 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3215__CLK
timestamp 1669390400
transform 1 0 14112 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3215__RN
timestamp 1669390400
transform 1 0 19152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3216__CLK
timestamp 1669390400
transform 1 0 14896 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3216__RN
timestamp 1669390400
transform 1 0 19376 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3217__CLK
timestamp 1669390400
transform 1 0 13552 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3217__RN
timestamp 1669390400
transform 1 0 14000 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3218__CLK
timestamp 1669390400
transform -1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3218__RN
timestamp 1669390400
transform -1 0 8176 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3219__CLK
timestamp 1669390400
transform 1 0 5600 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3219__RN
timestamp 1669390400
transform 1 0 12320 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3220__CLK
timestamp 1669390400
transform 1 0 10528 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3220__RN
timestamp 1669390400
transform 1 0 10976 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3221__CLK
timestamp 1669390400
transform -1 0 9744 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3221__RN
timestamp 1669390400
transform -1 0 10192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3222__CLK
timestamp 1669390400
transform 1 0 7952 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3222__RN
timestamp 1669390400
transform -1 0 7728 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3223__CLK
timestamp 1669390400
transform 1 0 8848 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3223__RN
timestamp 1669390400
transform 1 0 13664 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3224__CLK
timestamp 1669390400
transform 1 0 9632 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3224__RN
timestamp 1669390400
transform 1 0 10080 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3225__CLK
timestamp 1669390400
transform 1 0 9632 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3225__RN
timestamp 1669390400
transform -1 0 3472 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3226__CLK
timestamp 1669390400
transform -1 0 5152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3226__RN
timestamp 1669390400
transform 1 0 13552 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3227__CLK
timestamp 1669390400
transform 1 0 6384 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3227__RN
timestamp 1669390400
transform 1 0 12880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3228__CLK
timestamp 1669390400
transform 1 0 6832 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3228__RN
timestamp 1669390400
transform 1 0 11872 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3229__CLK
timestamp 1669390400
transform 1 0 10080 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3229__RN
timestamp 1669390400
transform 1 0 7728 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3230__CLK
timestamp 1669390400
transform 1 0 15344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3230__RN
timestamp 1669390400
transform 1 0 14000 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3231__CLK
timestamp 1669390400
transform 1 0 17584 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3231__RN
timestamp 1669390400
transform 1 0 18032 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3232__CLK
timestamp 1669390400
transform 1 0 15792 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3232__RN
timestamp 1669390400
transform 1 0 19712 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3233__CLK
timestamp 1669390400
transform 1 0 14896 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3233__RN
timestamp 1669390400
transform 1 0 19824 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1669390400
transform -1 0 11312 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_0__f_clk_I
timestamp 1669390400
transform 1 0 13552 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_1__f_clk_I
timestamp 1669390400
transform -1 0 16464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_2__f_clk_I
timestamp 1669390400
transform 1 0 7280 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_3__f_clk_I
timestamp 1669390400
transform 1 0 18480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout9_I
timestamp 1669390400
transform -1 0 17808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout10_I
timestamp 1669390400
transform 1 0 20160 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout11_I
timestamp 1669390400
transform -1 0 19824 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1669390400
transform -1 0 27328 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1669390400
transform -1 0 38640 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1669390400
transform 1 0 48720 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1669390400
transform 1 0 56560 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1669390400
transform -1 0 12992 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output6_I
timestamp 1669390400
transform 1 0 49840 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output8_I
timestamp 1669390400
transform 1 0 29792 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1568 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 3360 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 4256 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 4704 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5152 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37
timestamp 1669390400
transform 1 0 5488 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50
timestamp 1669390400
transform 1 0 6944 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54
timestamp 1669390400
transform 1 0 7392 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58
timestamp 1669390400
transform 1 0 7840 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66
timestamp 1669390400
transform 1 0 8736 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72
timestamp 1669390400
transform 1 0 9408 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75
timestamp 1669390400
transform 1 0 9744 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_79
timestamp 1669390400
transform 1 0 10192 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_95
timestamp 1669390400
transform 1 0 11984 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99
timestamp 1669390400
transform 1 0 12432 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_101
timestamp 1669390400
transform 1 0 12656 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1669390400
transform 1 0 12992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_107
timestamp 1669390400
transform 1 0 13328 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_124
timestamp 1669390400
transform 1 0 15232 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_132
timestamp 1669390400
transform 1 0 16128 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_135
timestamp 1669390400
transform 1 0 16464 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1669390400
transform 1 0 16912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_142
timestamp 1669390400
transform 1 0 17248 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_144
timestamp 1669390400
transform 1 0 17472 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_147
timestamp 1669390400
transform 1 0 17808 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_151
timestamp 1669390400
transform 1 0 18256 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_167
timestamp 1669390400
transform 1 0 20048 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_177
timestamp 1669390400
transform 1 0 21168 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_183
timestamp 1669390400
transform 1 0 21840 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_187
timestamp 1669390400
transform 1 0 22288 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_193
timestamp 1669390400
transform 1 0 22960 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_197
timestamp 1669390400
transform 1 0 23408 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_201
timestamp 1669390400
transform 1 0 23856 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_205
timestamp 1669390400
transform 1 0 24304 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1669390400
transform 1 0 24752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_212
timestamp 1669390400
transform 1 0 25088 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_216
timestamp 1669390400
transform 1 0 25536 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_220
timestamp 1669390400
transform 1 0 25984 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_224
timestamp 1669390400
transform 1 0 26432 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_228
timestamp 1669390400
transform 1 0 26880 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_232
timestamp 1669390400
transform 1 0 27328 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_236
timestamp 1669390400
transform 1 0 27776 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_240
timestamp 1669390400
transform 1 0 28224 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_244
timestamp 1669390400
transform 1 0 28672 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_247
timestamp 1669390400
transform 1 0 29008 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_250
timestamp 1669390400
transform 1 0 29344 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_254
timestamp 1669390400
transform 1 0 29792 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_264
timestamp 1669390400
transform 1 0 30912 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_278
timestamp 1669390400
transform 1 0 32480 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_282
timestamp 1669390400
transform 1 0 32928 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_285
timestamp 1669390400
transform 1 0 33264 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_289
timestamp 1669390400
transform 1 0 33712 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_293
timestamp 1669390400
transform 1 0 34160 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_297
timestamp 1669390400
transform 1 0 34608 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_301
timestamp 1669390400
transform 1 0 35056 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_305
timestamp 1669390400
transform 1 0 35504 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_309
timestamp 1669390400
transform 1 0 35952 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_313
timestamp 1669390400
transform 1 0 36400 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_317
timestamp 1669390400
transform 1 0 36848 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_326
timestamp 1669390400
transform 1 0 37856 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_330
timestamp 1669390400
transform 1 0 38304 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_333
timestamp 1669390400
transform 1 0 38640 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_343
timestamp 1669390400
transform 1 0 39760 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_349
timestamp 1669390400
transform 1 0 40432 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_352
timestamp 1669390400
transform 1 0 40768 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_358
timestamp 1669390400
transform 1 0 41440 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_365
timestamp 1669390400
transform 1 0 42224 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_381
timestamp 1669390400
transform 1 0 44016 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_387
timestamp 1669390400
transform 1 0 44688 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_403
timestamp 1669390400
transform 1 0 46480 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_419
timestamp 1669390400
transform 1 0 48272 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_422
timestamp 1669390400
transform 1 0 48608 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_425
timestamp 1669390400
transform 1 0 48944 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_441
timestamp 1669390400
transform 1 0 50736 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_449
timestamp 1669390400
transform 1 0 51632 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_453
timestamp 1669390400
transform 1 0 52080 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_457
timestamp 1669390400
transform 1 0 52528 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_473
timestamp 1669390400
transform 1 0 54320 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_487
timestamp 1669390400
transform 1 0 55888 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_489
timestamp 1669390400
transform 1 0 56112 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_492
timestamp 1669390400
transform 1 0 56448 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_495
timestamp 1669390400
transform 1 0 56784 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_511
timestamp 1669390400
transform 1 0 58576 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_2 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1568 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_34
timestamp 1669390400
transform 1 0 5152 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1669390400
transform 1 0 9184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_73
timestamp 1669390400
transform 1 0 9520 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_84
timestamp 1669390400
transform 1 0 10752 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_88
timestamp 1669390400
transform 1 0 11200 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_140
timestamp 1669390400
transform 1 0 17024 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_144
timestamp 1669390400
transform 1 0 17472 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_179
timestamp 1669390400
transform 1 0 21392 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_193
timestamp 1669390400
transform 1 0 22960 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_200
timestamp 1669390400
transform 1 0 23744 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_204
timestamp 1669390400
transform 1 0 24192 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_208
timestamp 1669390400
transform 1 0 24640 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1669390400
transform 1 0 25088 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_215
timestamp 1669390400
transform 1 0 25424 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_224
timestamp 1669390400
transform 1 0 26432 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_226
timestamp 1669390400
transform 1 0 26656 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_235
timestamp 1669390400
transform 1 0 27664 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_245
timestamp 1669390400
transform 1 0 28784 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_255
timestamp 1669390400
transform 1 0 29904 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_261
timestamp 1669390400
transform 1 0 30576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_265
timestamp 1669390400
transform 1 0 31024 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_279
timestamp 1669390400
transform 1 0 32592 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_283
timestamp 1669390400
transform 1 0 33040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_286
timestamp 1669390400
transform 1 0 33376 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_293
timestamp 1669390400
transform 1 0 34160 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_297
timestamp 1669390400
transform 1 0 34608 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_307
timestamp 1669390400
transform 1 0 35728 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_313
timestamp 1669390400
transform 1 0 36400 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_327
timestamp 1669390400
transform 1 0 37968 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_331
timestamp 1669390400
transform 1 0 38416 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_341
timestamp 1669390400
transform 1 0 39536 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_354
timestamp 1669390400
transform 1 0 40992 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_357
timestamp 1669390400
transform 1 0 41328 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_371
timestamp 1669390400
transform 1 0 42896 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_375
timestamp 1669390400
transform 1 0 43344 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_379
timestamp 1669390400
transform 1 0 43792 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_392
timestamp 1669390400
transform 1 0 45248 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_399
timestamp 1669390400
transform 1 0 46032 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_415
timestamp 1669390400
transform 1 0 47824 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_424
timestamp 1669390400
transform 1 0 48832 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_428 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 49280 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_492
timestamp 1669390400
transform 1 0 56448 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_496
timestamp 1669390400
transform 1 0 56896 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_499
timestamp 1669390400
transform 1 0 57232 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_507
timestamp 1669390400
transform 1 0 58128 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_511
timestamp 1669390400
transform 1 0 58576 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1669390400
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1669390400
transform 1 0 5152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_37
timestamp 1669390400
transform 1 0 5488 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_51
timestamp 1669390400
transform 1 0 7056 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1669390400
transform 1 0 13104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_108
timestamp 1669390400
transform 1 0 13440 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_111
timestamp 1669390400
transform 1 0 13776 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_113
timestamp 1669390400
transform 1 0 14000 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_116
timestamp 1669390400
transform 1 0 14336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_120
timestamp 1669390400
transform 1 0 14784 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_123
timestamp 1669390400
transform 1 0 15120 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_159
timestamp 1669390400
transform 1 0 19152 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_163
timestamp 1669390400
transform 1 0 19600 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_166
timestamp 1669390400
transform 1 0 19936 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1669390400
transform 1 0 21056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_179
timestamp 1669390400
transform 1 0 21392 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_203
timestamp 1669390400
transform 1 0 24080 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_207
timestamp 1669390400
transform 1 0 24528 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_220
timestamp 1669390400
transform 1 0 25984 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_222
timestamp 1669390400
transform 1 0 26208 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_225
timestamp 1669390400
transform 1 0 26544 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_237
timestamp 1669390400
transform 1 0 27888 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_247
timestamp 1669390400
transform 1 0 29008 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_250
timestamp 1669390400
transform 1 0 29344 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_289
timestamp 1669390400
transform 1 0 33712 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_291
timestamp 1669390400
transform 1 0 33936 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_294
timestamp 1669390400
transform 1 0 34272 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_308
timestamp 1669390400
transform 1 0 35840 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_318
timestamp 1669390400
transform 1 0 36960 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_321
timestamp 1669390400
transform 1 0 37296 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_334
timestamp 1669390400
transform 1 0 38752 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_346
timestamp 1669390400
transform 1 0 40096 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_350
timestamp 1669390400
transform 1 0 40544 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_352
timestamp 1669390400
transform 1 0 40768 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_364
timestamp 1669390400
transform 1 0 42112 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_374
timestamp 1669390400
transform 1 0 43232 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_376
timestamp 1669390400
transform 1 0 43456 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_389
timestamp 1669390400
transform 1 0 44912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_392
timestamp 1669390400
transform 1 0 45248 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_399
timestamp 1669390400
transform 1 0 46032 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_407
timestamp 1669390400
transform 1 0 46928 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_420
timestamp 1669390400
transform 1 0 48384 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_432
timestamp 1669390400
transform 1 0 49728 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_448
timestamp 1669390400
transform 1 0 51520 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_456
timestamp 1669390400
transform 1 0 52416 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_460
timestamp 1669390400
transform 1 0 52864 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_463
timestamp 1669390400
transform 1 0 53200 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_495
timestamp 1669390400
transform 1 0 56784 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_511
timestamp 1669390400
transform 1 0 58576 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_2
timestamp 1669390400
transform 1 0 1568 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_34
timestamp 1669390400
transform 1 0 5152 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1669390400
transform 1 0 9184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_73
timestamp 1669390400
transform 1 0 9520 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_76
timestamp 1669390400
transform 1 0 9856 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_114
timestamp 1669390400
transform 1 0 14112 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_118
timestamp 1669390400
transform 1 0 14560 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_122
timestamp 1669390400
transform 1 0 15008 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_125
timestamp 1669390400
transform 1 0 15344 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_129
timestamp 1669390400
transform 1 0 15792 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_139
timestamp 1669390400
transform 1 0 16912 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1669390400
transform 1 0 17136 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_144
timestamp 1669390400
transform 1 0 17472 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_179
timestamp 1669390400
transform 1 0 21392 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_189
timestamp 1669390400
transform 1 0 22512 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_200
timestamp 1669390400
transform 1 0 23744 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_210
timestamp 1669390400
transform 1 0 24864 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1669390400
transform 1 0 25088 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_215
timestamp 1669390400
transform 1 0 25424 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_221
timestamp 1669390400
transform 1 0 26096 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_231
timestamp 1669390400
transform 1 0 27216 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_239
timestamp 1669390400
transform 1 0 28112 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_241
timestamp 1669390400
transform 1 0 28336 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_244
timestamp 1669390400
transform 1 0 28672 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_252
timestamp 1669390400
transform 1 0 29568 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_256
timestamp 1669390400
transform 1 0 30016 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_259
timestamp 1669390400
transform 1 0 30352 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_266
timestamp 1669390400
transform 1 0 31136 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_280
timestamp 1669390400
transform 1 0 32704 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_286
timestamp 1669390400
transform 1 0 33376 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_293
timestamp 1669390400
transform 1 0 34160 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_297
timestamp 1669390400
transform 1 0 34608 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_310
timestamp 1669390400
transform 1 0 36064 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_324
timestamp 1669390400
transform 1 0 37632 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_332
timestamp 1669390400
transform 1 0 38528 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_336
timestamp 1669390400
transform 1 0 38976 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_347
timestamp 1669390400
transform 1 0 40208 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_357
timestamp 1669390400
transform 1 0 41328 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_366
timestamp 1669390400
transform 1 0 42336 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_376
timestamp 1669390400
transform 1 0 43456 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_388
timestamp 1669390400
transform 1 0 44800 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_395
timestamp 1669390400
transform 1 0 45584 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_404
timestamp 1669390400
transform 1 0 46592 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_419
timestamp 1669390400
transform 1 0 48272 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_423
timestamp 1669390400
transform 1 0 48720 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_425
timestamp 1669390400
transform 1 0 48944 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_428
timestamp 1669390400
transform 1 0 49280 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_492
timestamp 1669390400
transform 1 0 56448 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_496
timestamp 1669390400
transform 1 0 56896 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_499
timestamp 1669390400
transform 1 0 57232 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_507
timestamp 1669390400
transform 1 0 58128 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_511
timestamp 1669390400
transform 1 0 58576 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_2
timestamp 1669390400
transform 1 0 1568 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_18
timestamp 1669390400
transform 1 0 3360 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_26
timestamp 1669390400
transform 1 0 4256 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_28
timestamp 1669390400
transform 1 0 4480 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1669390400
transform 1 0 5152 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_37
timestamp 1669390400
transform 1 0 5488 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_40
timestamp 1669390400
transform 1 0 5824 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_44
timestamp 1669390400
transform 1 0 6272 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_51
timestamp 1669390400
transform 1 0 7056 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_57
timestamp 1669390400
transform 1 0 7728 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_61
timestamp 1669390400
transform 1 0 8176 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_65
timestamp 1669390400
transform 1 0 8624 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_69
timestamp 1669390400
transform 1 0 9072 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1669390400
transform 1 0 13104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_108
timestamp 1669390400
transform 1 0 13440 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_111
timestamp 1669390400
transform 1 0 13776 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_115
timestamp 1669390400
transform 1 0 14224 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_119
timestamp 1669390400
transform 1 0 14672 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_121
timestamp 1669390400
transform 1 0 14896 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_158
timestamp 1669390400
transform 1 0 19040 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_166
timestamp 1669390400
transform 1 0 19936 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_174
timestamp 1669390400
transform 1 0 20832 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1669390400
transform 1 0 21056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_179
timestamp 1669390400
transform 1 0 21392 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_186
timestamp 1669390400
transform 1 0 22176 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_188
timestamp 1669390400
transform 1 0 22400 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_191
timestamp 1669390400
transform 1 0 22736 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_195
timestamp 1669390400
transform 1 0 23184 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_199
timestamp 1669390400
transform 1 0 23632 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_209
timestamp 1669390400
transform 1 0 24752 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_213
timestamp 1669390400
transform 1 0 25200 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_216
timestamp 1669390400
transform 1 0 25536 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_232
timestamp 1669390400
transform 1 0 27328 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_236
timestamp 1669390400
transform 1 0 27776 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_240
timestamp 1669390400
transform 1 0 28224 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_246
timestamp 1669390400
transform 1 0 28896 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_250
timestamp 1669390400
transform 1 0 29344 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_256
timestamp 1669390400
transform 1 0 30016 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_260
timestamp 1669390400
transform 1 0 30464 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_264
timestamp 1669390400
transform 1 0 30912 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_268
timestamp 1669390400
transform 1 0 31360 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_277
timestamp 1669390400
transform 1 0 32368 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_287
timestamp 1669390400
transform 1 0 33488 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_291
timestamp 1669390400
transform 1 0 33936 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_307
timestamp 1669390400
transform 1 0 35728 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_311
timestamp 1669390400
transform 1 0 36176 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_321
timestamp 1669390400
transform 1 0 37296 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_353
timestamp 1669390400
transform 1 0 40880 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_369
timestamp 1669390400
transform 1 0 42672 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_377
timestamp 1669390400
transform 1 0 43568 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_380
timestamp 1669390400
transform 1 0 43904 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_388
timestamp 1669390400
transform 1 0 44800 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_392
timestamp 1669390400
transform 1 0 45248 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_395
timestamp 1669390400
transform 1 0 45584 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_459
timestamp 1669390400
transform 1 0 52752 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_463
timestamp 1669390400
transform 1 0 53200 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_481
timestamp 1669390400
transform 1 0 55216 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_485
timestamp 1669390400
transform 1 0 55664 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_501
timestamp 1669390400
transform 1 0 57456 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_509
timestamp 1669390400
transform 1 0 58352 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_2
timestamp 1669390400
transform 1 0 1568 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_36
timestamp 1669390400
transform 1 0 5376 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_38
timestamp 1669390400
transform 1 0 5600 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_45
timestamp 1669390400
transform 1 0 6384 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_53
timestamp 1669390400
transform 1 0 7280 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1669390400
transform 1 0 9184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_73
timestamp 1669390400
transform 1 0 9520 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_108
timestamp 1669390400
transform 1 0 13440 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_112
timestamp 1669390400
transform 1 0 13888 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_128
timestamp 1669390400
transform 1 0 15680 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_136
timestamp 1669390400
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_140
timestamp 1669390400
transform 1 0 17024 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_144
timestamp 1669390400
transform 1 0 17472 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_152
timestamp 1669390400
transform 1 0 18368 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_154
timestamp 1669390400
transform 1 0 18592 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_157
timestamp 1669390400
transform 1 0 18928 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_161
timestamp 1669390400
transform 1 0 19376 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_165
timestamp 1669390400
transform 1 0 19824 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_190
timestamp 1669390400
transform 1 0 22624 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_199
timestamp 1669390400
transform 1 0 23632 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_203
timestamp 1669390400
transform 1 0 24080 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_212
timestamp 1669390400
transform 1 0 25088 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_215
timestamp 1669390400
transform 1 0 25424 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_222
timestamp 1669390400
transform 1 0 26208 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_228
timestamp 1669390400
transform 1 0 26880 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_236
timestamp 1669390400
transform 1 0 27776 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_238
timestamp 1669390400
transform 1 0 28000 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_247
timestamp 1669390400
transform 1 0 29008 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_251
timestamp 1669390400
transform 1 0 29456 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_260
timestamp 1669390400
transform 1 0 30464 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_264
timestamp 1669390400
transform 1 0 30912 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_277
timestamp 1669390400
transform 1 0 32368 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_281
timestamp 1669390400
transform 1 0 32816 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_283
timestamp 1669390400
transform 1 0 33040 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_286
timestamp 1669390400
transform 1 0 33376 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_289
timestamp 1669390400
transform 1 0 33712 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_293
timestamp 1669390400
transform 1 0 34160 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_295
timestamp 1669390400
transform 1 0 34384 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_302
timestamp 1669390400
transform 1 0 35168 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_318
timestamp 1669390400
transform 1 0 36960 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_326
timestamp 1669390400
transform 1 0 37856 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_334
timestamp 1669390400
transform 1 0 38752 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_338
timestamp 1669390400
transform 1 0 39200 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_348
timestamp 1669390400
transform 1 0 40320 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_352
timestamp 1669390400
transform 1 0 40768 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_354
timestamp 1669390400
transform 1 0 40992 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_357
timestamp 1669390400
transform 1 0 41328 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_360
timestamp 1669390400
transform 1 0 41664 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_364
timestamp 1669390400
transform 1 0 42112 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_378
timestamp 1669390400
transform 1 0 43680 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_382
timestamp 1669390400
transform 1 0 44128 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_386
timestamp 1669390400
transform 1 0 44576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_390
timestamp 1669390400
transform 1 0 45024 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_392
timestamp 1669390400
transform 1 0 45248 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_395
timestamp 1669390400
transform 1 0 45584 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_409
timestamp 1669390400
transform 1 0 47152 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_425
timestamp 1669390400
transform 1 0 48944 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_428
timestamp 1669390400
transform 1 0 49280 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_432
timestamp 1669390400
transform 1 0 49728 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_446
timestamp 1669390400
transform 1 0 51296 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_454
timestamp 1669390400
transform 1 0 52192 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_458
timestamp 1669390400
transform 1 0 52640 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_460
timestamp 1669390400
transform 1 0 52864 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_466
timestamp 1669390400
transform 1 0 53536 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_470
timestamp 1669390400
transform 1 0 53984 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_477
timestamp 1669390400
transform 1 0 54768 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_489
timestamp 1669390400
transform 1 0 56112 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_499
timestamp 1669390400
transform 1 0 57232 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_507
timestamp 1669390400
transform 1 0 58128 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_511
timestamp 1669390400
transform 1 0 58576 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1669390400
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1669390400
transform 1 0 5152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_37
timestamp 1669390400
transform 1 0 5488 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_45
timestamp 1669390400
transform 1 0 6384 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_47
timestamp 1669390400
transform 1 0 6608 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_50
timestamp 1669390400
transform 1 0 6944 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_54
timestamp 1669390400
transform 1 0 7392 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_63
timestamp 1669390400
transform 1 0 8400 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_67
timestamp 1669390400
transform 1 0 8848 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1669390400
transform 1 0 13104 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_108
timestamp 1669390400
transform 1 0 13440 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_111
timestamp 1669390400
transform 1 0 13776 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_115
timestamp 1669390400
transform 1 0 14224 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_119
timestamp 1669390400
transform 1 0 14672 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_156
timestamp 1669390400
transform 1 0 18816 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_160
timestamp 1669390400
transform 1 0 19264 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_164
timestamp 1669390400
transform 1 0 19712 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_172
timestamp 1669390400
transform 1 0 20608 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1669390400
transform 1 0 21056 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_179
timestamp 1669390400
transform 1 0 21392 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_186
timestamp 1669390400
transform 1 0 22176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_198
timestamp 1669390400
transform 1 0 23520 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_200
timestamp 1669390400
transform 1 0 23744 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_213
timestamp 1669390400
transform 1 0 25200 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_217
timestamp 1669390400
transform 1 0 25648 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_227
timestamp 1669390400
transform 1 0 26768 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_247
timestamp 1669390400
transform 1 0 29008 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_250
timestamp 1669390400
transform 1 0 29344 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_256
timestamp 1669390400
transform 1 0 30016 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_263
timestamp 1669390400
transform 1 0 30800 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_265
timestamp 1669390400
transform 1 0 31024 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_268
timestamp 1669390400
transform 1 0 31360 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_270
timestamp 1669390400
transform 1 0 31584 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_279
timestamp 1669390400
transform 1 0 32592 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_283
timestamp 1669390400
transform 1 0 33040 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_287
timestamp 1669390400
transform 1 0 33488 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_299
timestamp 1669390400
transform 1 0 34832 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_307
timestamp 1669390400
transform 1 0 35728 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_311
timestamp 1669390400
transform 1 0 36176 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_321
timestamp 1669390400
transform 1 0 37296 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_334
timestamp 1669390400
transform 1 0 38752 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_346
timestamp 1669390400
transform 1 0 40096 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_356
timestamp 1669390400
transform 1 0 41216 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_360
timestamp 1669390400
transform 1 0 41664 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_364
timestamp 1669390400
transform 1 0 42112 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_375
timestamp 1669390400
transform 1 0 43344 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_389
timestamp 1669390400
transform 1 0 44912 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_392
timestamp 1669390400
transform 1 0 45248 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_396
timestamp 1669390400
transform 1 0 45696 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_400
timestamp 1669390400
transform 1 0 46144 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_417
timestamp 1669390400
transform 1 0 48048 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_421
timestamp 1669390400
transform 1 0 48496 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_434
timestamp 1669390400
transform 1 0 49952 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_436
timestamp 1669390400
transform 1 0 50176 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_460
timestamp 1669390400
transform 1 0 52864 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_463
timestamp 1669390400
transform 1 0 53200 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_480
timestamp 1669390400
transform 1 0 55104 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_482
timestamp 1669390400
transform 1 0 55328 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_501
timestamp 1669390400
transform 1 0 57456 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_505
timestamp 1669390400
transform 1 0 57904 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_2
timestamp 1669390400
transform 1 0 1568 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_18
timestamp 1669390400
transform 1 0 3360 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_22
timestamp 1669390400
transform 1 0 3808 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_24
timestamp 1669390400
transform 1 0 4032 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_29
timestamp 1669390400
transform 1 0 4592 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_33
timestamp 1669390400
transform 1 0 5040 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_69
timestamp 1669390400
transform 1 0 9072 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_73
timestamp 1669390400
transform 1 0 9520 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_80
timestamp 1669390400
transform 1 0 10304 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_84
timestamp 1669390400
transform 1 0 10752 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_88
timestamp 1669390400
transform 1 0 11200 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_96
timestamp 1669390400
transform 1 0 12096 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_100
timestamp 1669390400
transform 1 0 12544 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_102
timestamp 1669390400
transform 1 0 12768 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_105
timestamp 1669390400
transform 1 0 13104 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1669390400
transform 1 0 17136 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_144
timestamp 1669390400
transform 1 0 17472 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_147
timestamp 1669390400
transform 1 0 17808 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_151
timestamp 1669390400
transform 1 0 18256 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_155
timestamp 1669390400
transform 1 0 18704 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_171
timestamp 1669390400
transform 1 0 20496 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_175
timestamp 1669390400
transform 1 0 20944 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_179
timestamp 1669390400
transform 1 0 21392 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_186
timestamp 1669390400
transform 1 0 22176 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_196
timestamp 1669390400
transform 1 0 23296 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_200
timestamp 1669390400
transform 1 0 23744 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_204
timestamp 1669390400
transform 1 0 24192 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1669390400
transform 1 0 25088 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_215
timestamp 1669390400
transform 1 0 25424 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_219
timestamp 1669390400
transform 1 0 25872 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_221
timestamp 1669390400
transform 1 0 26096 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_224
timestamp 1669390400
transform 1 0 26432 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_228
timestamp 1669390400
transform 1 0 26880 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_232
timestamp 1669390400
transform 1 0 27328 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_236
timestamp 1669390400
transform 1 0 27776 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_244
timestamp 1669390400
transform 1 0 28672 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_250
timestamp 1669390400
transform 1 0 29344 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_266
timestamp 1669390400
transform 1 0 31136 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_274
timestamp 1669390400
transform 1 0 32032 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_282
timestamp 1669390400
transform 1 0 32928 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_286
timestamp 1669390400
transform 1 0 33376 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_288
timestamp 1669390400
transform 1 0 33600 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_291
timestamp 1669390400
transform 1 0 33936 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_295
timestamp 1669390400
transform 1 0 34384 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_298
timestamp 1669390400
transform 1 0 34720 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_302
timestamp 1669390400
transform 1 0 35168 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_308
timestamp 1669390400
transform 1 0 35840 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_314
timestamp 1669390400
transform 1 0 36512 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_328
timestamp 1669390400
transform 1 0 38080 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_332
timestamp 1669390400
transform 1 0 38528 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_339
timestamp 1669390400
transform 1 0 39312 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_341
timestamp 1669390400
transform 1 0 39536 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_354
timestamp 1669390400
transform 1 0 40992 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_357
timestamp 1669390400
transform 1 0 41328 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_366
timestamp 1669390400
transform 1 0 42336 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_376
timestamp 1669390400
transform 1 0 43456 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_382
timestamp 1669390400
transform 1 0 44128 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_392
timestamp 1669390400
transform 1 0 45248 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_396
timestamp 1669390400
transform 1 0 45696 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_406
timestamp 1669390400
transform 1 0 46816 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_416
timestamp 1669390400
transform 1 0 47936 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_424
timestamp 1669390400
transform 1 0 48832 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_428
timestamp 1669390400
transform 1 0 49280 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_435
timestamp 1669390400
transform 1 0 50064 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_445
timestamp 1669390400
transform 1 0 51184 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_452
timestamp 1669390400
transform 1 0 51968 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_456
timestamp 1669390400
transform 1 0 52416 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_469
timestamp 1669390400
transform 1 0 53872 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_479
timestamp 1669390400
transform 1 0 54992 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_483
timestamp 1669390400
transform 1 0 55440 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_496
timestamp 1669390400
transform 1 0 56896 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_499
timestamp 1669390400
transform 1 0 57232 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_510
timestamp 1669390400
transform 1 0 58464 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_512
timestamp 1669390400
transform 1 0 58688 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_2
timestamp 1669390400
transform 1 0 1568 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_18
timestamp 1669390400
transform 1 0 3360 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1669390400
transform 1 0 5152 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_37
timestamp 1669390400
transform 1 0 5488 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_44
timestamp 1669390400
transform 1 0 6272 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_60
timestamp 1669390400
transform 1 0 8064 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_69
timestamp 1669390400
transform 1 0 9072 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1669390400
transform 1 0 13104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_108
timestamp 1669390400
transform 1 0 13440 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_111
timestamp 1669390400
transform 1 0 13776 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_115
timestamp 1669390400
transform 1 0 14224 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_119
timestamp 1669390400
transform 1 0 14672 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_122
timestamp 1669390400
transform 1 0 15008 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_158
timestamp 1669390400
transform 1 0 19040 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_162
timestamp 1669390400
transform 1 0 19488 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_170
timestamp 1669390400
transform 1 0 20384 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_174
timestamp 1669390400
transform 1 0 20832 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1669390400
transform 1 0 21056 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_179
timestamp 1669390400
transform 1 0 21392 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_187
timestamp 1669390400
transform 1 0 22288 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_195
timestamp 1669390400
transform 1 0 23184 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_199
timestamp 1669390400
transform 1 0 23632 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_207
timestamp 1669390400
transform 1 0 24528 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_211
timestamp 1669390400
transform 1 0 24976 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_214
timestamp 1669390400
transform 1 0 25312 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_220
timestamp 1669390400
transform 1 0 25984 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_230
timestamp 1669390400
transform 1 0 27104 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_239
timestamp 1669390400
transform 1 0 28112 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_247
timestamp 1669390400
transform 1 0 29008 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_250
timestamp 1669390400
transform 1 0 29344 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_256
timestamp 1669390400
transform 1 0 30016 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_283
timestamp 1669390400
transform 1 0 33040 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_289
timestamp 1669390400
transform 1 0 33712 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_293
timestamp 1669390400
transform 1 0 34160 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_297
timestamp 1669390400
transform 1 0 34608 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_306
timestamp 1669390400
transform 1 0 35616 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_314
timestamp 1669390400
transform 1 0 36512 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_318
timestamp 1669390400
transform 1 0 36960 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_321
timestamp 1669390400
transform 1 0 37296 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_330
timestamp 1669390400
transform 1 0 38304 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_340
timestamp 1669390400
transform 1 0 39424 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_344
timestamp 1669390400
transform 1 0 39872 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_347
timestamp 1669390400
transform 1 0 40208 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_357
timestamp 1669390400
transform 1 0 41328 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_365
timestamp 1669390400
transform 1 0 42224 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_367
timestamp 1669390400
transform 1 0 42448 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_380
timestamp 1669390400
transform 1 0 43904 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_388
timestamp 1669390400
transform 1 0 44800 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_392
timestamp 1669390400
transform 1 0 45248 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_395
timestamp 1669390400
transform 1 0 45584 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_399
timestamp 1669390400
transform 1 0 46032 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_406
timestamp 1669390400
transform 1 0 46816 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_410
timestamp 1669390400
transform 1 0 47264 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_418
timestamp 1669390400
transform 1 0 48160 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_421
timestamp 1669390400
transform 1 0 48496 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_435
timestamp 1669390400
transform 1 0 50064 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_443
timestamp 1669390400
transform 1 0 50960 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_451
timestamp 1669390400
transform 1 0 51856 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_459
timestamp 1669390400
transform 1 0 52752 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_463
timestamp 1669390400
transform 1 0 53200 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_486
timestamp 1669390400
transform 1 0 55776 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_490
timestamp 1669390400
transform 1 0 56224 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_504
timestamp 1669390400
transform 1 0 57792 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_512
timestamp 1669390400
transform 1 0 58688 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_2
timestamp 1669390400
transform 1 0 1568 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_18
timestamp 1669390400
transform 1 0 3360 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_26
timestamp 1669390400
transform 1 0 4256 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_38
timestamp 1669390400
transform 1 0 5600 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_54
timestamp 1669390400
transform 1 0 7392 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_62
timestamp 1669390400
transform 1 0 8288 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_66
timestamp 1669390400
transform 1 0 8736 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1669390400
transform 1 0 9184 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_73
timestamp 1669390400
transform 1 0 9520 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_75
timestamp 1669390400
transform 1 0 9744 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_82
timestamp 1669390400
transform 1 0 10528 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_98
timestamp 1669390400
transform 1 0 12320 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_106
timestamp 1669390400
transform 1 0 13216 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1669390400
transform 1 0 17136 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_144
timestamp 1669390400
transform 1 0 17472 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_147
timestamp 1669390400
transform 1 0 17808 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_151
timestamp 1669390400
transform 1 0 18256 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_155
timestamp 1669390400
transform 1 0 18704 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_159
timestamp 1669390400
transform 1 0 19152 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_161
timestamp 1669390400
transform 1 0 19376 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_168
timestamp 1669390400
transform 1 0 20160 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_182
timestamp 1669390400
transform 1 0 21728 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_196
timestamp 1669390400
transform 1 0 23296 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_202
timestamp 1669390400
transform 1 0 23968 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_204
timestamp 1669390400
transform 1 0 24192 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1669390400
transform 1 0 25088 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_215
timestamp 1669390400
transform 1 0 25424 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_223
timestamp 1669390400
transform 1 0 26320 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_231
timestamp 1669390400
transform 1 0 27216 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_235
timestamp 1669390400
transform 1 0 27664 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_239
timestamp 1669390400
transform 1 0 28112 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_243
timestamp 1669390400
transform 1 0 28560 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_247
timestamp 1669390400
transform 1 0 29008 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_251
timestamp 1669390400
transform 1 0 29456 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_255
timestamp 1669390400
transform 1 0 29904 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_259
timestamp 1669390400
transform 1 0 30352 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_263
timestamp 1669390400
transform 1 0 30800 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_275
timestamp 1669390400
transform 1 0 32144 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_282
timestamp 1669390400
transform 1 0 32928 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_286
timestamp 1669390400
transform 1 0 33376 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_289
timestamp 1669390400
transform 1 0 33712 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_297
timestamp 1669390400
transform 1 0 34608 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_311
timestamp 1669390400
transform 1 0 36176 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_315
timestamp 1669390400
transform 1 0 36624 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_319
timestamp 1669390400
transform 1 0 37072 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_321
timestamp 1669390400
transform 1 0 37296 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_330
timestamp 1669390400
transform 1 0 38304 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_340
timestamp 1669390400
transform 1 0 39424 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_344
timestamp 1669390400
transform 1 0 39872 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_348
timestamp 1669390400
transform 1 0 40320 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_352
timestamp 1669390400
transform 1 0 40768 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_354
timestamp 1669390400
transform 1 0 40992 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_357
timestamp 1669390400
transform 1 0 41328 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_360
timestamp 1669390400
transform 1 0 41664 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_364
timestamp 1669390400
transform 1 0 42112 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_367
timestamp 1669390400
transform 1 0 42448 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_371
timestamp 1669390400
transform 1 0 42896 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_375
timestamp 1669390400
transform 1 0 43344 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_385
timestamp 1669390400
transform 1 0 44464 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_389
timestamp 1669390400
transform 1 0 44912 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_393
timestamp 1669390400
transform 1 0 45360 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_397
timestamp 1669390400
transform 1 0 45808 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_399
timestamp 1669390400
transform 1 0 46032 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_413
timestamp 1669390400
transform 1 0 47600 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_421
timestamp 1669390400
transform 1 0 48496 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_425
timestamp 1669390400
transform 1 0 48944 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_428
timestamp 1669390400
transform 1 0 49280 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_435
timestamp 1669390400
transform 1 0 50064 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_437
timestamp 1669390400
transform 1 0 50288 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_450
timestamp 1669390400
transform 1 0 51744 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_458
timestamp 1669390400
transform 1 0 52640 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_472
timestamp 1669390400
transform 1 0 54208 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_482
timestamp 1669390400
transform 1 0 55328 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_489
timestamp 1669390400
transform 1 0 56112 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_499
timestamp 1669390400
transform 1 0 57232 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_507
timestamp 1669390400
transform 1 0 58128 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_511
timestamp 1669390400
transform 1 0 58576 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_2
timestamp 1669390400
transform 1 0 1568 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_18
timestamp 1669390400
transform 1 0 3360 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_26
timestamp 1669390400
transform 1 0 4256 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_30
timestamp 1669390400
transform 1 0 4704 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1669390400
transform 1 0 5152 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_37
timestamp 1669390400
transform 1 0 5488 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_44
timestamp 1669390400
transform 1 0 6272 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_52
timestamp 1669390400
transform 1 0 7168 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_56
timestamp 1669390400
transform 1 0 7616 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_58
timestamp 1669390400
transform 1 0 7840 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_61
timestamp 1669390400
transform 1 0 8176 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_71
timestamp 1669390400
transform 1 0 9296 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_85
timestamp 1669390400
transform 1 0 10864 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_89
timestamp 1669390400
transform 1 0 11312 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_93
timestamp 1669390400
transform 1 0 11760 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1669390400
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1669390400
transform 1 0 13104 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_108
timestamp 1669390400
transform 1 0 13440 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_116
timestamp 1669390400
transform 1 0 14336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_120
timestamp 1669390400
transform 1 0 14784 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_123
timestamp 1669390400
transform 1 0 15120 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_161
timestamp 1669390400
transform 1 0 19376 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_165
timestamp 1669390400
transform 1 0 19824 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_173
timestamp 1669390400
transform 1 0 20720 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_179
timestamp 1669390400
transform 1 0 21392 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_183
timestamp 1669390400
transform 1 0 21840 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_193
timestamp 1669390400
transform 1 0 22960 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_197
timestamp 1669390400
transform 1 0 23408 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_201
timestamp 1669390400
transform 1 0 23856 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_203
timestamp 1669390400
transform 1 0 24080 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_206
timestamp 1669390400
transform 1 0 24416 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_215
timestamp 1669390400
transform 1 0 25424 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_227
timestamp 1669390400
transform 1 0 26768 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_234
timestamp 1669390400
transform 1 0 27552 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_238
timestamp 1669390400
transform 1 0 28000 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_240
timestamp 1669390400
transform 1 0 28224 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_243
timestamp 1669390400
transform 1 0 28560 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_247
timestamp 1669390400
transform 1 0 29008 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_250
timestamp 1669390400
transform 1 0 29344 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_263
timestamp 1669390400
transform 1 0 30800 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_267
timestamp 1669390400
transform 1 0 31248 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_277
timestamp 1669390400
transform 1 0 32368 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_281
timestamp 1669390400
transform 1 0 32816 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_284
timestamp 1669390400
transform 1 0 33152 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_296
timestamp 1669390400
transform 1 0 34496 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_313
timestamp 1669390400
transform 1 0 36400 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_317
timestamp 1669390400
transform 1 0 36848 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_321
timestamp 1669390400
transform 1 0 37296 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_325
timestamp 1669390400
transform 1 0 37744 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_339
timestamp 1669390400
transform 1 0 39312 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_352
timestamp 1669390400
transform 1 0 40768 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_358
timestamp 1669390400
transform 1 0 41440 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_362
timestamp 1669390400
transform 1 0 41888 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_366
timestamp 1669390400
transform 1 0 42336 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_368
timestamp 1669390400
transform 1 0 42560 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_375
timestamp 1669390400
transform 1 0 43344 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_389
timestamp 1669390400
transform 1 0 44912 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_392
timestamp 1669390400
transform 1 0 45248 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_401
timestamp 1669390400
transform 1 0 46256 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_411
timestamp 1669390400
transform 1 0 47376 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_427
timestamp 1669390400
transform 1 0 49168 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_435
timestamp 1669390400
transform 1 0 50064 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_437
timestamp 1669390400
transform 1 0 50288 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_451
timestamp 1669390400
transform 1 0 51856 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_459
timestamp 1669390400
transform 1 0 52752 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_463
timestamp 1669390400
transform 1 0 53200 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_467
timestamp 1669390400
transform 1 0 53648 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_485
timestamp 1669390400
transform 1 0 55664 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_489
timestamp 1669390400
transform 1 0 56112 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_498
timestamp 1669390400
transform 1 0 57120 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_506
timestamp 1669390400
transform 1 0 58016 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_510
timestamp 1669390400
transform 1 0 58464 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_512
timestamp 1669390400
transform 1 0 58688 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_2
timestamp 1669390400
transform 1 0 1568 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_18
timestamp 1669390400
transform 1 0 3360 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_31
timestamp 1669390400
transform 1 0 4816 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_35
timestamp 1669390400
transform 1 0 5264 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_70
timestamp 1669390400
transform 1 0 9184 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_73
timestamp 1669390400
transform 1 0 9520 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_76
timestamp 1669390400
transform 1 0 9856 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_80
timestamp 1669390400
transform 1 0 10304 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_82
timestamp 1669390400
transform 1 0 10528 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_85
timestamp 1669390400
transform 1 0 10864 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_89
timestamp 1669390400
transform 1 0 11312 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1669390400
transform 1 0 17136 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_144
timestamp 1669390400
transform 1 0 17472 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_166
timestamp 1669390400
transform 1 0 19936 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_170
timestamp 1669390400
transform 1 0 20384 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_184
timestamp 1669390400
transform 1 0 21952 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_194
timestamp 1669390400
transform 1 0 23072 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_201
timestamp 1669390400
transform 1 0 23856 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_203
timestamp 1669390400
transform 1 0 24080 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_208
timestamp 1669390400
transform 1 0 24640 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_212
timestamp 1669390400
transform 1 0 25088 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_215
timestamp 1669390400
transform 1 0 25424 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_221
timestamp 1669390400
transform 1 0 26096 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_225
timestamp 1669390400
transform 1 0 26544 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_229
timestamp 1669390400
transform 1 0 26992 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_232
timestamp 1669390400
transform 1 0 27328 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_236
timestamp 1669390400
transform 1 0 27776 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_240
timestamp 1669390400
transform 1 0 28224 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_248
timestamp 1669390400
transform 1 0 29120 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_262
timestamp 1669390400
transform 1 0 30688 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_270
timestamp 1669390400
transform 1 0 31584 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_274
timestamp 1669390400
transform 1 0 32032 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_278
timestamp 1669390400
transform 1 0 32480 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_280
timestamp 1669390400
transform 1 0 32704 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_283
timestamp 1669390400
transform 1 0 33040 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_286
timestamp 1669390400
transform 1 0 33376 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_289
timestamp 1669390400
transform 1 0 33712 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_293
timestamp 1669390400
transform 1 0 34160 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_295
timestamp 1669390400
transform 1 0 34384 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_302
timestamp 1669390400
transform 1 0 35168 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_306
timestamp 1669390400
transform 1 0 35616 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_324
timestamp 1669390400
transform 1 0 37632 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_328
timestamp 1669390400
transform 1 0 38080 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_332
timestamp 1669390400
transform 1 0 38528 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_342
timestamp 1669390400
transform 1 0 39648 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_354
timestamp 1669390400
transform 1 0 40992 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_357
timestamp 1669390400
transform 1 0 41328 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_366
timestamp 1669390400
transform 1 0 42336 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_370
timestamp 1669390400
transform 1 0 42784 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_374
timestamp 1669390400
transform 1 0 43232 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_378
timestamp 1669390400
transform 1 0 43680 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_382
timestamp 1669390400
transform 1 0 44128 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_390
timestamp 1669390400
transform 1 0 45024 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_393
timestamp 1669390400
transform 1 0 45360 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_399
timestamp 1669390400
transform 1 0 46032 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_407
timestamp 1669390400
transform 1 0 46928 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_416
timestamp 1669390400
transform 1 0 47936 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_424
timestamp 1669390400
transform 1 0 48832 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_428
timestamp 1669390400
transform 1 0 49280 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_435
timestamp 1669390400
transform 1 0 50064 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_451
timestamp 1669390400
transform 1 0 51856 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_459
timestamp 1669390400
transform 1 0 52752 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_463
timestamp 1669390400
transform 1 0 53200 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_465
timestamp 1669390400
transform 1 0 53424 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_472
timestamp 1669390400
transform 1 0 54208 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_480
timestamp 1669390400
transform 1 0 55104 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_482
timestamp 1669390400
transform 1 0 55328 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_496
timestamp 1669390400
transform 1 0 56896 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_499
timestamp 1669390400
transform 1 0 57232 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_505
timestamp 1669390400
transform 1 0 57904 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_2
timestamp 1669390400
transform 1 0 1568 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_23
timestamp 1669390400
transform 1 0 3920 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_32
timestamp 1669390400
transform 1 0 4928 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1669390400
transform 1 0 5152 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_37
timestamp 1669390400
transform 1 0 5488 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_72
timestamp 1669390400
transform 1 0 9408 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_74
timestamp 1669390400
transform 1 0 9632 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_83
timestamp 1669390400
transform 1 0 10640 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_87
timestamp 1669390400
transform 1 0 11088 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_91
timestamp 1669390400
transform 1 0 11536 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_93
timestamp 1669390400
transform 1 0 11760 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_96
timestamp 1669390400
transform 1 0 12096 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_100
timestamp 1669390400
transform 1 0 12544 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_102
timestamp 1669390400
transform 1 0 12768 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_105
timestamp 1669390400
transform 1 0 13104 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_108
timestamp 1669390400
transform 1 0 13440 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_111
timestamp 1669390400
transform 1 0 13776 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_113
timestamp 1669390400
transform 1 0 14000 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_116
timestamp 1669390400
transform 1 0 14336 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_120
timestamp 1669390400
transform 1 0 14784 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_124
timestamp 1669390400
transform 1 0 15232 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_159
timestamp 1669390400
transform 1 0 19152 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_175
timestamp 1669390400
transform 1 0 20944 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_179
timestamp 1669390400
transform 1 0 21392 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_203
timestamp 1669390400
transform 1 0 24080 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_207
timestamp 1669390400
transform 1 0 24528 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_211
timestamp 1669390400
transform 1 0 24976 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_217
timestamp 1669390400
transform 1 0 25648 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_227
timestamp 1669390400
transform 1 0 26768 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_235
timestamp 1669390400
transform 1 0 27664 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_239
timestamp 1669390400
transform 1 0 28112 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_243
timestamp 1669390400
transform 1 0 28560 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_247
timestamp 1669390400
transform 1 0 29008 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_250
timestamp 1669390400
transform 1 0 29344 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_259
timestamp 1669390400
transform 1 0 30352 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_269
timestamp 1669390400
transform 1 0 31472 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_273
timestamp 1669390400
transform 1 0 31920 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_277
timestamp 1669390400
transform 1 0 32368 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_281
timestamp 1669390400
transform 1 0 32816 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_283
timestamp 1669390400
transform 1 0 33040 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_297
timestamp 1669390400
transform 1 0 34608 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_301
timestamp 1669390400
transform 1 0 35056 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_317
timestamp 1669390400
transform 1 0 36848 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_321
timestamp 1669390400
transform 1 0 37296 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_329
timestamp 1669390400
transform 1 0 38192 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_333
timestamp 1669390400
transform 1 0 38640 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_337
timestamp 1669390400
transform 1 0 39088 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_343
timestamp 1669390400
transform 1 0 39760 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_353
timestamp 1669390400
transform 1 0 40880 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_360
timestamp 1669390400
transform 1 0 41664 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_364
timestamp 1669390400
transform 1 0 42112 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_368
timestamp 1669390400
transform 1 0 42560 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_381
timestamp 1669390400
transform 1 0 44016 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_389
timestamp 1669390400
transform 1 0 44912 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_392
timestamp 1669390400
transform 1 0 45248 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_394
timestamp 1669390400
transform 1 0 45472 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_397
timestamp 1669390400
transform 1 0 45808 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_423
timestamp 1669390400
transform 1 0 48720 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_425
timestamp 1669390400
transform 1 0 48944 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_438
timestamp 1669390400
transform 1 0 50400 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_448
timestamp 1669390400
transform 1 0 51520 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_460
timestamp 1669390400
transform 1 0 52864 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_463
timestamp 1669390400
transform 1 0 53200 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_479
timestamp 1669390400
transform 1 0 54992 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_487
timestamp 1669390400
transform 1 0 55888 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_494
timestamp 1669390400
transform 1 0 56672 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_510
timestamp 1669390400
transform 1 0 58464 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_512
timestamp 1669390400
transform 1 0 58688 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_2
timestamp 1669390400
transform 1 0 1568 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_18
timestamp 1669390400
transform 1 0 3360 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_32
timestamp 1669390400
transform 1 0 4928 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_68
timestamp 1669390400
transform 1 0 8960 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1669390400
transform 1 0 9184 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_73
timestamp 1669390400
transform 1 0 9520 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_76
timestamp 1669390400
transform 1 0 9856 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_80
timestamp 1669390400
transform 1 0 10304 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_116
timestamp 1669390400
transform 1 0 14336 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_120
timestamp 1669390400
transform 1 0 14784 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_123
timestamp 1669390400
transform 1 0 15120 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_127
timestamp 1669390400
transform 1 0 15568 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_131
timestamp 1669390400
transform 1 0 16016 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_135
timestamp 1669390400
transform 1 0 16464 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_139
timestamp 1669390400
transform 1 0 16912 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_141
timestamp 1669390400
transform 1 0 17136 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_144
timestamp 1669390400
transform 1 0 17472 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_152
timestamp 1669390400
transform 1 0 18368 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_156
timestamp 1669390400
transform 1 0 18816 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_158
timestamp 1669390400
transform 1 0 19040 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_161
timestamp 1669390400
transform 1 0 19376 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_165
timestamp 1669390400
transform 1 0 19824 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_181
timestamp 1669390400
transform 1 0 21616 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_185
timestamp 1669390400
transform 1 0 22064 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_195
timestamp 1669390400
transform 1 0 23184 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_199
timestamp 1669390400
transform 1 0 23632 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_203
timestamp 1669390400
transform 1 0 24080 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1669390400
transform 1 0 25088 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_215
timestamp 1669390400
transform 1 0 25424 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_241
timestamp 1669390400
transform 1 0 28336 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_245
timestamp 1669390400
transform 1 0 28784 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_249
timestamp 1669390400
transform 1 0 29232 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_251
timestamp 1669390400
transform 1 0 29456 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_254
timestamp 1669390400
transform 1 0 29792 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_258
timestamp 1669390400
transform 1 0 30240 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_266
timestamp 1669390400
transform 1 0 31136 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_268
timestamp 1669390400
transform 1 0 31360 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_271
timestamp 1669390400
transform 1 0 31696 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_273
timestamp 1669390400
transform 1 0 31920 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_283
timestamp 1669390400
transform 1 0 33040 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_286
timestamp 1669390400
transform 1 0 33376 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_302
timestamp 1669390400
transform 1 0 35168 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_306
timestamp 1669390400
transform 1 0 35616 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_322
timestamp 1669390400
transform 1 0 37408 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_332
timestamp 1669390400
transform 1 0 38528 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_340
timestamp 1669390400
transform 1 0 39424 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_342
timestamp 1669390400
transform 1 0 39648 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_345
timestamp 1669390400
transform 1 0 39984 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_353
timestamp 1669390400
transform 1 0 40880 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_357
timestamp 1669390400
transform 1 0 41328 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_360
timestamp 1669390400
transform 1 0 41664 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_364
timestamp 1669390400
transform 1 0 42112 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_380
timestamp 1669390400
transform 1 0 43904 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_384
timestamp 1669390400
transform 1 0 44352 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_392
timestamp 1669390400
transform 1 0 45248 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_394
timestamp 1669390400
transform 1 0 45472 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_397
timestamp 1669390400
transform 1 0 45808 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_401
timestamp 1669390400
transform 1 0 46256 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_409
timestamp 1669390400
transform 1 0 47152 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_416
timestamp 1669390400
transform 1 0 47936 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_420
timestamp 1669390400
transform 1 0 48384 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_424
timestamp 1669390400
transform 1 0 48832 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_428
timestamp 1669390400
transform 1 0 49280 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_444
timestamp 1669390400
transform 1 0 51072 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_448
timestamp 1669390400
transform 1 0 51520 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_478
timestamp 1669390400
transform 1 0 54880 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_480
timestamp 1669390400
transform 1 0 55104 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_483
timestamp 1669390400
transform 1 0 55440 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_487
timestamp 1669390400
transform 1 0 55888 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_495
timestamp 1669390400
transform 1 0 56784 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_499
timestamp 1669390400
transform 1 0 57232 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_507
timestamp 1669390400
transform 1 0 58128 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_511
timestamp 1669390400
transform 1 0 58576 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_2
timestamp 1669390400
transform 1 0 1568 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_18
timestamp 1669390400
transform 1 0 3360 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_26
timestamp 1669390400
transform 1 0 4256 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_30
timestamp 1669390400
transform 1 0 4704 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1669390400
transform 1 0 5152 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_37
timestamp 1669390400
transform 1 0 5488 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_40
timestamp 1669390400
transform 1 0 5824 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_44
timestamp 1669390400
transform 1 0 6272 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_47
timestamp 1669390400
transform 1 0 6608 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_51
timestamp 1669390400
transform 1 0 7056 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_55
timestamp 1669390400
transform 1 0 7504 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_59
timestamp 1669390400
transform 1 0 7952 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_63
timestamp 1669390400
transform 1 0 8400 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_65
timestamp 1669390400
transform 1 0 8624 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_68
timestamp 1669390400
transform 1 0 8960 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_70
timestamp 1669390400
transform 1 0 9184 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1669390400
transform 1 0 13104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_108
timestamp 1669390400
transform 1 0 13440 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_111
timestamp 1669390400
transform 1 0 13776 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_115
timestamp 1669390400
transform 1 0 14224 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_119
timestamp 1669390400
transform 1 0 14672 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_123
timestamp 1669390400
transform 1 0 15120 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_159
timestamp 1669390400
transform 1 0 19152 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_163
timestamp 1669390400
transform 1 0 19600 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_171
timestamp 1669390400
transform 1 0 20496 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_175
timestamp 1669390400
transform 1 0 20944 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_179
timestamp 1669390400
transform 1 0 21392 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_186
timestamp 1669390400
transform 1 0 22176 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_188
timestamp 1669390400
transform 1 0 22400 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_195
timestamp 1669390400
transform 1 0 23184 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_199
timestamp 1669390400
transform 1 0 23632 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_202
timestamp 1669390400
transform 1 0 23968 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_206
timestamp 1669390400
transform 1 0 24416 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_214
timestamp 1669390400
transform 1 0 25312 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_218
timestamp 1669390400
transform 1 0 25760 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_221
timestamp 1669390400
transform 1 0 26096 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_231
timestamp 1669390400
transform 1 0 27216 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_238
timestamp 1669390400
transform 1 0 28000 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_240
timestamp 1669390400
transform 1 0 28224 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_243
timestamp 1669390400
transform 1 0 28560 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_247
timestamp 1669390400
transform 1 0 29008 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_250
timestamp 1669390400
transform 1 0 29344 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_262
timestamp 1669390400
transform 1 0 30688 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_266
timestamp 1669390400
transform 1 0 31136 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_270
timestamp 1669390400
transform 1 0 31584 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_274
timestamp 1669390400
transform 1 0 32032 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_276
timestamp 1669390400
transform 1 0 32256 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_286
timestamp 1669390400
transform 1 0 33376 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_298
timestamp 1669390400
transform 1 0 34720 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_306
timestamp 1669390400
transform 1 0 35616 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_310
timestamp 1669390400
transform 1 0 36064 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_314
timestamp 1669390400
transform 1 0 36512 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_318
timestamp 1669390400
transform 1 0 36960 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_321
timestamp 1669390400
transform 1 0 37296 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_345
timestamp 1669390400
transform 1 0 39984 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_361
timestamp 1669390400
transform 1 0 41776 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_365
timestamp 1669390400
transform 1 0 42224 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_375
timestamp 1669390400
transform 1 0 43344 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_389
timestamp 1669390400
transform 1 0 44912 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_392
timestamp 1669390400
transform 1 0 45248 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_400
timestamp 1669390400
transform 1 0 46144 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_413
timestamp 1669390400
transform 1 0 47600 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_417
timestamp 1669390400
transform 1 0 48048 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_421
timestamp 1669390400
transform 1 0 48496 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_425
timestamp 1669390400
transform 1 0 48944 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_440
timestamp 1669390400
transform 1 0 50624 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_456
timestamp 1669390400
transform 1 0 52416 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_460
timestamp 1669390400
transform 1 0 52864 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_463
timestamp 1669390400
transform 1 0 53200 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_465
timestamp 1669390400
transform 1 0 53424 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_478
timestamp 1669390400
transform 1 0 54880 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_482
timestamp 1669390400
transform 1 0 55328 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_495
timestamp 1669390400
transform 1 0 56784 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_497
timestamp 1669390400
transform 1 0 57008 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_500
timestamp 1669390400
transform 1 0 57344 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_508
timestamp 1669390400
transform 1 0 58240 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_512
timestamp 1669390400
transform 1 0 58688 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_2
timestamp 1669390400
transform 1 0 1568 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_18
timestamp 1669390400
transform 1 0 3360 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_70
timestamp 1669390400
transform 1 0 9184 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_73
timestamp 1669390400
transform 1 0 9520 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_76
timestamp 1669390400
transform 1 0 9856 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_80
timestamp 1669390400
transform 1 0 10304 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_83
timestamp 1669390400
transform 1 0 10640 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_87
timestamp 1669390400
transform 1 0 11088 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_89
timestamp 1669390400
transform 1 0 11312 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_140
timestamp 1669390400
transform 1 0 17024 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_144
timestamp 1669390400
transform 1 0 17472 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_147
timestamp 1669390400
transform 1 0 17808 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_151
timestamp 1669390400
transform 1 0 18256 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_155
timestamp 1669390400
transform 1 0 18704 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_159
timestamp 1669390400
transform 1 0 19152 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_162
timestamp 1669390400
transform 1 0 19488 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_166
timestamp 1669390400
transform 1 0 19936 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_170
timestamp 1669390400
transform 1 0 20384 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_183
timestamp 1669390400
transform 1 0 21840 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_197
timestamp 1669390400
transform 1 0 23408 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_203
timestamp 1669390400
transform 1 0 24080 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_205
timestamp 1669390400
transform 1 0 24304 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_208
timestamp 1669390400
transform 1 0 24640 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_212
timestamp 1669390400
transform 1 0 25088 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_215
timestamp 1669390400
transform 1 0 25424 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_219
timestamp 1669390400
transform 1 0 25872 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_223
timestamp 1669390400
transform 1 0 26320 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_227
timestamp 1669390400
transform 1 0 26768 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_231
timestamp 1669390400
transform 1 0 27216 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_235
timestamp 1669390400
transform 1 0 27664 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_239
timestamp 1669390400
transform 1 0 28112 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_243
timestamp 1669390400
transform 1 0 28560 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_247
timestamp 1669390400
transform 1 0 29008 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_251
timestamp 1669390400
transform 1 0 29456 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_255
timestamp 1669390400
transform 1 0 29904 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_266
timestamp 1669390400
transform 1 0 31136 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_273
timestamp 1669390400
transform 1 0 31920 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_277
timestamp 1669390400
transform 1 0 32368 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_281
timestamp 1669390400
transform 1 0 32816 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_283
timestamp 1669390400
transform 1 0 33040 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_286
timestamp 1669390400
transform 1 0 33376 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_289
timestamp 1669390400
transform 1 0 33712 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_293
timestamp 1669390400
transform 1 0 34160 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_297
timestamp 1669390400
transform 1 0 34608 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_303
timestamp 1669390400
transform 1 0 35280 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_305
timestamp 1669390400
transform 1 0 35504 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_314
timestamp 1669390400
transform 1 0 36512 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_324
timestamp 1669390400
transform 1 0 37632 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_332
timestamp 1669390400
transform 1 0 38528 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_336
timestamp 1669390400
transform 1 0 38976 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_340
timestamp 1669390400
transform 1 0 39424 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_354
timestamp 1669390400
transform 1 0 40992 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_357
timestamp 1669390400
transform 1 0 41328 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_363
timestamp 1669390400
transform 1 0 42000 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_373
timestamp 1669390400
transform 1 0 43120 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_383
timestamp 1669390400
transform 1 0 44240 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_387
timestamp 1669390400
transform 1 0 44688 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_389
timestamp 1669390400
transform 1 0 44912 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_392
timestamp 1669390400
transform 1 0 45248 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_402
timestamp 1669390400
transform 1 0 46368 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_412
timestamp 1669390400
transform 1 0 47488 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_416
timestamp 1669390400
transform 1 0 47936 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_418
timestamp 1669390400
transform 1 0 48160 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_425
timestamp 1669390400
transform 1 0 48944 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_428
timestamp 1669390400
transform 1 0 49280 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_437
timestamp 1669390400
transform 1 0 50288 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_453
timestamp 1669390400
transform 1 0 52080 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_469
timestamp 1669390400
transform 1 0 53872 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_479
timestamp 1669390400
transform 1 0 54992 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_496
timestamp 1669390400
transform 1 0 56896 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_499
timestamp 1669390400
transform 1 0 57232 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_512
timestamp 1669390400
transform 1 0 58688 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_2
timestamp 1669390400
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_34
timestamp 1669390400
transform 1 0 5152 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_37
timestamp 1669390400
transform 1 0 5488 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_39
timestamp 1669390400
transform 1 0 5712 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_42
timestamp 1669390400
transform 1 0 6048 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_46
timestamp 1669390400
transform 1 0 6496 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_50
timestamp 1669390400
transform 1 0 6944 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_54
timestamp 1669390400
transform 1 0 7392 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_58
timestamp 1669390400
transform 1 0 7840 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_94
timestamp 1669390400
transform 1 0 11872 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_98
timestamp 1669390400
transform 1 0 12320 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_101
timestamp 1669390400
transform 1 0 12656 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1669390400
transform 1 0 13104 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_108
timestamp 1669390400
transform 1 0 13440 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_111
timestamp 1669390400
transform 1 0 13776 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_115
timestamp 1669390400
transform 1 0 14224 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_119
timestamp 1669390400
transform 1 0 14672 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_123
timestamp 1669390400
transform 1 0 15120 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_159
timestamp 1669390400
transform 1 0 19152 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_163
timestamp 1669390400
transform 1 0 19600 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_167
timestamp 1669390400
transform 1 0 20048 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_169
timestamp 1669390400
transform 1 0 20272 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_172
timestamp 1669390400
transform 1 0 20608 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_176
timestamp 1669390400
transform 1 0 21056 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_179
timestamp 1669390400
transform 1 0 21392 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_183
timestamp 1669390400
transform 1 0 21840 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_193
timestamp 1669390400
transform 1 0 22960 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_197
timestamp 1669390400
transform 1 0 23408 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_201
timestamp 1669390400
transform 1 0 23856 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_207
timestamp 1669390400
transform 1 0 24528 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_211
timestamp 1669390400
transform 1 0 24976 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_225
timestamp 1669390400
transform 1 0 26544 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_229
timestamp 1669390400
transform 1 0 26992 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_236
timestamp 1669390400
transform 1 0 27776 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_238
timestamp 1669390400
transform 1 0 28000 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_241
timestamp 1669390400
transform 1 0 28336 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_245
timestamp 1669390400
transform 1 0 28784 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_247
timestamp 1669390400
transform 1 0 29008 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_250
timestamp 1669390400
transform 1 0 29344 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_255
timestamp 1669390400
transform 1 0 29904 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_263
timestamp 1669390400
transform 1 0 30800 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_270
timestamp 1669390400
transform 1 0 31584 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_274
timestamp 1669390400
transform 1 0 32032 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_278
timestamp 1669390400
transform 1 0 32480 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_282
timestamp 1669390400
transform 1 0 32928 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_286
timestamp 1669390400
transform 1 0 33376 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_290
timestamp 1669390400
transform 1 0 33824 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_296
timestamp 1669390400
transform 1 0 34496 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_300
timestamp 1669390400
transform 1 0 34944 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_302
timestamp 1669390400
transform 1 0 35168 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_311
timestamp 1669390400
transform 1 0 36176 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_315
timestamp 1669390400
transform 1 0 36624 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_321
timestamp 1669390400
transform 1 0 37296 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_324
timestamp 1669390400
transform 1 0 37632 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_328
timestamp 1669390400
transform 1 0 38080 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_330
timestamp 1669390400
transform 1 0 38304 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_333
timestamp 1669390400
transform 1 0 38640 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_340
timestamp 1669390400
transform 1 0 39424 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_354
timestamp 1669390400
transform 1 0 40992 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_358
timestamp 1669390400
transform 1 0 41440 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_362
timestamp 1669390400
transform 1 0 41888 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_366
timestamp 1669390400
transform 1 0 42336 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_373
timestamp 1669390400
transform 1 0 43120 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_383
timestamp 1669390400
transform 1 0 44240 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_387
timestamp 1669390400
transform 1 0 44688 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_389
timestamp 1669390400
transform 1 0 44912 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_392
timestamp 1669390400
transform 1 0 45248 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_394
timestamp 1669390400
transform 1 0 45472 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_401
timestamp 1669390400
transform 1 0 46256 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_407
timestamp 1669390400
transform 1 0 46928 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_423
timestamp 1669390400
transform 1 0 48720 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_429
timestamp 1669390400
transform 1 0 49392 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_445
timestamp 1669390400
transform 1 0 51184 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_453
timestamp 1669390400
transform 1 0 52080 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_460
timestamp 1669390400
transform 1 0 52864 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_463
timestamp 1669390400
transform 1 0 53200 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_470
timestamp 1669390400
transform 1 0 53984 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_512
timestamp 1669390400
transform 1 0 58688 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_2
timestamp 1669390400
transform 1 0 1568 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_18
timestamp 1669390400
transform 1 0 3360 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_26
timestamp 1669390400
transform 1 0 4256 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_30
timestamp 1669390400
transform 1 0 4704 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_34
timestamp 1669390400
transform 1 0 5152 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_70
timestamp 1669390400
transform 1 0 9184 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_73
timestamp 1669390400
transform 1 0 9520 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_76
timestamp 1669390400
transform 1 0 9856 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_80
timestamp 1669390400
transform 1 0 10304 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_84
timestamp 1669390400
transform 1 0 10752 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_86
timestamp 1669390400
transform 1 0 10976 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_123
timestamp 1669390400
transform 1 0 15120 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_129
timestamp 1669390400
transform 1 0 15792 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_133
timestamp 1669390400
transform 1 0 16240 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_137
timestamp 1669390400
transform 1 0 16688 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_141
timestamp 1669390400
transform 1 0 17136 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_144
timestamp 1669390400
transform 1 0 17472 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_147
timestamp 1669390400
transform 1 0 17808 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_151
timestamp 1669390400
transform 1 0 18256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_157
timestamp 1669390400
transform 1 0 18928 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_161
timestamp 1669390400
transform 1 0 19376 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_163
timestamp 1669390400
transform 1 0 19600 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_166
timestamp 1669390400
transform 1 0 19936 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_172
timestamp 1669390400
transform 1 0 20608 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_176
timestamp 1669390400
transform 1 0 21056 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_180
timestamp 1669390400
transform 1 0 21504 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_188
timestamp 1669390400
transform 1 0 22400 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_192
timestamp 1669390400
transform 1 0 22848 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_195
timestamp 1669390400
transform 1 0 23184 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_199
timestamp 1669390400
transform 1 0 23632 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_203
timestamp 1669390400
transform 1 0 24080 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_205
timestamp 1669390400
transform 1 0 24304 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_208
timestamp 1669390400
transform 1 0 24640 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_212
timestamp 1669390400
transform 1 0 25088 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_215
timestamp 1669390400
transform 1 0 25424 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_219
timestamp 1669390400
transform 1 0 25872 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_223
timestamp 1669390400
transform 1 0 26320 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_237
timestamp 1669390400
transform 1 0 27888 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_247
timestamp 1669390400
transform 1 0 29008 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_249
timestamp 1669390400
transform 1 0 29232 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_252
timestamp 1669390400
transform 1 0 29568 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_262
timestamp 1669390400
transform 1 0 30688 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_266
timestamp 1669390400
transform 1 0 31136 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_270
timestamp 1669390400
transform 1 0 31584 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_274
timestamp 1669390400
transform 1 0 32032 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_283
timestamp 1669390400
transform 1 0 33040 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_286
timestamp 1669390400
transform 1 0 33376 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_296
timestamp 1669390400
transform 1 0 34496 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_300
timestamp 1669390400
transform 1 0 34944 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_312
timestamp 1669390400
transform 1 0 36288 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_316
timestamp 1669390400
transform 1 0 36736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_332
timestamp 1669390400
transform 1 0 38528 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_336
timestamp 1669390400
transform 1 0 38976 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_340
timestamp 1669390400
transform 1 0 39424 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_343
timestamp 1669390400
transform 1 0 39760 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_352
timestamp 1669390400
transform 1 0 40768 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_354
timestamp 1669390400
transform 1 0 40992 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_357
timestamp 1669390400
transform 1 0 41328 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_360
timestamp 1669390400
transform 1 0 41664 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_364
timestamp 1669390400
transform 1 0 42112 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_377
timestamp 1669390400
transform 1 0 43568 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_381
timestamp 1669390400
transform 1 0 44016 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_385
timestamp 1669390400
transform 1 0 44464 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_389
timestamp 1669390400
transform 1 0 44912 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_393
timestamp 1669390400
transform 1 0 45360 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_397
timestamp 1669390400
transform 1 0 45808 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_413
timestamp 1669390400
transform 1 0 47600 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_421
timestamp 1669390400
transform 1 0 48496 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_425
timestamp 1669390400
transform 1 0 48944 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_428
timestamp 1669390400
transform 1 0 49280 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_430
timestamp 1669390400
transform 1 0 49504 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_443
timestamp 1669390400
transform 1 0 50960 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_447
timestamp 1669390400
transform 1 0 51408 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_449
timestamp 1669390400
transform 1 0 51632 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_462
timestamp 1669390400
transform 1 0 53088 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_472
timestamp 1669390400
transform 1 0 54208 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_476
timestamp 1669390400
transform 1 0 54656 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_496
timestamp 1669390400
transform 1 0 56896 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_499
timestamp 1669390400
transform 1 0 57232 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_512
timestamp 1669390400
transform 1 0 58688 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_2
timestamp 1669390400
transform 1 0 1568 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_18
timestamp 1669390400
transform 1 0 3360 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_22
timestamp 1669390400
transform 1 0 3808 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_26
timestamp 1669390400
transform 1 0 4256 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_30
timestamp 1669390400
transform 1 0 4704 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_34
timestamp 1669390400
transform 1 0 5152 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_37
timestamp 1669390400
transform 1 0 5488 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_40
timestamp 1669390400
transform 1 0 5824 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_44
timestamp 1669390400
transform 1 0 6272 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_48
timestamp 1669390400
transform 1 0 6720 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_52
timestamp 1669390400
transform 1 0 7168 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_56
timestamp 1669390400
transform 1 0 7616 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_60
timestamp 1669390400
transform 1 0 8064 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_62
timestamp 1669390400
transform 1 0 8288 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_65
timestamp 1669390400
transform 1 0 8624 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_69
timestamp 1669390400
transform 1 0 9072 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_105
timestamp 1669390400
transform 1 0 13104 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_108
timestamp 1669390400
transform 1 0 13440 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_111
timestamp 1669390400
transform 1 0 13776 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_113
timestamp 1669390400
transform 1 0 14000 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_116
timestamp 1669390400
transform 1 0 14336 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_120
timestamp 1669390400
transform 1 0 14784 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_124
timestamp 1669390400
transform 1 0 15232 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_160
timestamp 1669390400
transform 1 0 19264 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_164
timestamp 1669390400
transform 1 0 19712 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_168
timestamp 1669390400
transform 1 0 20160 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_172
timestamp 1669390400
transform 1 0 20608 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_176
timestamp 1669390400
transform 1 0 21056 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_179
timestamp 1669390400
transform 1 0 21392 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_181
timestamp 1669390400
transform 1 0 21616 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_190
timestamp 1669390400
transform 1 0 22624 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_196
timestamp 1669390400
transform 1 0 23296 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_202
timestamp 1669390400
transform 1 0 23968 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_204
timestamp 1669390400
transform 1 0 24192 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_207
timestamp 1669390400
transform 1 0 24528 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_211
timestamp 1669390400
transform 1 0 24976 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_221
timestamp 1669390400
transform 1 0 26096 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_231
timestamp 1669390400
transform 1 0 27216 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_235
timestamp 1669390400
transform 1 0 27664 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_237
timestamp 1669390400
transform 1 0 27888 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_240
timestamp 1669390400
transform 1 0 28224 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_246
timestamp 1669390400
transform 1 0 28896 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_250
timestamp 1669390400
transform 1 0 29344 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_269
timestamp 1669390400
transform 1 0 31472 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_273
timestamp 1669390400
transform 1 0 31920 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_289
timestamp 1669390400
transform 1 0 33712 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_303
timestamp 1669390400
transform 1 0 35280 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_314
timestamp 1669390400
transform 1 0 36512 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_318
timestamp 1669390400
transform 1 0 36960 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_321
timestamp 1669390400
transform 1 0 37296 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_329
timestamp 1669390400
transform 1 0 38192 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_344
timestamp 1669390400
transform 1 0 39872 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_351
timestamp 1669390400
transform 1 0 40656 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_355
timestamp 1669390400
transform 1 0 41104 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_359
timestamp 1669390400
transform 1 0 41552 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_373
timestamp 1669390400
transform 1 0 43120 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_388
timestamp 1669390400
transform 1 0 44800 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_392
timestamp 1669390400
transform 1 0 45248 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_413
timestamp 1669390400
transform 1 0 47600 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_421
timestamp 1669390400
transform 1 0 48496 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_428
timestamp 1669390400
transform 1 0 49280 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_432
timestamp 1669390400
transform 1 0 49728 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_437
timestamp 1669390400
transform 1 0 50288 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_454
timestamp 1669390400
transform 1 0 52192 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_458
timestamp 1669390400
transform 1 0 52640 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_460
timestamp 1669390400
transform 1 0 52864 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_463
timestamp 1669390400
transform 1 0 53200 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_466
timestamp 1669390400
transform 1 0 53536 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_470
timestamp 1669390400
transform 1 0 53984 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_478
timestamp 1669390400
transform 1 0 54880 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_512
timestamp 1669390400
transform 1 0 58688 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_2
timestamp 1669390400
transform 1 0 1568 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_10
timestamp 1669390400
transform 1 0 2464 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_14
timestamp 1669390400
transform 1 0 2912 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_16
timestamp 1669390400
transform 1 0 3136 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_19
timestamp 1669390400
transform 1 0 3472 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_23
timestamp 1669390400
transform 1 0 3920 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_27
timestamp 1669390400
transform 1 0 4368 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_31
timestamp 1669390400
transform 1 0 4816 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_67
timestamp 1669390400
transform 1 0 8848 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_73
timestamp 1669390400
transform 1 0 9520 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_79
timestamp 1669390400
transform 1 0 10192 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_83
timestamp 1669390400
transform 1 0 10640 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_87
timestamp 1669390400
transform 1 0 11088 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_90
timestamp 1669390400
transform 1 0 11424 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_94
timestamp 1669390400
transform 1 0 11872 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_98
timestamp 1669390400
transform 1 0 12320 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_102
timestamp 1669390400
transform 1 0 12768 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_106
timestamp 1669390400
transform 1 0 13216 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_141
timestamp 1669390400
transform 1 0 17136 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_144
timestamp 1669390400
transform 1 0 17472 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_146
timestamp 1669390400
transform 1 0 17696 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_149
timestamp 1669390400
transform 1 0 18032 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_153
timestamp 1669390400
transform 1 0 18480 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_157
timestamp 1669390400
transform 1 0 18928 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_161
timestamp 1669390400
transform 1 0 19376 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_165
timestamp 1669390400
transform 1 0 19824 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_169
timestamp 1669390400
transform 1 0 20272 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_171
timestamp 1669390400
transform 1 0 20496 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_195
timestamp 1669390400
transform 1 0 23184 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_203
timestamp 1669390400
transform 1 0 24080 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_205
timestamp 1669390400
transform 1 0 24304 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_212
timestamp 1669390400
transform 1 0 25088 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_215
timestamp 1669390400
transform 1 0 25424 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_224
timestamp 1669390400
transform 1 0 26432 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_232
timestamp 1669390400
transform 1 0 27328 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_239
timestamp 1669390400
transform 1 0 28112 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_243
timestamp 1669390400
transform 1 0 28560 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_247
timestamp 1669390400
transform 1 0 29008 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_249
timestamp 1669390400
transform 1 0 29232 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_262
timestamp 1669390400
transform 1 0 30688 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_266
timestamp 1669390400
transform 1 0 31136 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_268
timestamp 1669390400
transform 1 0 31360 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_271
timestamp 1669390400
transform 1 0 31696 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_282
timestamp 1669390400
transform 1 0 32928 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_286
timestamp 1669390400
transform 1 0 33376 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_289
timestamp 1669390400
transform 1 0 33712 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_291
timestamp 1669390400
transform 1 0 33936 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_300
timestamp 1669390400
transform 1 0 34944 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_304
timestamp 1669390400
transform 1 0 35392 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_308
timestamp 1669390400
transform 1 0 35840 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_312
timestamp 1669390400
transform 1 0 36288 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_316
timestamp 1669390400
transform 1 0 36736 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_320
timestamp 1669390400
transform 1 0 37184 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_324
timestamp 1669390400
transform 1 0 37632 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_328
timestamp 1669390400
transform 1 0 38080 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_330
timestamp 1669390400
transform 1 0 38304 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_339
timestamp 1669390400
transform 1 0 39312 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_349
timestamp 1669390400
transform 1 0 40432 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_351
timestamp 1669390400
transform 1 0 40656 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_354
timestamp 1669390400
transform 1 0 40992 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_357
timestamp 1669390400
transform 1 0 41328 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_368
timestamp 1669390400
transform 1 0 42560 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_372
timestamp 1669390400
transform 1 0 43008 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_374
timestamp 1669390400
transform 1 0 43232 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_383
timestamp 1669390400
transform 1 0 44240 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_387
timestamp 1669390400
transform 1 0 44688 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_391
timestamp 1669390400
transform 1 0 45136 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_405
timestamp 1669390400
transform 1 0 46704 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_425
timestamp 1669390400
transform 1 0 48944 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_428
timestamp 1669390400
transform 1 0 49280 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_442
timestamp 1669390400
transform 1 0 50848 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_461
timestamp 1669390400
transform 1 0 52976 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_492
timestamp 1669390400
transform 1 0 56448 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_496
timestamp 1669390400
transform 1 0 56896 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_499
timestamp 1669390400
transform 1 0 57232 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_510
timestamp 1669390400
transform 1 0 58464 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_512
timestamp 1669390400
transform 1 0 58688 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_2
timestamp 1669390400
transform 1 0 1568 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_6
timestamp 1669390400
transform 1 0 2016 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_10
timestamp 1669390400
transform 1 0 2464 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_14
timestamp 1669390400
transform 1 0 2912 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_18
timestamp 1669390400
transform 1 0 3360 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_22
timestamp 1669390400
transform 1 0 3808 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_26
timestamp 1669390400
transform 1 0 4256 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_30
timestamp 1669390400
transform 1 0 4704 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_34
timestamp 1669390400
transform 1 0 5152 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_37
timestamp 1669390400
transform 1 0 5488 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_41
timestamp 1669390400
transform 1 0 5936 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_45
timestamp 1669390400
transform 1 0 6384 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_49
timestamp 1669390400
transform 1 0 6832 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_53
timestamp 1669390400
transform 1 0 7280 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_57
timestamp 1669390400
transform 1 0 7728 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_61
timestamp 1669390400
transform 1 0 8176 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_65
timestamp 1669390400
transform 1 0 8624 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_69
timestamp 1669390400
transform 1 0 9072 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_71
timestamp 1669390400
transform 1 0 9296 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_78
timestamp 1669390400
transform 1 0 10080 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_80
timestamp 1669390400
transform 1 0 10304 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_83
timestamp 1669390400
transform 1 0 10640 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_87
timestamp 1669390400
transform 1 0 11088 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_91
timestamp 1669390400
transform 1 0 11536 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_97
timestamp 1669390400
transform 1 0 12208 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_101
timestamp 1669390400
transform 1 0 12656 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_105
timestamp 1669390400
transform 1 0 13104 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_108
timestamp 1669390400
transform 1 0 13440 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_111
timestamp 1669390400
transform 1 0 13776 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_117
timestamp 1669390400
transform 1 0 14448 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_121
timestamp 1669390400
transform 1 0 14896 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_159
timestamp 1669390400
transform 1 0 19152 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_163
timestamp 1669390400
transform 1 0 19600 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_165
timestamp 1669390400
transform 1 0 19824 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_168
timestamp 1669390400
transform 1 0 20160 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_172
timestamp 1669390400
transform 1 0 20608 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_176
timestamp 1669390400
transform 1 0 21056 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_179
timestamp 1669390400
transform 1 0 21392 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_189
timestamp 1669390400
transform 1 0 22512 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_196
timestamp 1669390400
transform 1 0 23296 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_202
timestamp 1669390400
transform 1 0 23968 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_227
timestamp 1669390400
transform 1 0 26768 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_231
timestamp 1669390400
transform 1 0 27216 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_235
timestamp 1669390400
transform 1 0 27664 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_239
timestamp 1669390400
transform 1 0 28112 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_243
timestamp 1669390400
transform 1 0 28560 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_247
timestamp 1669390400
transform 1 0 29008 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_250
timestamp 1669390400
transform 1 0 29344 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_253
timestamp 1669390400
transform 1 0 29680 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_257
timestamp 1669390400
transform 1 0 30128 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_260
timestamp 1669390400
transform 1 0 30464 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_264
timestamp 1669390400
transform 1 0 30912 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_268
timestamp 1669390400
transform 1 0 31360 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_272
timestamp 1669390400
transform 1 0 31808 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_276
timestamp 1669390400
transform 1 0 32256 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_280
timestamp 1669390400
transform 1 0 32704 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_284
timestamp 1669390400
transform 1 0 33152 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_288
timestamp 1669390400
transform 1 0 33600 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_292
timestamp 1669390400
transform 1 0 34048 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_296
timestamp 1669390400
transform 1 0 34496 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_300
timestamp 1669390400
transform 1 0 34944 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_304
timestamp 1669390400
transform 1 0 35392 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_317
timestamp 1669390400
transform 1 0 36848 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_321
timestamp 1669390400
transform 1 0 37296 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_324
timestamp 1669390400
transform 1 0 37632 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_328
timestamp 1669390400
transform 1 0 38080 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_332
timestamp 1669390400
transform 1 0 38528 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_336
timestamp 1669390400
transform 1 0 38976 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_338
timestamp 1669390400
transform 1 0 39200 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_341
timestamp 1669390400
transform 1 0 39536 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_345
timestamp 1669390400
transform 1 0 39984 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_348
timestamp 1669390400
transform 1 0 40320 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_352
timestamp 1669390400
transform 1 0 40768 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_355
timestamp 1669390400
transform 1 0 41104 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_362
timestamp 1669390400
transform 1 0 41888 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_364
timestamp 1669390400
transform 1 0 42112 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_378
timestamp 1669390400
transform 1 0 43680 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_385
timestamp 1669390400
transform 1 0 44464 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_389
timestamp 1669390400
transform 1 0 44912 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_392
timestamp 1669390400
transform 1 0 45248 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_404
timestamp 1669390400
transform 1 0 46592 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_414
timestamp 1669390400
transform 1 0 47712 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_422
timestamp 1669390400
transform 1 0 48608 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_424
timestamp 1669390400
transform 1 0 48832 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_430
timestamp 1669390400
transform 1 0 49504 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_432
timestamp 1669390400
transform 1 0 49728 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_441
timestamp 1669390400
transform 1 0 50736 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_450
timestamp 1669390400
transform 1 0 51744 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_460
timestamp 1669390400
transform 1 0 52864 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_463
timestamp 1669390400
transform 1 0 53200 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_465
timestamp 1669390400
transform 1 0 53424 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_474
timestamp 1669390400
transform 1 0 54432 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_512
timestamp 1669390400
transform 1 0 58688 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_2
timestamp 1669390400
transform 1 0 1568 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_5
timestamp 1669390400
transform 1 0 1904 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_9
timestamp 1669390400
transform 1 0 2352 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_13
timestamp 1669390400
transform 1 0 2800 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_17
timestamp 1669390400
transform 1 0 3248 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_21
timestamp 1669390400
transform 1 0 3696 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_25
timestamp 1669390400
transform 1 0 4144 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_29
timestamp 1669390400
transform 1 0 4592 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_37
timestamp 1669390400
transform 1 0 5488 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_45
timestamp 1669390400
transform 1 0 6384 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_47
timestamp 1669390400
transform 1 0 6608 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_59
timestamp 1669390400
transform 1 0 7952 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_63
timestamp 1669390400
transform 1 0 8400 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_67
timestamp 1669390400
transform 1 0 8848 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_70
timestamp 1669390400
transform 1 0 9184 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_73
timestamp 1669390400
transform 1 0 9520 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_75
timestamp 1669390400
transform 1 0 9744 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_88
timestamp 1669390400
transform 1 0 11200 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_90
timestamp 1669390400
transform 1 0 11424 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_97
timestamp 1669390400
transform 1 0 12208 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_111
timestamp 1669390400
transform 1 0 13776 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_115
timestamp 1669390400
transform 1 0 14224 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_118
timestamp 1669390400
transform 1 0 14560 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_122
timestamp 1669390400
transform 1 0 15008 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_125
timestamp 1669390400
transform 1 0 15344 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_129
timestamp 1669390400
transform 1 0 15792 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_133
timestamp 1669390400
transform 1 0 16240 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_137
timestamp 1669390400
transform 1 0 16688 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_141
timestamp 1669390400
transform 1 0 17136 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_144
timestamp 1669390400
transform 1 0 17472 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_146
timestamp 1669390400
transform 1 0 17696 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_149
timestamp 1669390400
transform 1 0 18032 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_153
timestamp 1669390400
transform 1 0 18480 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_157
timestamp 1669390400
transform 1 0 18928 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_161
timestamp 1669390400
transform 1 0 19376 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_173
timestamp 1669390400
transform 1 0 20720 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_182
timestamp 1669390400
transform 1 0 21728 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_188
timestamp 1669390400
transform 1 0 22400 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_192
timestamp 1669390400
transform 1 0 22848 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_195
timestamp 1669390400
transform 1 0 23184 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_202
timestamp 1669390400
transform 1 0 23968 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_208
timestamp 1669390400
transform 1 0 24640 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_212
timestamp 1669390400
transform 1 0 25088 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_215
timestamp 1669390400
transform 1 0 25424 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_222
timestamp 1669390400
transform 1 0 26208 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_226
timestamp 1669390400
transform 1 0 26656 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_230
timestamp 1669390400
transform 1 0 27104 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_233
timestamp 1669390400
transform 1 0 27440 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_241
timestamp 1669390400
transform 1 0 28336 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_251
timestamp 1669390400
transform 1 0 29456 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_266
timestamp 1669390400
transform 1 0 31136 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_275
timestamp 1669390400
transform 1 0 32144 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_283
timestamp 1669390400
transform 1 0 33040 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_286
timestamp 1669390400
transform 1 0 33376 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_306
timestamp 1669390400
transform 1 0 35616 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_310
timestamp 1669390400
transform 1 0 36064 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_317
timestamp 1669390400
transform 1 0 36848 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_342
timestamp 1669390400
transform 1 0 39648 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_346
timestamp 1669390400
transform 1 0 40096 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_350
timestamp 1669390400
transform 1 0 40544 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_354
timestamp 1669390400
transform 1 0 40992 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_357
timestamp 1669390400
transform 1 0 41328 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_373
timestamp 1669390400
transform 1 0 43120 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_389
timestamp 1669390400
transform 1 0 44912 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_397
timestamp 1669390400
transform 1 0 45808 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_400
timestamp 1669390400
transform 1 0 46144 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_408
timestamp 1669390400
transform 1 0 47040 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_412
timestamp 1669390400
transform 1 0 47488 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_416
timestamp 1669390400
transform 1 0 47936 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_420
timestamp 1669390400
transform 1 0 48384 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_424
timestamp 1669390400
transform 1 0 48832 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_428
timestamp 1669390400
transform 1 0 49280 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_444
timestamp 1669390400
transform 1 0 51072 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_452
timestamp 1669390400
transform 1 0 51968 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_456
timestamp 1669390400
transform 1 0 52416 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_481
timestamp 1669390400
transform 1 0 55216 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_485
timestamp 1669390400
transform 1 0 55664 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_496
timestamp 1669390400
transform 1 0 56896 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_499
timestamp 1669390400
transform 1 0 57232 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_510
timestamp 1669390400
transform 1 0 58464 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_512
timestamp 1669390400
transform 1 0 58688 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_2
timestamp 1669390400
transform 1 0 1568 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_6
timestamp 1669390400
transform 1 0 2016 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_10
timestamp 1669390400
transform 1 0 2464 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_14
timestamp 1669390400
transform 1 0 2912 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_18
timestamp 1669390400
transform 1 0 3360 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_22
timestamp 1669390400
transform 1 0 3808 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_26
timestamp 1669390400
transform 1 0 4256 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_30
timestamp 1669390400
transform 1 0 4704 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_34
timestamp 1669390400
transform 1 0 5152 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_37
timestamp 1669390400
transform 1 0 5488 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_40
timestamp 1669390400
transform 1 0 5824 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_44
timestamp 1669390400
transform 1 0 6272 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_58
timestamp 1669390400
transform 1 0 7840 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_62
timestamp 1669390400
transform 1 0 8288 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_65
timestamp 1669390400
transform 1 0 8624 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_80
timestamp 1669390400
transform 1 0 10304 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_95
timestamp 1669390400
transform 1 0 11984 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_99
timestamp 1669390400
transform 1 0 12432 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_105
timestamp 1669390400
transform 1 0 13104 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_108
timestamp 1669390400
transform 1 0 13440 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_115
timestamp 1669390400
transform 1 0 14224 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_125
timestamp 1669390400
transform 1 0 15344 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_127
timestamp 1669390400
transform 1 0 15568 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_130
timestamp 1669390400
transform 1 0 15904 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_138
timestamp 1669390400
transform 1 0 16800 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_140
timestamp 1669390400
transform 1 0 17024 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_143
timestamp 1669390400
transform 1 0 17360 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_147
timestamp 1669390400
transform 1 0 17808 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_151
timestamp 1669390400
transform 1 0 18256 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_155
timestamp 1669390400
transform 1 0 18704 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_159
timestamp 1669390400
transform 1 0 19152 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_175
timestamp 1669390400
transform 1 0 20944 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_179
timestamp 1669390400
transform 1 0 21392 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_192
timestamp 1669390400
transform 1 0 22848 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_199
timestamp 1669390400
transform 1 0 23632 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_207
timestamp 1669390400
transform 1 0 24528 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_213
timestamp 1669390400
transform 1 0 25200 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_217
timestamp 1669390400
transform 1 0 25648 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_221
timestamp 1669390400
transform 1 0 26096 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_234
timestamp 1669390400
transform 1 0 27552 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_247
timestamp 1669390400
transform 1 0 29008 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_250
timestamp 1669390400
transform 1 0 29344 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_267
timestamp 1669390400
transform 1 0 31248 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_275
timestamp 1669390400
transform 1 0 32144 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_300
timestamp 1669390400
transform 1 0 34944 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_313
timestamp 1669390400
transform 1 0 36400 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_317
timestamp 1669390400
transform 1 0 36848 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_321
timestamp 1669390400
transform 1 0 37296 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_330
timestamp 1669390400
transform 1 0 38304 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_334
timestamp 1669390400
transform 1 0 38752 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_338
timestamp 1669390400
transform 1 0 39200 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_342
timestamp 1669390400
transform 1 0 39648 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_346
timestamp 1669390400
transform 1 0 40096 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_357
timestamp 1669390400
transform 1 0 41328 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_361
timestamp 1669390400
transform 1 0 41776 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_370
timestamp 1669390400
transform 1 0 42784 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_374
timestamp 1669390400
transform 1 0 43232 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_392
timestamp 1669390400
transform 1 0 45248 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_398
timestamp 1669390400
transform 1 0 45920 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_424
timestamp 1669390400
transform 1 0 48832 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_426
timestamp 1669390400
transform 1 0 49056 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_429
timestamp 1669390400
transform 1 0 49392 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_433
timestamp 1669390400
transform 1 0 49840 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_435
timestamp 1669390400
transform 1 0 50064 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_448
timestamp 1669390400
transform 1 0 51520 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_456
timestamp 1669390400
transform 1 0 52416 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_460
timestamp 1669390400
transform 1 0 52864 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_463
timestamp 1669390400
transform 1 0 53200 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_467
timestamp 1669390400
transform 1 0 53648 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_470
timestamp 1669390400
transform 1 0 53984 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_477
timestamp 1669390400
transform 1 0 54768 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_512
timestamp 1669390400
transform 1 0 58688 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_2
timestamp 1669390400
transform 1 0 1568 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_5
timestamp 1669390400
transform 1 0 1904 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_9
timestamp 1669390400
transform 1 0 2352 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_13
timestamp 1669390400
transform 1 0 2800 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_17
timestamp 1669390400
transform 1 0 3248 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_21
timestamp 1669390400
transform 1 0 3696 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_25
timestamp 1669390400
transform 1 0 4144 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_29
timestamp 1669390400
transform 1 0 4592 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_33
timestamp 1669390400
transform 1 0 5040 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_37
timestamp 1669390400
transform 1 0 5488 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_45
timestamp 1669390400
transform 1 0 6384 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_49
timestamp 1669390400
transform 1 0 6832 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_55
timestamp 1669390400
transform 1 0 7504 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_66
timestamp 1669390400
transform 1 0 8736 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_70
timestamp 1669390400
transform 1 0 9184 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_73
timestamp 1669390400
transform 1 0 9520 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_75
timestamp 1669390400
transform 1 0 9744 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_78
timestamp 1669390400
transform 1 0 10080 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_85
timestamp 1669390400
transform 1 0 10864 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_91
timestamp 1669390400
transform 1 0 11536 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_95
timestamp 1669390400
transform 1 0 11984 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_111
timestamp 1669390400
transform 1 0 13776 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_115
timestamp 1669390400
transform 1 0 14224 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_118
timestamp 1669390400
transform 1 0 14560 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_132
timestamp 1669390400
transform 1 0 16128 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_134
timestamp 1669390400
transform 1 0 16352 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_141
timestamp 1669390400
transform 1 0 17136 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_144
timestamp 1669390400
transform 1 0 17472 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_151
timestamp 1669390400
transform 1 0 18256 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_161
timestamp 1669390400
transform 1 0 19376 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_165
timestamp 1669390400
transform 1 0 19824 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_173
timestamp 1669390400
transform 1 0 20720 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_175
timestamp 1669390400
transform 1 0 20944 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_191
timestamp 1669390400
transform 1 0 22736 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_212
timestamp 1669390400
transform 1 0 25088 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_215
timestamp 1669390400
transform 1 0 25424 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_219
timestamp 1669390400
transform 1 0 25872 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_239
timestamp 1669390400
transform 1 0 28112 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_243
timestamp 1669390400
transform 1 0 28560 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_254
timestamp 1669390400
transform 1 0 29792 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_266
timestamp 1669390400
transform 1 0 31136 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_272
timestamp 1669390400
transform 1 0 31808 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_276
timestamp 1669390400
transform 1 0 32256 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_283
timestamp 1669390400
transform 1 0 33040 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_286
timestamp 1669390400
transform 1 0 33376 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_297
timestamp 1669390400
transform 1 0 34608 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_301
timestamp 1669390400
transform 1 0 35056 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_305
timestamp 1669390400
transform 1 0 35504 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_316
timestamp 1669390400
transform 1 0 36736 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_323
timestamp 1669390400
transform 1 0 37520 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_327
timestamp 1669390400
transform 1 0 37968 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_331
timestamp 1669390400
transform 1 0 38416 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_333
timestamp 1669390400
transform 1 0 38640 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_340
timestamp 1669390400
transform 1 0 39424 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_352
timestamp 1669390400
transform 1 0 40768 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_354
timestamp 1669390400
transform 1 0 40992 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_357
timestamp 1669390400
transform 1 0 41328 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_360
timestamp 1669390400
transform 1 0 41664 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_364
timestamp 1669390400
transform 1 0 42112 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_370
timestamp 1669390400
transform 1 0 42784 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_382
timestamp 1669390400
transform 1 0 44128 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_392
timestamp 1669390400
transform 1 0 45248 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_406
timestamp 1669390400
transform 1 0 46816 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_416
timestamp 1669390400
transform 1 0 47936 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_423
timestamp 1669390400
transform 1 0 48720 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_425
timestamp 1669390400
transform 1 0 48944 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_428
timestamp 1669390400
transform 1 0 49280 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_441
timestamp 1669390400
transform 1 0 50736 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_451
timestamp 1669390400
transform 1 0 51856 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_455
timestamp 1669390400
transform 1 0 52304 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_463
timestamp 1669390400
transform 1 0 53200 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_473
timestamp 1669390400
transform 1 0 54320 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_477
timestamp 1669390400
transform 1 0 54768 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_486
timestamp 1669390400
transform 1 0 55776 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_496
timestamp 1669390400
transform 1 0 56896 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_499
timestamp 1669390400
transform 1 0 57232 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_508
timestamp 1669390400
transform 1 0 58240 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_512
timestamp 1669390400
transform 1 0 58688 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_2
timestamp 1669390400
transform 1 0 1568 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_5
timestamp 1669390400
transform 1 0 1904 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_9
timestamp 1669390400
transform 1 0 2352 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_13
timestamp 1669390400
transform 1 0 2800 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_17
timestamp 1669390400
transform 1 0 3248 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_21
timestamp 1669390400
transform 1 0 3696 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_25
timestamp 1669390400
transform 1 0 4144 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_29
timestamp 1669390400
transform 1 0 4592 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_33
timestamp 1669390400
transform 1 0 5040 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_37
timestamp 1669390400
transform 1 0 5488 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_43
timestamp 1669390400
transform 1 0 6160 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_47
timestamp 1669390400
transform 1 0 6608 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_51
timestamp 1669390400
transform 1 0 7056 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_66
timestamp 1669390400
transform 1 0 8736 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_76
timestamp 1669390400
transform 1 0 9856 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_80
timestamp 1669390400
transform 1 0 10304 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_84
timestamp 1669390400
transform 1 0 10752 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_86
timestamp 1669390400
transform 1 0 10976 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_89
timestamp 1669390400
transform 1 0 11312 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_93
timestamp 1669390400
transform 1 0 11760 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_103
timestamp 1669390400
transform 1 0 12880 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_105
timestamp 1669390400
transform 1 0 13104 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_108
timestamp 1669390400
transform 1 0 13440 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_114
timestamp 1669390400
transform 1 0 14112 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_118
timestamp 1669390400
transform 1 0 14560 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_121
timestamp 1669390400
transform 1 0 14896 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_125
timestamp 1669390400
transform 1 0 15344 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_129
timestamp 1669390400
transform 1 0 15792 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_145
timestamp 1669390400
transform 1 0 17584 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_159
timestamp 1669390400
transform 1 0 19152 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_169
timestamp 1669390400
transform 1 0 20272 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_176
timestamp 1669390400
transform 1 0 21056 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_179
timestamp 1669390400
transform 1 0 21392 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_186
timestamp 1669390400
transform 1 0 22176 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_188
timestamp 1669390400
transform 1 0 22400 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_191
timestamp 1669390400
transform 1 0 22736 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_201
timestamp 1669390400
transform 1 0 23856 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_229
timestamp 1669390400
transform 1 0 26992 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_239
timestamp 1669390400
transform 1 0 28112 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_243
timestamp 1669390400
transform 1 0 28560 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_247
timestamp 1669390400
transform 1 0 29008 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_250
timestamp 1669390400
transform 1 0 29344 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_254
timestamp 1669390400
transform 1 0 29792 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_266
timestamp 1669390400
transform 1 0 31136 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_272
timestamp 1669390400
transform 1 0 31808 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_274
timestamp 1669390400
transform 1 0 32032 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_277
timestamp 1669390400
transform 1 0 32368 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_281
timestamp 1669390400
transform 1 0 32816 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_285
timestamp 1669390400
transform 1 0 33264 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_296
timestamp 1669390400
transform 1 0 34496 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_300
timestamp 1669390400
transform 1 0 34944 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_304
timestamp 1669390400
transform 1 0 35392 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_308
timestamp 1669390400
transform 1 0 35840 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_312
timestamp 1669390400
transform 1 0 36288 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_316
timestamp 1669390400
transform 1 0 36736 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_318
timestamp 1669390400
transform 1 0 36960 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_321
timestamp 1669390400
transform 1 0 37296 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_324
timestamp 1669390400
transform 1 0 37632 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_328
timestamp 1669390400
transform 1 0 38080 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_332
timestamp 1669390400
transform 1 0 38528 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_336
timestamp 1669390400
transform 1 0 38976 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_340
timestamp 1669390400
transform 1 0 39424 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_344
timestamp 1669390400
transform 1 0 39872 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_352
timestamp 1669390400
transform 1 0 40768 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_356
timestamp 1669390400
transform 1 0 41216 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_360
timestamp 1669390400
transform 1 0 41664 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_364
timestamp 1669390400
transform 1 0 42112 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_368
timestamp 1669390400
transform 1 0 42560 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_372
timestamp 1669390400
transform 1 0 43008 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_376
timestamp 1669390400
transform 1 0 43456 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_382
timestamp 1669390400
transform 1 0 44128 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_389
timestamp 1669390400
transform 1 0 44912 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_392
timestamp 1669390400
transform 1 0 45248 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_402
timestamp 1669390400
transform 1 0 46368 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_410
timestamp 1669390400
transform 1 0 47264 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_416
timestamp 1669390400
transform 1 0 47936 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_420
timestamp 1669390400
transform 1 0 48384 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_424
timestamp 1669390400
transform 1 0 48832 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_432
timestamp 1669390400
transform 1 0 49728 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_434
timestamp 1669390400
transform 1 0 49952 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_447
timestamp 1669390400
transform 1 0 51408 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_457
timestamp 1669390400
transform 1 0 52528 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_463
timestamp 1669390400
transform 1 0 53200 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_482
timestamp 1669390400
transform 1 0 55328 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_512
timestamp 1669390400
transform 1 0 58688 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_2
timestamp 1669390400
transform 1 0 1568 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_4
timestamp 1669390400
transform 1 0 1792 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_7
timestamp 1669390400
transform 1 0 2128 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_11
timestamp 1669390400
transform 1 0 2576 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_15
timestamp 1669390400
transform 1 0 3024 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_19
timestamp 1669390400
transform 1 0 3472 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_23
timestamp 1669390400
transform 1 0 3920 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_27
timestamp 1669390400
transform 1 0 4368 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_31
timestamp 1669390400
transform 1 0 4816 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_35
timestamp 1669390400
transform 1 0 5264 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_39
timestamp 1669390400
transform 1 0 5712 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_43
timestamp 1669390400
transform 1 0 6160 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_55
timestamp 1669390400
transform 1 0 7504 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_70
timestamp 1669390400
transform 1 0 9184 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_73
timestamp 1669390400
transform 1 0 9520 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_76
timestamp 1669390400
transform 1 0 9856 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_80
timestamp 1669390400
transform 1 0 10304 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_86
timestamp 1669390400
transform 1 0 10976 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_90
timestamp 1669390400
transform 1 0 11424 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_94
timestamp 1669390400
transform 1 0 11872 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_98
timestamp 1669390400
transform 1 0 12320 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_105
timestamp 1669390400
transform 1 0 13104 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_107
timestamp 1669390400
transform 1 0 13328 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_110
timestamp 1669390400
transform 1 0 13664 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_114
timestamp 1669390400
transform 1 0 14112 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_118
timestamp 1669390400
transform 1 0 14560 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_120
timestamp 1669390400
transform 1 0 14784 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_123
timestamp 1669390400
transform 1 0 15120 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_133
timestamp 1669390400
transform 1 0 16240 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_141
timestamp 1669390400
transform 1 0 17136 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_144
timestamp 1669390400
transform 1 0 17472 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_151
timestamp 1669390400
transform 1 0 18256 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_155
timestamp 1669390400
transform 1 0 18704 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_159
timestamp 1669390400
transform 1 0 19152 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_163
timestamp 1669390400
transform 1 0 19600 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_167
timestamp 1669390400
transform 1 0 20048 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_175
timestamp 1669390400
transform 1 0 20944 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_203
timestamp 1669390400
transform 1 0 24080 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_212
timestamp 1669390400
transform 1 0 25088 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_215
timestamp 1669390400
transform 1 0 25424 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_228
timestamp 1669390400
transform 1 0 26880 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_256
timestamp 1669390400
transform 1 0 30016 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_270
timestamp 1669390400
transform 1 0 31584 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_281
timestamp 1669390400
transform 1 0 32816 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_283
timestamp 1669390400
transform 1 0 33040 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_286
timestamp 1669390400
transform 1 0 33376 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_289
timestamp 1669390400
transform 1 0 33712 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_293
timestamp 1669390400
transform 1 0 34160 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_303
timestamp 1669390400
transform 1 0 35280 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_313
timestamp 1669390400
transform 1 0 36400 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_321
timestamp 1669390400
transform 1 0 37296 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_323
timestamp 1669390400
transform 1 0 37520 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_336
timestamp 1669390400
transform 1 0 38976 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_340
timestamp 1669390400
transform 1 0 39424 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_350
timestamp 1669390400
transform 1 0 40544 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_354
timestamp 1669390400
transform 1 0 40992 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_357
timestamp 1669390400
transform 1 0 41328 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_370
timestamp 1669390400
transform 1 0 42784 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_384
timestamp 1669390400
transform 1 0 44352 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_398
timestamp 1669390400
transform 1 0 45920 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_400
timestamp 1669390400
transform 1 0 46144 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_403
timestamp 1669390400
transform 1 0 46480 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_417
timestamp 1669390400
transform 1 0 48048 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_421
timestamp 1669390400
transform 1 0 48496 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_425
timestamp 1669390400
transform 1 0 48944 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_428
timestamp 1669390400
transform 1 0 49280 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_436
timestamp 1669390400
transform 1 0 50176 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_440
timestamp 1669390400
transform 1 0 50624 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_447
timestamp 1669390400
transform 1 0 51408 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_468
timestamp 1669390400
transform 1 0 53760 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_483
timestamp 1669390400
transform 1 0 55440 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_487
timestamp 1669390400
transform 1 0 55888 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_491
timestamp 1669390400
transform 1 0 56336 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_495
timestamp 1669390400
transform 1 0 56784 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_499
timestamp 1669390400
transform 1 0 57232 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_507
timestamp 1669390400
transform 1 0 58128 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_511
timestamp 1669390400
transform 1 0 58576 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_2
timestamp 1669390400
transform 1 0 1568 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_6
timestamp 1669390400
transform 1 0 2016 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_10
timestamp 1669390400
transform 1 0 2464 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_14
timestamp 1669390400
transform 1 0 2912 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_18
timestamp 1669390400
transform 1 0 3360 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_22
timestamp 1669390400
transform 1 0 3808 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_26
timestamp 1669390400
transform 1 0 4256 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_30
timestamp 1669390400
transform 1 0 4704 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_34
timestamp 1669390400
transform 1 0 5152 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_37
timestamp 1669390400
transform 1 0 5488 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_59
timestamp 1669390400
transform 1 0 7952 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_84
timestamp 1669390400
transform 1 0 10752 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_86
timestamp 1669390400
transform 1 0 10976 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_94
timestamp 1669390400
transform 1 0 11872 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_98
timestamp 1669390400
transform 1 0 12320 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_101
timestamp 1669390400
transform 1 0 12656 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_105
timestamp 1669390400
transform 1 0 13104 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_108
timestamp 1669390400
transform 1 0 13440 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_130
timestamp 1669390400
transform 1 0 15904 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_132
timestamp 1669390400
transform 1 0 16128 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_135
timestamp 1669390400
transform 1 0 16464 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_147
timestamp 1669390400
transform 1 0 17808 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_149
timestamp 1669390400
transform 1 0 18032 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_152
timestamp 1669390400
transform 1 0 18368 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_156
timestamp 1669390400
transform 1 0 18816 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_160
timestamp 1669390400
transform 1 0 19264 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_164
timestamp 1669390400
transform 1 0 19712 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_176
timestamp 1669390400
transform 1 0 21056 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_179
timestamp 1669390400
transform 1 0 21392 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_188
timestamp 1669390400
transform 1 0 22400 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_194
timestamp 1669390400
transform 1 0 23072 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_202
timestamp 1669390400
transform 1 0 23968 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_230
timestamp 1669390400
transform 1 0 27104 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_245
timestamp 1669390400
transform 1 0 28784 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_247
timestamp 1669390400
transform 1 0 29008 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_250
timestamp 1669390400
transform 1 0 29344 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_284
timestamp 1669390400
transform 1 0 33152 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_288
timestamp 1669390400
transform 1 0 33600 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_292
timestamp 1669390400
transform 1 0 34048 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_294
timestamp 1669390400
transform 1 0 34272 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_318
timestamp 1669390400
transform 1 0 36960 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_321
timestamp 1669390400
transform 1 0 37296 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_334
timestamp 1669390400
transform 1 0 38752 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_338
timestamp 1669390400
transform 1 0 39200 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_342
timestamp 1669390400
transform 1 0 39648 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_346
timestamp 1669390400
transform 1 0 40096 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_350
timestamp 1669390400
transform 1 0 40544 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_360
timestamp 1669390400
transform 1 0 41664 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_364
timestamp 1669390400
transform 1 0 42112 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_26_374
timestamp 1669390400
transform 1 0 43232 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_382
timestamp 1669390400
transform 1 0 44128 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_386
timestamp 1669390400
transform 1 0 44576 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_392
timestamp 1669390400
transform 1 0 45248 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_405
timestamp 1669390400
transform 1 0 46704 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_409
timestamp 1669390400
transform 1 0 47152 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_411
timestamp 1669390400
transform 1 0 47376 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_414
timestamp 1669390400
transform 1 0 47712 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_418
timestamp 1669390400
transform 1 0 48160 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_442
timestamp 1669390400
transform 1 0 50848 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_458
timestamp 1669390400
transform 1 0 52640 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_460
timestamp 1669390400
transform 1 0 52864 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_463
timestamp 1669390400
transform 1 0 53200 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_482
timestamp 1669390400
transform 1 0 55328 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_507
timestamp 1669390400
transform 1 0 58128 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_511
timestamp 1669390400
transform 1 0 58576 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_2
timestamp 1669390400
transform 1 0 1568 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_6
timestamp 1669390400
transform 1 0 2016 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_10
timestamp 1669390400
transform 1 0 2464 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_14
timestamp 1669390400
transform 1 0 2912 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_18
timestamp 1669390400
transform 1 0 3360 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_22
timestamp 1669390400
transform 1 0 3808 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_46
timestamp 1669390400
transform 1 0 6496 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_69
timestamp 1669390400
transform 1 0 9072 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_73
timestamp 1669390400
transform 1 0 9520 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_89
timestamp 1669390400
transform 1 0 11312 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_99
timestamp 1669390400
transform 1 0 12432 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_103
timestamp 1669390400
transform 1 0 12880 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_122
timestamp 1669390400
transform 1 0 15008 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_126
timestamp 1669390400
transform 1 0 15456 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_129
timestamp 1669390400
transform 1 0 15792 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_133
timestamp 1669390400
transform 1 0 16240 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_137
timestamp 1669390400
transform 1 0 16688 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_141
timestamp 1669390400
transform 1 0 17136 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_144
timestamp 1669390400
transform 1 0 17472 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_157
timestamp 1669390400
transform 1 0 18928 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_167
timestamp 1669390400
transform 1 0 20048 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_187
timestamp 1669390400
transform 1 0 22288 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_189
timestamp 1669390400
transform 1 0 22512 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1669390400
transform 1 0 25088 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_215
timestamp 1669390400
transform 1 0 25424 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_219
timestamp 1669390400
transform 1 0 25872 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_238
timestamp 1669390400
transform 1 0 28000 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_249
timestamp 1669390400
transform 1 0 29232 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_253
timestamp 1669390400
transform 1 0 29680 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_257
timestamp 1669390400
transform 1 0 30128 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_261
timestamp 1669390400
transform 1 0 30576 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_265
timestamp 1669390400
transform 1 0 31024 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_269
timestamp 1669390400
transform 1 0 31472 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_273
timestamp 1669390400
transform 1 0 31920 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_276
timestamp 1669390400
transform 1 0 32256 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_280
timestamp 1669390400
transform 1 0 32704 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_286
timestamp 1669390400
transform 1 0 33376 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_303
timestamp 1669390400
transform 1 0 35280 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_313
timestamp 1669390400
transform 1 0 36400 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_317
timestamp 1669390400
transform 1 0 36848 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_343
timestamp 1669390400
transform 1 0 39760 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_347
timestamp 1669390400
transform 1 0 40208 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_351
timestamp 1669390400
transform 1 0 40656 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_357
timestamp 1669390400
transform 1 0 41328 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_360
timestamp 1669390400
transform 1 0 41664 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_364
timestamp 1669390400
transform 1 0 42112 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_368
timestamp 1669390400
transform 1 0 42560 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_382
timestamp 1669390400
transform 1 0 44128 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_386
timestamp 1669390400
transform 1 0 44576 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_388
timestamp 1669390400
transform 1 0 44800 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_391
timestamp 1669390400
transform 1 0 45136 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_395
timestamp 1669390400
transform 1 0 45584 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_412
timestamp 1669390400
transform 1 0 47488 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_416
timestamp 1669390400
transform 1 0 47936 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_425
timestamp 1669390400
transform 1 0 48944 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_428
timestamp 1669390400
transform 1 0 49280 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_438
timestamp 1669390400
transform 1 0 50400 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_454
timestamp 1669390400
transform 1 0 52192 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_466
timestamp 1669390400
transform 1 0 53536 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_487
timestamp 1669390400
transform 1 0 55888 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_495
timestamp 1669390400
transform 1 0 56784 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_499
timestamp 1669390400
transform 1 0 57232 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_508
timestamp 1669390400
transform 1 0 58240 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_512
timestamp 1669390400
transform 1 0 58688 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_2
timestamp 1669390400
transform 1 0 1568 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_4
timestamp 1669390400
transform 1 0 1792 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_7
timestamp 1669390400
transform 1 0 2128 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_11
timestamp 1669390400
transform 1 0 2576 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_15
timestamp 1669390400
transform 1 0 3024 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_34
timestamp 1669390400
transform 1 0 5152 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_37
timestamp 1669390400
transform 1 0 5488 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_41
timestamp 1669390400
transform 1 0 5936 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_51
timestamp 1669390400
transform 1 0 7056 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_63
timestamp 1669390400
transform 1 0 8400 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_65
timestamp 1669390400
transform 1 0 8624 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_68
timestamp 1669390400
transform 1 0 8960 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_72
timestamp 1669390400
transform 1 0 9408 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_76
timestamp 1669390400
transform 1 0 9856 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_86
timestamp 1669390400
transform 1 0 10976 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_97
timestamp 1669390400
transform 1 0 12208 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_101
timestamp 1669390400
transform 1 0 12656 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_105
timestamp 1669390400
transform 1 0 13104 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_108
timestamp 1669390400
transform 1 0 13440 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_112
timestamp 1669390400
transform 1 0 13888 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_116
timestamp 1669390400
transform 1 0 14336 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_136
timestamp 1669390400
transform 1 0 16576 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_138
timestamp 1669390400
transform 1 0 16800 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_141
timestamp 1669390400
transform 1 0 17136 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_161
timestamp 1669390400
transform 1 0 19376 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_173
timestamp 1669390400
transform 1 0 20720 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_179
timestamp 1669390400
transform 1 0 21392 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_181
timestamp 1669390400
transform 1 0 21616 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_190
timestamp 1669390400
transform 1 0 22624 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_192
timestamp 1669390400
transform 1 0 22848 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_195
timestamp 1669390400
transform 1 0 23184 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_199
timestamp 1669390400
transform 1 0 23632 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_223
timestamp 1669390400
transform 1 0 26320 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_229
timestamp 1669390400
transform 1 0 26992 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_245
timestamp 1669390400
transform 1 0 28784 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_247
timestamp 1669390400
transform 1 0 29008 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_250
timestamp 1669390400
transform 1 0 29344 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_256
timestamp 1669390400
transform 1 0 30016 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_268
timestamp 1669390400
transform 1 0 31360 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_287
timestamp 1669390400
transform 1 0 33488 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_301
timestamp 1669390400
transform 1 0 35056 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_311
timestamp 1669390400
transform 1 0 36176 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_315
timestamp 1669390400
transform 1 0 36624 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_321
timestamp 1669390400
transform 1 0 37296 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_324
timestamp 1669390400
transform 1 0 37632 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_328
timestamp 1669390400
transform 1 0 38080 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_332
timestamp 1669390400
transform 1 0 38528 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_336
timestamp 1669390400
transform 1 0 38976 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_340
timestamp 1669390400
transform 1 0 39424 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_344
timestamp 1669390400
transform 1 0 39872 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_361
timestamp 1669390400
transform 1 0 41776 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_376
timestamp 1669390400
transform 1 0 43456 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_384
timestamp 1669390400
transform 1 0 44352 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_388
timestamp 1669390400
transform 1 0 44800 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_392
timestamp 1669390400
transform 1 0 45248 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_399
timestamp 1669390400
transform 1 0 46032 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_403
timestamp 1669390400
transform 1 0 46480 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_420
timestamp 1669390400
transform 1 0 48384 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_434
timestamp 1669390400
transform 1 0 49952 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_444
timestamp 1669390400
transform 1 0 51072 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_448
timestamp 1669390400
transform 1 0 51520 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_456
timestamp 1669390400
transform 1 0 52416 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_460
timestamp 1669390400
transform 1 0 52864 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_463
timestamp 1669390400
transform 1 0 53200 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_476
timestamp 1669390400
transform 1 0 54656 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_490
timestamp 1669390400
transform 1 0 56224 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_494
timestamp 1669390400
transform 1 0 56672 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_508
timestamp 1669390400
transform 1 0 58240 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_512
timestamp 1669390400
transform 1 0 58688 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_2
timestamp 1669390400
transform 1 0 1568 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_4
timestamp 1669390400
transform 1 0 1792 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_7
timestamp 1669390400
transform 1 0 2128 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_11
timestamp 1669390400
transform 1 0 2576 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_15
timestamp 1669390400
transform 1 0 3024 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_19
timestamp 1669390400
transform 1 0 3472 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_23
timestamp 1669390400
transform 1 0 3920 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_27
timestamp 1669390400
transform 1 0 4368 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_47
timestamp 1669390400
transform 1 0 6608 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_70
timestamp 1669390400
transform 1 0 9184 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_73
timestamp 1669390400
transform 1 0 9520 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_77
timestamp 1669390400
transform 1 0 9968 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_81
timestamp 1669390400
transform 1 0 10416 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_94
timestamp 1669390400
transform 1 0 11872 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_98
timestamp 1669390400
transform 1 0 12320 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_118
timestamp 1669390400
transform 1 0 14560 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_120
timestamp 1669390400
transform 1 0 14784 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_138
timestamp 1669390400
transform 1 0 16800 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_144
timestamp 1669390400
transform 1 0 17472 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_170
timestamp 1669390400
transform 1 0 20384 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_176
timestamp 1669390400
transform 1 0 21056 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_195
timestamp 1669390400
transform 1 0 23184 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_202
timestamp 1669390400
transform 1 0 23968 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_208
timestamp 1669390400
transform 1 0 24640 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1669390400
transform 1 0 25088 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_215
timestamp 1669390400
transform 1 0 25424 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_224
timestamp 1669390400
transform 1 0 26432 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_226
timestamp 1669390400
transform 1 0 26656 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_236
timestamp 1669390400
transform 1 0 27776 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_247
timestamp 1669390400
transform 1 0 29008 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_261
timestamp 1669390400
transform 1 0 30576 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_265
timestamp 1669390400
transform 1 0 31024 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_269
timestamp 1669390400
transform 1 0 31472 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_273
timestamp 1669390400
transform 1 0 31920 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_277
timestamp 1669390400
transform 1 0 32368 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_283
timestamp 1669390400
transform 1 0 33040 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_286
timestamp 1669390400
transform 1 0 33376 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_296
timestamp 1669390400
transform 1 0 34496 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_306
timestamp 1669390400
transform 1 0 35616 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_310
timestamp 1669390400
transform 1 0 36064 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_314
timestamp 1669390400
transform 1 0 36512 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_318
timestamp 1669390400
transform 1 0 36960 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_322
timestamp 1669390400
transform 1 0 37408 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_326
timestamp 1669390400
transform 1 0 37856 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_330
timestamp 1669390400
transform 1 0 38304 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_334
timestamp 1669390400
transform 1 0 38752 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_336
timestamp 1669390400
transform 1 0 38976 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_353
timestamp 1669390400
transform 1 0 40880 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_357
timestamp 1669390400
transform 1 0 41328 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_370
timestamp 1669390400
transform 1 0 42784 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_372
timestamp 1669390400
transform 1 0 43008 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_381
timestamp 1669390400
transform 1 0 44016 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_385
timestamp 1669390400
transform 1 0 44464 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_389
timestamp 1669390400
transform 1 0 44912 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_397
timestamp 1669390400
transform 1 0 45808 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_401
timestamp 1669390400
transform 1 0 46256 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_405
timestamp 1669390400
transform 1 0 46704 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_409
timestamp 1669390400
transform 1 0 47152 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_413
timestamp 1669390400
transform 1 0 47600 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_417
timestamp 1669390400
transform 1 0 48048 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_421
timestamp 1669390400
transform 1 0 48496 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_425
timestamp 1669390400
transform 1 0 48944 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_428
timestamp 1669390400
transform 1 0 49280 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_431
timestamp 1669390400
transform 1 0 49616 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_435
timestamp 1669390400
transform 1 0 50064 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_439
timestamp 1669390400
transform 1 0 50512 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_447
timestamp 1669390400
transform 1 0 51408 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_451
timestamp 1669390400
transform 1 0 51856 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_455
timestamp 1669390400
transform 1 0 52304 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_470
timestamp 1669390400
transform 1 0 53984 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_478
timestamp 1669390400
transform 1 0 54880 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_486
timestamp 1669390400
transform 1 0 55776 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_496
timestamp 1669390400
transform 1 0 56896 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_499
timestamp 1669390400
transform 1 0 57232 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_512
timestamp 1669390400
transform 1 0 58688 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_2
timestamp 1669390400
transform 1 0 1568 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_6
timestamp 1669390400
transform 1 0 2016 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_30
timestamp 1669390400
transform 1 0 4704 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_34
timestamp 1669390400
transform 1 0 5152 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_37
timestamp 1669390400
transform 1 0 5488 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_56
timestamp 1669390400
transform 1 0 7616 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_58
timestamp 1669390400
transform 1 0 7840 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_61
timestamp 1669390400
transform 1 0 8176 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_65
timestamp 1669390400
transform 1 0 8624 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_77
timestamp 1669390400
transform 1 0 9968 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_79
timestamp 1669390400
transform 1 0 10192 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_82
timestamp 1669390400
transform 1 0 10528 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_92
timestamp 1669390400
transform 1 0 11648 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_102
timestamp 1669390400
transform 1 0 12768 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_108
timestamp 1669390400
transform 1 0 13440 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_120
timestamp 1669390400
transform 1 0 14784 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_126
timestamp 1669390400
transform 1 0 15456 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_130
timestamp 1669390400
transform 1 0 15904 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_169
timestamp 1669390400
transform 1 0 20272 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_173
timestamp 1669390400
transform 1 0 20720 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_176
timestamp 1669390400
transform 1 0 21056 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_179
timestamp 1669390400
transform 1 0 21392 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_196
timestamp 1669390400
transform 1 0 23296 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_212
timestamp 1669390400
transform 1 0 25088 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_226
timestamp 1669390400
transform 1 0 26656 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_236
timestamp 1669390400
transform 1 0 27776 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_247
timestamp 1669390400
transform 1 0 29008 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_250
timestamp 1669390400
transform 1 0 29344 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_253
timestamp 1669390400
transform 1 0 29680 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_257
timestamp 1669390400
transform 1 0 30128 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_259
timestamp 1669390400
transform 1 0 30352 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_307
timestamp 1669390400
transform 1 0 35728 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_318
timestamp 1669390400
transform 1 0 36960 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_321
timestamp 1669390400
transform 1 0 37296 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_348
timestamp 1669390400
transform 1 0 40320 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_355
timestamp 1669390400
transform 1 0 41104 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_359
timestamp 1669390400
transform 1 0 41552 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_363
timestamp 1669390400
transform 1 0 42000 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_367
timestamp 1669390400
transform 1 0 42448 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_371
timestamp 1669390400
transform 1 0 42896 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_375
timestamp 1669390400
transform 1 0 43344 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_379
timestamp 1669390400
transform 1 0 43792 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_383
timestamp 1669390400
transform 1 0 44240 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_387
timestamp 1669390400
transform 1 0 44688 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_389
timestamp 1669390400
transform 1 0 44912 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_392
timestamp 1669390400
transform 1 0 45248 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_404
timestamp 1669390400
transform 1 0 46592 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_416
timestamp 1669390400
transform 1 0 47936 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_423
timestamp 1669390400
transform 1 0 48720 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_427
timestamp 1669390400
transform 1 0 49168 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_435
timestamp 1669390400
transform 1 0 50064 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_449
timestamp 1669390400
transform 1 0 51632 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_451
timestamp 1669390400
transform 1 0 51856 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_454
timestamp 1669390400
transform 1 0 52192 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_460
timestamp 1669390400
transform 1 0 52864 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_463
timestamp 1669390400
transform 1 0 53200 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_472
timestamp 1669390400
transform 1 0 54208 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_488
timestamp 1669390400
transform 1 0 56000 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_496
timestamp 1669390400
transform 1 0 56896 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_510
timestamp 1669390400
transform 1 0 58464 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_512
timestamp 1669390400
transform 1 0 58688 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_2
timestamp 1669390400
transform 1 0 1568 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_6
timestamp 1669390400
transform 1 0 2016 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_30
timestamp 1669390400
transform 1 0 4704 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_44
timestamp 1669390400
transform 1 0 6272 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_70
timestamp 1669390400
transform 1 0 9184 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_73
timestamp 1669390400
transform 1 0 9520 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_101
timestamp 1669390400
transform 1 0 12656 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_105
timestamp 1669390400
transform 1 0 13104 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_108
timestamp 1669390400
transform 1 0 13440 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_112
timestamp 1669390400
transform 1 0 13888 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_116
timestamp 1669390400
transform 1 0 14336 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_131
timestamp 1669390400
transform 1 0 16016 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_137
timestamp 1669390400
transform 1 0 16688 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_141
timestamp 1669390400
transform 1 0 17136 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_144
timestamp 1669390400
transform 1 0 17472 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_150
timestamp 1669390400
transform 1 0 18144 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_171
timestamp 1669390400
transform 1 0 20496 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_183
timestamp 1669390400
transform 1 0 21840 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_185
timestamp 1669390400
transform 1 0 22064 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_188
timestamp 1669390400
transform 1 0 22400 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_192
timestamp 1669390400
transform 1 0 22848 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_196
timestamp 1669390400
transform 1 0 23296 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_200
timestamp 1669390400
transform 1 0 23744 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_204
timestamp 1669390400
transform 1 0 24192 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_208
timestamp 1669390400
transform 1 0 24640 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1669390400
transform 1 0 25088 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_215
timestamp 1669390400
transform 1 0 25424 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_222
timestamp 1669390400
transform 1 0 26208 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_226
timestamp 1669390400
transform 1 0 26656 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_246
timestamp 1669390400
transform 1 0 28896 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_252
timestamp 1669390400
transform 1 0 29568 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_278
timestamp 1669390400
transform 1 0 32480 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_282
timestamp 1669390400
transform 1 0 32928 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_286
timestamp 1669390400
transform 1 0 33376 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_297
timestamp 1669390400
transform 1 0 34608 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_301
timestamp 1669390400
transform 1 0 35056 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_314
timestamp 1669390400
transform 1 0 36512 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_316
timestamp 1669390400
transform 1 0 36736 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_326
timestamp 1669390400
transform 1 0 37856 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_330
timestamp 1669390400
transform 1 0 38304 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_334
timestamp 1669390400
transform 1 0 38752 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_347
timestamp 1669390400
transform 1 0 40208 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_351
timestamp 1669390400
transform 1 0 40656 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_357
timestamp 1669390400
transform 1 0 41328 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_360
timestamp 1669390400
transform 1 0 41664 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_364
timestamp 1669390400
transform 1 0 42112 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_366
timestamp 1669390400
transform 1 0 42336 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_391
timestamp 1669390400
transform 1 0 45136 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_393
timestamp 1669390400
transform 1 0 45360 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_400
timestamp 1669390400
transform 1 0 46144 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_416
timestamp 1669390400
transform 1 0 47936 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_420
timestamp 1669390400
transform 1 0 48384 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_424
timestamp 1669390400
transform 1 0 48832 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_428
timestamp 1669390400
transform 1 0 49280 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_452
timestamp 1669390400
transform 1 0 51968 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_466
timestamp 1669390400
transform 1 0 53536 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_482
timestamp 1669390400
transform 1 0 55328 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_490
timestamp 1669390400
transform 1 0 56224 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_494
timestamp 1669390400
transform 1 0 56672 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_496
timestamp 1669390400
transform 1 0 56896 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_499
timestamp 1669390400
transform 1 0 57232 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_507
timestamp 1669390400
transform 1 0 58128 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_511
timestamp 1669390400
transform 1 0 58576 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_2
timestamp 1669390400
transform 1 0 1568 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_4
timestamp 1669390400
transform 1 0 1792 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_7
timestamp 1669390400
transform 1 0 2128 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_26
timestamp 1669390400
transform 1 0 4256 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_30
timestamp 1669390400
transform 1 0 4704 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_34
timestamp 1669390400
transform 1 0 5152 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_37
timestamp 1669390400
transform 1 0 5488 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_39
timestamp 1669390400
transform 1 0 5712 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_42
timestamp 1669390400
transform 1 0 6048 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_46
timestamp 1669390400
transform 1 0 6496 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_64
timestamp 1669390400
transform 1 0 8512 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_68
timestamp 1669390400
transform 1 0 8960 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_77
timestamp 1669390400
transform 1 0 9968 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_89
timestamp 1669390400
transform 1 0 11312 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_95
timestamp 1669390400
transform 1 0 11984 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_105
timestamp 1669390400
transform 1 0 13104 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_108
timestamp 1669390400
transform 1 0 13440 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_111
timestamp 1669390400
transform 1 0 13776 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_130
timestamp 1669390400
transform 1 0 15904 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_134
timestamp 1669390400
transform 1 0 16352 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_149
timestamp 1669390400
transform 1 0 18032 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_167
timestamp 1669390400
transform 1 0 20048 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_169
timestamp 1669390400
transform 1 0 20272 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_172
timestamp 1669390400
transform 1 0 20608 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_176
timestamp 1669390400
transform 1 0 21056 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_179
timestamp 1669390400
transform 1 0 21392 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_190
timestamp 1669390400
transform 1 0 22624 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_210
timestamp 1669390400
transform 1 0 24864 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_212
timestamp 1669390400
transform 1 0 25088 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_215
timestamp 1669390400
transform 1 0 25424 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_219
timestamp 1669390400
transform 1 0 25872 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_231
timestamp 1669390400
transform 1 0 27216 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_245
timestamp 1669390400
transform 1 0 28784 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_247
timestamp 1669390400
transform 1 0 29008 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_250
timestamp 1669390400
transform 1 0 29344 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_260
timestamp 1669390400
transform 1 0 30464 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_287
timestamp 1669390400
transform 1 0 33488 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_304
timestamp 1669390400
transform 1 0 35392 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_306
timestamp 1669390400
transform 1 0 35616 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_313
timestamp 1669390400
transform 1 0 36400 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_317
timestamp 1669390400
transform 1 0 36848 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_321
timestamp 1669390400
transform 1 0 37296 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_324
timestamp 1669390400
transform 1 0 37632 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_328
timestamp 1669390400
transform 1 0 38080 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_332
timestamp 1669390400
transform 1 0 38528 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_336
timestamp 1669390400
transform 1 0 38976 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_338
timestamp 1669390400
transform 1 0 39200 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_346
timestamp 1669390400
transform 1 0 40096 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_350
timestamp 1669390400
transform 1 0 40544 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_354
timestamp 1669390400
transform 1 0 40992 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_363
timestamp 1669390400
transform 1 0 42000 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_373
timestamp 1669390400
transform 1 0 43120 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_383
timestamp 1669390400
transform 1 0 44240 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_387
timestamp 1669390400
transform 1 0 44688 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_389
timestamp 1669390400
transform 1 0 44912 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_392
timestamp 1669390400
transform 1 0 45248 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_395
timestamp 1669390400
transform 1 0 45584 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_399
timestamp 1669390400
transform 1 0 46032 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_403
timestamp 1669390400
transform 1 0 46480 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_420
timestamp 1669390400
transform 1 0 48384 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_424
timestamp 1669390400
transform 1 0 48832 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_430
timestamp 1669390400
transform 1 0 49504 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_440
timestamp 1669390400
transform 1 0 50624 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_448
timestamp 1669390400
transform 1 0 51520 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_460
timestamp 1669390400
transform 1 0 52864 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_463
timestamp 1669390400
transform 1 0 53200 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_466
timestamp 1669390400
transform 1 0 53536 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_470
timestamp 1669390400
transform 1 0 53984 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_474
timestamp 1669390400
transform 1 0 54432 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_500
timestamp 1669390400
transform 1 0 57344 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_510
timestamp 1669390400
transform 1 0 58464 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_512
timestamp 1669390400
transform 1 0 58688 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_2
timestamp 1669390400
transform 1 0 1568 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_4
timestamp 1669390400
transform 1 0 1792 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_22
timestamp 1669390400
transform 1 0 3808 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_39
timestamp 1669390400
transform 1 0 5712 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_43
timestamp 1669390400
transform 1 0 6160 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_69
timestamp 1669390400
transform 1 0 9072 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_73
timestamp 1669390400
transform 1 0 9520 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_79
timestamp 1669390400
transform 1 0 10192 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_94
timestamp 1669390400
transform 1 0 11872 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_98
timestamp 1669390400
transform 1 0 12320 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_108
timestamp 1669390400
transform 1 0 13440 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_120
timestamp 1669390400
transform 1 0 14784 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_127
timestamp 1669390400
transform 1 0 15568 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_133
timestamp 1669390400
transform 1 0 16240 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_137
timestamp 1669390400
transform 1 0 16688 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_141
timestamp 1669390400
transform 1 0 17136 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_144
timestamp 1669390400
transform 1 0 17472 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_146
timestamp 1669390400
transform 1 0 17696 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_153
timestamp 1669390400
transform 1 0 18480 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_157
timestamp 1669390400
transform 1 0 18928 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_165
timestamp 1669390400
transform 1 0 19824 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_167
timestamp 1669390400
transform 1 0 20048 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_185
timestamp 1669390400
transform 1 0 22064 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_187
timestamp 1669390400
transform 1 0 22288 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_190
timestamp 1669390400
transform 1 0 22624 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_210
timestamp 1669390400
transform 1 0 24864 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1669390400
transform 1 0 25088 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_215
timestamp 1669390400
transform 1 0 25424 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_226
timestamp 1669390400
transform 1 0 26656 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_233
timestamp 1669390400
transform 1 0 27440 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_250
timestamp 1669390400
transform 1 0 29344 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_256
timestamp 1669390400
transform 1 0 30016 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_283
timestamp 1669390400
transform 1 0 33040 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_286
timestamp 1669390400
transform 1 0 33376 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_293
timestamp 1669390400
transform 1 0 34160 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_304
timestamp 1669390400
transform 1 0 35392 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_311
timestamp 1669390400
transform 1 0 36176 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_315
timestamp 1669390400
transform 1 0 36624 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_319
timestamp 1669390400
transform 1 0 37072 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_333
timestamp 1669390400
transform 1 0 38640 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_337
timestamp 1669390400
transform 1 0 39088 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_341
timestamp 1669390400
transform 1 0 39536 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_354
timestamp 1669390400
transform 1 0 40992 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_357
timestamp 1669390400
transform 1 0 41328 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_370
timestamp 1669390400
transform 1 0 42784 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_378
timestamp 1669390400
transform 1 0 43680 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_382
timestamp 1669390400
transform 1 0 44128 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_386
timestamp 1669390400
transform 1 0 44576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_390
timestamp 1669390400
transform 1 0 45024 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_393
timestamp 1669390400
transform 1 0 45360 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_397
timestamp 1669390400
transform 1 0 45808 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_405
timestamp 1669390400
transform 1 0 46704 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_409
timestamp 1669390400
transform 1 0 47152 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_413
timestamp 1669390400
transform 1 0 47600 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_416
timestamp 1669390400
transform 1 0 47936 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_424
timestamp 1669390400
transform 1 0 48832 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_428
timestamp 1669390400
transform 1 0 49280 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_444
timestamp 1669390400
transform 1 0 51072 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_448
timestamp 1669390400
transform 1 0 51520 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_450
timestamp 1669390400
transform 1 0 51744 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_463
timestamp 1669390400
transform 1 0 53200 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_477
timestamp 1669390400
transform 1 0 54768 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_487
timestamp 1669390400
transform 1 0 55888 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_491
timestamp 1669390400
transform 1 0 56336 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_493
timestamp 1669390400
transform 1 0 56560 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_496
timestamp 1669390400
transform 1 0 56896 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_499
timestamp 1669390400
transform 1 0 57232 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_508
timestamp 1669390400
transform 1 0 58240 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_512
timestamp 1669390400
transform 1 0 58688 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_2
timestamp 1669390400
transform 1 0 1568 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_5
timestamp 1669390400
transform 1 0 1904 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_25
timestamp 1669390400
transform 1 0 4144 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_34
timestamp 1669390400
transform 1 0 5152 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_37
timestamp 1669390400
transform 1 0 5488 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_39
timestamp 1669390400
transform 1 0 5712 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_55
timestamp 1669390400
transform 1 0 7504 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_67
timestamp 1669390400
transform 1 0 8848 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_79
timestamp 1669390400
transform 1 0 10192 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_83
timestamp 1669390400
transform 1 0 10640 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_97
timestamp 1669390400
transform 1 0 12208 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_101
timestamp 1669390400
transform 1 0 12656 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_105
timestamp 1669390400
transform 1 0 13104 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_108
timestamp 1669390400
transform 1 0 13440 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_111
timestamp 1669390400
transform 1 0 13776 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_131
timestamp 1669390400
transform 1 0 16016 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_143
timestamp 1669390400
transform 1 0 17360 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_154
timestamp 1669390400
transform 1 0 18592 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_168
timestamp 1669390400
transform 1 0 20160 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_172
timestamp 1669390400
transform 1 0 20608 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_176
timestamp 1669390400
transform 1 0 21056 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_179
timestamp 1669390400
transform 1 0 21392 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_182
timestamp 1669390400
transform 1 0 21728 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_186
timestamp 1669390400
transform 1 0 22176 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_206
timestamp 1669390400
transform 1 0 24416 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_222
timestamp 1669390400
transform 1 0 26208 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_228
timestamp 1669390400
transform 1 0 26880 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_247
timestamp 1669390400
transform 1 0 29008 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_250
timestamp 1669390400
transform 1 0 29344 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_253
timestamp 1669390400
transform 1 0 29680 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_302
timestamp 1669390400
transform 1 0 35168 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_314
timestamp 1669390400
transform 1 0 36512 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_318
timestamp 1669390400
transform 1 0 36960 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_321
timestamp 1669390400
transform 1 0 37296 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_328
timestamp 1669390400
transform 1 0 38080 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_330
timestamp 1669390400
transform 1 0 38304 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_354
timestamp 1669390400
transform 1 0 40992 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_358
timestamp 1669390400
transform 1 0 41440 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_362
timestamp 1669390400
transform 1 0 41888 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_366
timestamp 1669390400
transform 1 0 42336 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_370
timestamp 1669390400
transform 1 0 42784 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_374
timestamp 1669390400
transform 1 0 43232 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_378
timestamp 1669390400
transform 1 0 43680 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_382
timestamp 1669390400
transform 1 0 44128 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_392
timestamp 1669390400
transform 1 0 45248 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_396
timestamp 1669390400
transform 1 0 45696 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_400
timestamp 1669390400
transform 1 0 46144 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_404
timestamp 1669390400
transform 1 0 46592 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_414
timestamp 1669390400
transform 1 0 47712 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_422
timestamp 1669390400
transform 1 0 48608 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_426
timestamp 1669390400
transform 1 0 49056 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_429
timestamp 1669390400
transform 1 0 49392 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_443
timestamp 1669390400
transform 1 0 50960 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_447
timestamp 1669390400
transform 1 0 51408 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_455
timestamp 1669390400
transform 1 0 52304 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_457
timestamp 1669390400
transform 1 0 52528 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_460
timestamp 1669390400
transform 1 0 52864 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_463
timestamp 1669390400
transform 1 0 53200 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_472
timestamp 1669390400
transform 1 0 54208 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_476
timestamp 1669390400
transform 1 0 54656 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_480
timestamp 1669390400
transform 1 0 55104 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_490
timestamp 1669390400
transform 1 0 56224 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_494
timestamp 1669390400
transform 1 0 56672 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_509
timestamp 1669390400
transform 1 0 58352 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_2
timestamp 1669390400
transform 1 0 1568 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_6
timestamp 1669390400
transform 1 0 2016 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_10
timestamp 1669390400
transform 1 0 2464 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_14
timestamp 1669390400
transform 1 0 2912 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_43
timestamp 1669390400
transform 1 0 6160 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_58
timestamp 1669390400
transform 1 0 7840 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_70
timestamp 1669390400
transform 1 0 9184 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_73
timestamp 1669390400
transform 1 0 9520 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_82
timestamp 1669390400
transform 1 0 10528 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_92
timestamp 1669390400
transform 1 0 11648 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_98
timestamp 1669390400
transform 1 0 12320 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_102
timestamp 1669390400
transform 1 0 12768 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_106
timestamp 1669390400
transform 1 0 13216 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_118
timestamp 1669390400
transform 1 0 14560 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_130
timestamp 1669390400
transform 1 0 15904 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_134
timestamp 1669390400
transform 1 0 16352 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_137
timestamp 1669390400
transform 1 0 16688 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_141
timestamp 1669390400
transform 1 0 17136 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_144
timestamp 1669390400
transform 1 0 17472 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_146
timestamp 1669390400
transform 1 0 17696 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_149
timestamp 1669390400
transform 1 0 18032 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_153
timestamp 1669390400
transform 1 0 18480 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_157
timestamp 1669390400
transform 1 0 18928 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_176
timestamp 1669390400
transform 1 0 21056 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_185
timestamp 1669390400
transform 1 0 22064 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_189
timestamp 1669390400
transform 1 0 22512 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_192
timestamp 1669390400
transform 1 0 22848 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_196
timestamp 1669390400
transform 1 0 23296 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_200
timestamp 1669390400
transform 1 0 23744 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_204
timestamp 1669390400
transform 1 0 24192 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_208
timestamp 1669390400
transform 1 0 24640 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_212
timestamp 1669390400
transform 1 0 25088 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_215
timestamp 1669390400
transform 1 0 25424 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_226
timestamp 1669390400
transform 1 0 26656 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_230
timestamp 1669390400
transform 1 0 27104 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_257
timestamp 1669390400
transform 1 0 30128 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_267
timestamp 1669390400
transform 1 0 31248 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_271
timestamp 1669390400
transform 1 0 31696 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_274
timestamp 1669390400
transform 1 0 32032 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_283
timestamp 1669390400
transform 1 0 33040 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_286
timestamp 1669390400
transform 1 0 33376 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_312
timestamp 1669390400
transform 1 0 36288 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_326
timestamp 1669390400
transform 1 0 37856 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_330
timestamp 1669390400
transform 1 0 38304 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_340
timestamp 1669390400
transform 1 0 39424 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_348
timestamp 1669390400
transform 1 0 40320 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_352
timestamp 1669390400
transform 1 0 40768 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_354
timestamp 1669390400
transform 1 0 40992 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_357
timestamp 1669390400
transform 1 0 41328 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_371
timestamp 1669390400
transform 1 0 42896 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_381
timestamp 1669390400
transform 1 0 44016 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_385
timestamp 1669390400
transform 1 0 44464 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_389
timestamp 1669390400
transform 1 0 44912 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_391
timestamp 1669390400
transform 1 0 45136 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_405
timestamp 1669390400
transform 1 0 46704 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_411
timestamp 1669390400
transform 1 0 47376 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_415
timestamp 1669390400
transform 1 0 47824 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_425
timestamp 1669390400
transform 1 0 48944 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_428
timestamp 1669390400
transform 1 0 49280 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_435
timestamp 1669390400
transform 1 0 50064 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_437
timestamp 1669390400
transform 1 0 50288 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_450
timestamp 1669390400
transform 1 0 51744 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_454
timestamp 1669390400
transform 1 0 52192 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_460
timestamp 1669390400
transform 1 0 52864 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_464
timestamp 1669390400
transform 1 0 53312 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_472
timestamp 1669390400
transform 1 0 54208 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_478
timestamp 1669390400
transform 1 0 54880 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_482
timestamp 1669390400
transform 1 0 55328 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_492
timestamp 1669390400
transform 1 0 56448 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_496
timestamp 1669390400
transform 1 0 56896 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_499
timestamp 1669390400
transform 1 0 57232 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_508
timestamp 1669390400
transform 1 0 58240 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_512
timestamp 1669390400
transform 1 0 58688 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_2
timestamp 1669390400
transform 1 0 1568 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_6
timestamp 1669390400
transform 1 0 2016 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_10
timestamp 1669390400
transform 1 0 2464 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_14
timestamp 1669390400
transform 1 0 2912 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_24
timestamp 1669390400
transform 1 0 4032 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_30
timestamp 1669390400
transform 1 0 4704 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1669390400
transform 1 0 5152 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_37
timestamp 1669390400
transform 1 0 5488 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_41
timestamp 1669390400
transform 1 0 5936 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_53
timestamp 1669390400
transform 1 0 7280 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_63
timestamp 1669390400
transform 1 0 8400 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_67
timestamp 1669390400
transform 1 0 8848 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_93
timestamp 1669390400
transform 1 0 11760 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_97
timestamp 1669390400
transform 1 0 12208 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_101
timestamp 1669390400
transform 1 0 12656 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_105
timestamp 1669390400
transform 1 0 13104 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_108
timestamp 1669390400
transform 1 0 13440 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_116
timestamp 1669390400
transform 1 0 14336 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_120
timestamp 1669390400
transform 1 0 14784 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_133
timestamp 1669390400
transform 1 0 16240 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_137
timestamp 1669390400
transform 1 0 16688 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_140
timestamp 1669390400
transform 1 0 17024 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_144
timestamp 1669390400
transform 1 0 17472 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_148
timestamp 1669390400
transform 1 0 17920 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_152
timestamp 1669390400
transform 1 0 18368 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_156
timestamp 1669390400
transform 1 0 18816 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_160
timestamp 1669390400
transform 1 0 19264 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_164
timestamp 1669390400
transform 1 0 19712 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_174
timestamp 1669390400
transform 1 0 20832 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_176
timestamp 1669390400
transform 1 0 21056 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_179
timestamp 1669390400
transform 1 0 21392 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_189
timestamp 1669390400
transform 1 0 22512 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_191
timestamp 1669390400
transform 1 0 22736 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_194
timestamp 1669390400
transform 1 0 23072 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_208
timestamp 1669390400
transform 1 0 24640 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_210
timestamp 1669390400
transform 1 0 24864 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_213
timestamp 1669390400
transform 1 0 25200 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_217
timestamp 1669390400
transform 1 0 25648 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_234
timestamp 1669390400
transform 1 0 27552 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_236
timestamp 1669390400
transform 1 0 27776 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_239
timestamp 1669390400
transform 1 0 28112 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_243
timestamp 1669390400
transform 1 0 28560 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_247
timestamp 1669390400
transform 1 0 29008 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_250
timestamp 1669390400
transform 1 0 29344 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_260
timestamp 1669390400
transform 1 0 30464 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_264
timestamp 1669390400
transform 1 0 30912 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_268
timestamp 1669390400
transform 1 0 31360 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_276
timestamp 1669390400
transform 1 0 32256 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_318
timestamp 1669390400
transform 1 0 36960 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_321
timestamp 1669390400
transform 1 0 37296 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_327
timestamp 1669390400
transform 1 0 37968 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_367
timestamp 1669390400
transform 1 0 42448 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_374
timestamp 1669390400
transform 1 0 43232 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_389
timestamp 1669390400
transform 1 0 44912 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_392
timestamp 1669390400
transform 1 0 45248 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_401
timestamp 1669390400
transform 1 0 46256 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_405
timestamp 1669390400
transform 1 0 46704 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_407
timestamp 1669390400
transform 1 0 46928 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_410
timestamp 1669390400
transform 1 0 47264 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_414
timestamp 1669390400
transform 1 0 47712 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_428
timestamp 1669390400
transform 1 0 49280 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_442
timestamp 1669390400
transform 1 0 50848 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_446
timestamp 1669390400
transform 1 0 51296 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_460
timestamp 1669390400
transform 1 0 52864 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_463
timestamp 1669390400
transform 1 0 53200 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_472
timestamp 1669390400
transform 1 0 54208 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_476
timestamp 1669390400
transform 1 0 54656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_488
timestamp 1669390400
transform 1 0 56000 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_496
timestamp 1669390400
transform 1 0 56896 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_510
timestamp 1669390400
transform 1 0 58464 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_512
timestamp 1669390400
transform 1 0 58688 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_2
timestamp 1669390400
transform 1 0 1568 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_6
timestamp 1669390400
transform 1 0 2016 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_16
timestamp 1669390400
transform 1 0 3136 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_20
timestamp 1669390400
transform 1 0 3584 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_35
timestamp 1669390400
transform 1 0 5264 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_39
timestamp 1669390400
transform 1 0 5712 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_46
timestamp 1669390400
transform 1 0 6496 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_58
timestamp 1669390400
transform 1 0 7840 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_62
timestamp 1669390400
transform 1 0 8288 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_66
timestamp 1669390400
transform 1 0 8736 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_70
timestamp 1669390400
transform 1 0 9184 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_73
timestamp 1669390400
transform 1 0 9520 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_89
timestamp 1669390400
transform 1 0 11312 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_104
timestamp 1669390400
transform 1 0 12992 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_106
timestamp 1669390400
transform 1 0 13216 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_112
timestamp 1669390400
transform 1 0 13888 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_122
timestamp 1669390400
transform 1 0 15008 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_124
timestamp 1669390400
transform 1 0 15232 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_127
timestamp 1669390400
transform 1 0 15568 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_131
timestamp 1669390400
transform 1 0 16016 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_141
timestamp 1669390400
transform 1 0 17136 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_144
timestamp 1669390400
transform 1 0 17472 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_157
timestamp 1669390400
transform 1 0 18928 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_163
timestamp 1669390400
transform 1 0 19600 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_188
timestamp 1669390400
transform 1 0 22400 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_199
timestamp 1669390400
transform 1 0 23632 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_201
timestamp 1669390400
transform 1 0 23856 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_212
timestamp 1669390400
transform 1 0 25088 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_215
timestamp 1669390400
transform 1 0 25424 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_231
timestamp 1669390400
transform 1 0 27216 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_241
timestamp 1669390400
transform 1 0 28336 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_267
timestamp 1669390400
transform 1 0 31248 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_274
timestamp 1669390400
transform 1 0 32032 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_278
timestamp 1669390400
transform 1 0 32480 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_282
timestamp 1669390400
transform 1 0 32928 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_286
timestamp 1669390400
transform 1 0 33376 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_289
timestamp 1669390400
transform 1 0 33712 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_293
timestamp 1669390400
transform 1 0 34160 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_299
timestamp 1669390400
transform 1 0 34832 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_316
timestamp 1669390400
transform 1 0 36736 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_320
timestamp 1669390400
transform 1 0 37184 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_324
timestamp 1669390400
transform 1 0 37632 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_333
timestamp 1669390400
transform 1 0 38640 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_340
timestamp 1669390400
transform 1 0 39424 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_354
timestamp 1669390400
transform 1 0 40992 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_357
timestamp 1669390400
transform 1 0 41328 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_365
timestamp 1669390400
transform 1 0 42224 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_379
timestamp 1669390400
transform 1 0 43792 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_383
timestamp 1669390400
transform 1 0 44240 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_392
timestamp 1669390400
transform 1 0 45248 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_396
timestamp 1669390400
transform 1 0 45696 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_412
timestamp 1669390400
transform 1 0 47488 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_420
timestamp 1669390400
transform 1 0 48384 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_424
timestamp 1669390400
transform 1 0 48832 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_428
timestamp 1669390400
transform 1 0 49280 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_432
timestamp 1669390400
transform 1 0 49728 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_435
timestamp 1669390400
transform 1 0 50064 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_445
timestamp 1669390400
transform 1 0 51184 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_449
timestamp 1669390400
transform 1 0 51632 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_457
timestamp 1669390400
transform 1 0 52528 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_461
timestamp 1669390400
transform 1 0 52976 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_463
timestamp 1669390400
transform 1 0 53200 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_476
timestamp 1669390400
transform 1 0 54656 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_490
timestamp 1669390400
transform 1 0 56224 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_494
timestamp 1669390400
transform 1 0 56672 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_496
timestamp 1669390400
transform 1 0 56896 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_499
timestamp 1669390400
transform 1 0 57232 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_506
timestamp 1669390400
transform 1 0 58016 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_510
timestamp 1669390400
transform 1 0 58464 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_512
timestamp 1669390400
transform 1 0 58688 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_2
timestamp 1669390400
transform 1 0 1568 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_4
timestamp 1669390400
transform 1 0 1792 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_15
timestamp 1669390400
transform 1 0 3024 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_31
timestamp 1669390400
transform 1 0 4816 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_37
timestamp 1669390400
transform 1 0 5488 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_53
timestamp 1669390400
transform 1 0 7280 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_55
timestamp 1669390400
transform 1 0 7504 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_66
timestamp 1669390400
transform 1 0 8736 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_72
timestamp 1669390400
transform 1 0 9408 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_79
timestamp 1669390400
transform 1 0 10192 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_95
timestamp 1669390400
transform 1 0 11984 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_101
timestamp 1669390400
transform 1 0 12656 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_105
timestamp 1669390400
transform 1 0 13104 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_108
timestamp 1669390400
transform 1 0 13440 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_124
timestamp 1669390400
transform 1 0 15232 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_138
timestamp 1669390400
transform 1 0 16800 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_150
timestamp 1669390400
transform 1 0 18144 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_160
timestamp 1669390400
transform 1 0 19264 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_168
timestamp 1669390400
transform 1 0 20160 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_172
timestamp 1669390400
transform 1 0 20608 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_176
timestamp 1669390400
transform 1 0 21056 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_179
timestamp 1669390400
transform 1 0 21392 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_190
timestamp 1669390400
transform 1 0 22624 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_197
timestamp 1669390400
transform 1 0 23408 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_201
timestamp 1669390400
transform 1 0 23856 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_220
timestamp 1669390400
transform 1 0 25984 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_224
timestamp 1669390400
transform 1 0 26432 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_228
timestamp 1669390400
transform 1 0 26880 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_245
timestamp 1669390400
transform 1 0 28784 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_247
timestamp 1669390400
transform 1 0 29008 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_250
timestamp 1669390400
transform 1 0 29344 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_252
timestamp 1669390400
transform 1 0 29568 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_255
timestamp 1669390400
transform 1 0 29904 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_280
timestamp 1669390400
transform 1 0 32704 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_284
timestamp 1669390400
transform 1 0 33152 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_288
timestamp 1669390400
transform 1 0 33600 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_292
timestamp 1669390400
transform 1 0 34048 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_296
timestamp 1669390400
transform 1 0 34496 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_300
timestamp 1669390400
transform 1 0 34944 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_304
timestamp 1669390400
transform 1 0 35392 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_316
timestamp 1669390400
transform 1 0 36736 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_318
timestamp 1669390400
transform 1 0 36960 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_321
timestamp 1669390400
transform 1 0 37296 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_324
timestamp 1669390400
transform 1 0 37632 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_328
timestamp 1669390400
transform 1 0 38080 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_339
timestamp 1669390400
transform 1 0 39312 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_343
timestamp 1669390400
transform 1 0 39760 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_350
timestamp 1669390400
transform 1 0 40544 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_357
timestamp 1669390400
transform 1 0 41328 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_361
timestamp 1669390400
transform 1 0 41776 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_365
timestamp 1669390400
transform 1 0 42224 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_369
timestamp 1669390400
transform 1 0 42672 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_373
timestamp 1669390400
transform 1 0 43120 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_377
timestamp 1669390400
transform 1 0 43568 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_381
timestamp 1669390400
transform 1 0 44016 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_385
timestamp 1669390400
transform 1 0 44464 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_389
timestamp 1669390400
transform 1 0 44912 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_392
timestamp 1669390400
transform 1 0 45248 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_396
timestamp 1669390400
transform 1 0 45696 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_400
timestamp 1669390400
transform 1 0 46144 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_406
timestamp 1669390400
transform 1 0 46816 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_410
timestamp 1669390400
transform 1 0 47264 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_418
timestamp 1669390400
transform 1 0 48160 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_422
timestamp 1669390400
transform 1 0 48608 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_424
timestamp 1669390400
transform 1 0 48832 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_427
timestamp 1669390400
transform 1 0 49168 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_431
timestamp 1669390400
transform 1 0 49616 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_447
timestamp 1669390400
transform 1 0 51408 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_455
timestamp 1669390400
transform 1 0 52304 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_459
timestamp 1669390400
transform 1 0 52752 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_463
timestamp 1669390400
transform 1 0 53200 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_471
timestamp 1669390400
transform 1 0 54096 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_475
timestamp 1669390400
transform 1 0 54544 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_478
timestamp 1669390400
transform 1 0 54880 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_498
timestamp 1669390400
transform 1 0 57120 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_508
timestamp 1669390400
transform 1 0 58240 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_512
timestamp 1669390400
transform 1 0 58688 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_2
timestamp 1669390400
transform 1 0 1568 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_4
timestamp 1669390400
transform 1 0 1792 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_7
timestamp 1669390400
transform 1 0 2128 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_11
timestamp 1669390400
transform 1 0 2576 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_21
timestamp 1669390400
transform 1 0 3696 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_31
timestamp 1669390400
transform 1 0 4816 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_39
timestamp 1669390400
transform 1 0 5712 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_43
timestamp 1669390400
transform 1 0 6160 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_47
timestamp 1669390400
transform 1 0 6608 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_62
timestamp 1669390400
transform 1 0 8288 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_66
timestamp 1669390400
transform 1 0 8736 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_70
timestamp 1669390400
transform 1 0 9184 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_73
timestamp 1669390400
transform 1 0 9520 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_89
timestamp 1669390400
transform 1 0 11312 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_95
timestamp 1669390400
transform 1 0 11984 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_99
timestamp 1669390400
transform 1 0 12432 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_124
timestamp 1669390400
transform 1 0 15232 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_135
timestamp 1669390400
transform 1 0 16464 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_141
timestamp 1669390400
transform 1 0 17136 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_144
timestamp 1669390400
transform 1 0 17472 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_150
timestamp 1669390400
transform 1 0 18144 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_154
timestamp 1669390400
transform 1 0 18592 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_157
timestamp 1669390400
transform 1 0 18928 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_161
timestamp 1669390400
transform 1 0 19376 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_163
timestamp 1669390400
transform 1 0 19600 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_166
timestamp 1669390400
transform 1 0 19936 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_170
timestamp 1669390400
transform 1 0 20384 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_174
timestamp 1669390400
transform 1 0 20832 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_184
timestamp 1669390400
transform 1 0 21952 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_188
timestamp 1669390400
transform 1 0 22400 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_192
timestamp 1669390400
transform 1 0 22848 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_196
timestamp 1669390400
transform 1 0 23296 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_200
timestamp 1669390400
transform 1 0 23744 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_204
timestamp 1669390400
transform 1 0 24192 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_208
timestamp 1669390400
transform 1 0 24640 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_212
timestamp 1669390400
transform 1 0 25088 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_215
timestamp 1669390400
transform 1 0 25424 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_218
timestamp 1669390400
transform 1 0 25760 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_222
timestamp 1669390400
transform 1 0 26208 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_226
timestamp 1669390400
transform 1 0 26656 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_240
timestamp 1669390400
transform 1 0 28224 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_252
timestamp 1669390400
transform 1 0 29568 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_256
timestamp 1669390400
transform 1 0 30016 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_264
timestamp 1669390400
transform 1 0 30912 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_266
timestamp 1669390400
transform 1 0 31136 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_281
timestamp 1669390400
transform 1 0 32816 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_283
timestamp 1669390400
transform 1 0 33040 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_286
timestamp 1669390400
transform 1 0 33376 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_289
timestamp 1669390400
transform 1 0 33712 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_305
timestamp 1669390400
transform 1 0 35504 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_309
timestamp 1669390400
transform 1 0 35952 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_313
timestamp 1669390400
transform 1 0 36400 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_317
timestamp 1669390400
transform 1 0 36848 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_321
timestamp 1669390400
transform 1 0 37296 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_325
timestamp 1669390400
transform 1 0 37744 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_350
timestamp 1669390400
transform 1 0 40544 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_354
timestamp 1669390400
transform 1 0 40992 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_357
timestamp 1669390400
transform 1 0 41328 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_360
timestamp 1669390400
transform 1 0 41664 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_387
timestamp 1669390400
transform 1 0 44688 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_391
timestamp 1669390400
transform 1 0 45136 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_395
timestamp 1669390400
transform 1 0 45584 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_409
timestamp 1669390400
transform 1 0 47152 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_423
timestamp 1669390400
transform 1 0 48720 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_425
timestamp 1669390400
transform 1 0 48944 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_428
timestamp 1669390400
transform 1 0 49280 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_441
timestamp 1669390400
transform 1 0 50736 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_443
timestamp 1669390400
transform 1 0 50960 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_446
timestamp 1669390400
transform 1 0 51296 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_450
timestamp 1669390400
transform 1 0 51744 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_456
timestamp 1669390400
transform 1 0 52416 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_460
timestamp 1669390400
transform 1 0 52864 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_472
timestamp 1669390400
transform 1 0 54208 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_480
timestamp 1669390400
transform 1 0 55104 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_484
timestamp 1669390400
transform 1 0 55552 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_494
timestamp 1669390400
transform 1 0 56672 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_496
timestamp 1669390400
transform 1 0 56896 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_499
timestamp 1669390400
transform 1 0 57232 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_512
timestamp 1669390400
transform 1 0 58688 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_2
timestamp 1669390400
transform 1 0 1568 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_5
timestamp 1669390400
transform 1 0 1904 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_15
timestamp 1669390400
transform 1 0 3024 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_29
timestamp 1669390400
transform 1 0 4592 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_31
timestamp 1669390400
transform 1 0 4816 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_34
timestamp 1669390400
transform 1 0 5152 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_37
timestamp 1669390400
transform 1 0 5488 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_45
timestamp 1669390400
transform 1 0 6384 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_56
timestamp 1669390400
transform 1 0 7616 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_68
timestamp 1669390400
transform 1 0 8960 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_72
timestamp 1669390400
transform 1 0 9408 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_75
timestamp 1669390400
transform 1 0 9744 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_90
timestamp 1669390400
transform 1 0 11424 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_92
timestamp 1669390400
transform 1 0 11648 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_103
timestamp 1669390400
transform 1 0 12880 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1669390400
transform 1 0 13104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_108
timestamp 1669390400
transform 1 0 13440 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_119
timestamp 1669390400
transform 1 0 14672 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_121
timestamp 1669390400
transform 1 0 14896 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_124
timestamp 1669390400
transform 1 0 15232 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_128
timestamp 1669390400
transform 1 0 15680 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_132
timestamp 1669390400
transform 1 0 16128 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_140
timestamp 1669390400
transform 1 0 17024 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_146
timestamp 1669390400
transform 1 0 17696 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_150
timestamp 1669390400
transform 1 0 18144 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_154
timestamp 1669390400
transform 1 0 18592 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_164
timestamp 1669390400
transform 1 0 19712 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_176
timestamp 1669390400
transform 1 0 21056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_179
timestamp 1669390400
transform 1 0 21392 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_182
timestamp 1669390400
transform 1 0 21728 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_186
timestamp 1669390400
transform 1 0 22176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_192
timestamp 1669390400
transform 1 0 22848 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_196
timestamp 1669390400
transform 1 0 23296 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_200
timestamp 1669390400
transform 1 0 23744 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_220
timestamp 1669390400
transform 1 0 25984 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_222
timestamp 1669390400
transform 1 0 26208 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_225
timestamp 1669390400
transform 1 0 26544 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_235
timestamp 1669390400
transform 1 0 27664 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_245
timestamp 1669390400
transform 1 0 28784 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_247
timestamp 1669390400
transform 1 0 29008 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_250
timestamp 1669390400
transform 1 0 29344 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_260
timestamp 1669390400
transform 1 0 30464 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_272
timestamp 1669390400
transform 1 0 31808 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_282
timestamp 1669390400
transform 1 0 32928 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_289
timestamp 1669390400
transform 1 0 33712 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_306
timestamp 1669390400
transform 1 0 35616 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_313
timestamp 1669390400
transform 1 0 36400 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_317
timestamp 1669390400
transform 1 0 36848 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_321
timestamp 1669390400
transform 1 0 37296 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_330
timestamp 1669390400
transform 1 0 38304 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_338
timestamp 1669390400
transform 1 0 39200 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_342
timestamp 1669390400
transform 1 0 39648 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_346
timestamp 1669390400
transform 1 0 40096 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_350
timestamp 1669390400
transform 1 0 40544 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_354
timestamp 1669390400
transform 1 0 40992 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_358
timestamp 1669390400
transform 1 0 41440 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_365
timestamp 1669390400
transform 1 0 42224 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_375
timestamp 1669390400
transform 1 0 43344 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_382
timestamp 1669390400
transform 1 0 44128 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_386
timestamp 1669390400
transform 1 0 44576 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_392
timestamp 1669390400
transform 1 0 45248 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_405
timestamp 1669390400
transform 1 0 46704 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_415
timestamp 1669390400
transform 1 0 47824 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_417
timestamp 1669390400
transform 1 0 48048 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_441
timestamp 1669390400
transform 1 0 50736 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_445
timestamp 1669390400
transform 1 0 51184 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_459
timestamp 1669390400
transform 1 0 52752 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_463
timestamp 1669390400
transform 1 0 53200 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_476
timestamp 1669390400
transform 1 0 54656 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_484
timestamp 1669390400
transform 1 0 55552 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_488
timestamp 1669390400
transform 1 0 56000 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_502
timestamp 1669390400
transform 1 0 57568 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_510
timestamp 1669390400
transform 1 0 58464 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_512
timestamp 1669390400
transform 1 0 58688 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_2
timestamp 1669390400
transform 1 0 1568 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_8
timestamp 1669390400
transform 1 0 2240 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_12
timestamp 1669390400
transform 1 0 2688 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_33
timestamp 1669390400
transform 1 0 5040 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_40
timestamp 1669390400
transform 1 0 5824 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_50
timestamp 1669390400
transform 1 0 6944 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_54
timestamp 1669390400
transform 1 0 7392 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_58
timestamp 1669390400
transform 1 0 7840 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_62
timestamp 1669390400
transform 1 0 8288 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_66
timestamp 1669390400
transform 1 0 8736 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_70
timestamp 1669390400
transform 1 0 9184 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_73
timestamp 1669390400
transform 1 0 9520 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_89
timestamp 1669390400
transform 1 0 11312 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_101
timestamp 1669390400
transform 1 0 12656 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_103
timestamp 1669390400
transform 1 0 12880 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_106
timestamp 1669390400
transform 1 0 13216 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_113
timestamp 1669390400
transform 1 0 14000 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_117
timestamp 1669390400
transform 1 0 14448 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_128
timestamp 1669390400
transform 1 0 15680 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_141
timestamp 1669390400
transform 1 0 17136 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_144
timestamp 1669390400
transform 1 0 17472 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_156
timestamp 1669390400
transform 1 0 18816 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_160
timestamp 1669390400
transform 1 0 19264 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_163
timestamp 1669390400
transform 1 0 19600 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_173
timestamp 1669390400
transform 1 0 20720 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_183
timestamp 1669390400
transform 1 0 21840 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_185
timestamp 1669390400
transform 1 0 22064 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_188
timestamp 1669390400
transform 1 0 22400 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_192
timestamp 1669390400
transform 1 0 22848 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_212
timestamp 1669390400
transform 1 0 25088 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_215
timestamp 1669390400
transform 1 0 25424 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_225
timestamp 1669390400
transform 1 0 26544 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_229
timestamp 1669390400
transform 1 0 26992 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_249
timestamp 1669390400
transform 1 0 29232 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_266
timestamp 1669390400
transform 1 0 31136 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_276
timestamp 1669390400
transform 1 0 32256 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_280
timestamp 1669390400
transform 1 0 32704 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_286
timestamp 1669390400
transform 1 0 33376 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_293
timestamp 1669390400
transform 1 0 34160 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_295
timestamp 1669390400
transform 1 0 34384 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_305
timestamp 1669390400
transform 1 0 35504 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_309
timestamp 1669390400
transform 1 0 35952 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_313
timestamp 1669390400
transform 1 0 36400 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_315
timestamp 1669390400
transform 1 0 36624 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_326
timestamp 1669390400
transform 1 0 37856 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_330
timestamp 1669390400
transform 1 0 38304 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_334
timestamp 1669390400
transform 1 0 38752 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_338
timestamp 1669390400
transform 1 0 39200 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_346
timestamp 1669390400
transform 1 0 40096 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_354
timestamp 1669390400
transform 1 0 40992 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_357
timestamp 1669390400
transform 1 0 41328 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_370
timestamp 1669390400
transform 1 0 42784 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_374
timestamp 1669390400
transform 1 0 43232 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_378
timestamp 1669390400
transform 1 0 43680 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_382
timestamp 1669390400
transform 1 0 44128 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_386
timestamp 1669390400
transform 1 0 44576 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_390
timestamp 1669390400
transform 1 0 45024 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_398
timestamp 1669390400
transform 1 0 45920 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_402
timestamp 1669390400
transform 1 0 46368 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_406
timestamp 1669390400
transform 1 0 46816 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_416
timestamp 1669390400
transform 1 0 47936 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_420
timestamp 1669390400
transform 1 0 48384 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_424
timestamp 1669390400
transform 1 0 48832 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_428
timestamp 1669390400
transform 1 0 49280 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_435
timestamp 1669390400
transform 1 0 50064 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_437
timestamp 1669390400
transform 1 0 50288 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_450
timestamp 1669390400
transform 1 0 51744 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_454
timestamp 1669390400
transform 1 0 52192 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_458
timestamp 1669390400
transform 1 0 52640 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_471
timestamp 1669390400
transform 1 0 54096 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_486
timestamp 1669390400
transform 1 0 55776 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_496
timestamp 1669390400
transform 1 0 56896 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_499
timestamp 1669390400
transform 1 0 57232 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_508
timestamp 1669390400
transform 1 0 58240 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_512
timestamp 1669390400
transform 1 0 58688 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_2
timestamp 1669390400
transform 1 0 1568 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_5
timestamp 1669390400
transform 1 0 1904 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_9
timestamp 1669390400
transform 1 0 2352 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_34
timestamp 1669390400
transform 1 0 5152 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_37
timestamp 1669390400
transform 1 0 5488 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_49
timestamp 1669390400
transform 1 0 6832 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_61
timestamp 1669390400
transform 1 0 8176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_65
timestamp 1669390400
transform 1 0 8624 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_74
timestamp 1669390400
transform 1 0 9632 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_88
timestamp 1669390400
transform 1 0 11200 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_98
timestamp 1669390400
transform 1 0 12320 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_102
timestamp 1669390400
transform 1 0 12768 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_105
timestamp 1669390400
transform 1 0 13104 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_108
timestamp 1669390400
transform 1 0 13440 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_132
timestamp 1669390400
transform 1 0 16128 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_134
timestamp 1669390400
transform 1 0 16352 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_140
timestamp 1669390400
transform 1 0 17024 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_154
timestamp 1669390400
transform 1 0 18592 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_164
timestamp 1669390400
transform 1 0 19712 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_168
timestamp 1669390400
transform 1 0 20160 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_172
timestamp 1669390400
transform 1 0 20608 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_176
timestamp 1669390400
transform 1 0 21056 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_179
timestamp 1669390400
transform 1 0 21392 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_188
timestamp 1669390400
transform 1 0 22400 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_195
timestamp 1669390400
transform 1 0 23184 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_197
timestamp 1669390400
transform 1 0 23408 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_200
timestamp 1669390400
transform 1 0 23744 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_204
timestamp 1669390400
transform 1 0 24192 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_208
timestamp 1669390400
transform 1 0 24640 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_215
timestamp 1669390400
transform 1 0 25424 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_227
timestamp 1669390400
transform 1 0 26768 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_247
timestamp 1669390400
transform 1 0 29008 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_250
timestamp 1669390400
transform 1 0 29344 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_259
timestamp 1669390400
transform 1 0 30352 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_263
timestamp 1669390400
transform 1 0 30800 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_266
timestamp 1669390400
transform 1 0 31136 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_276
timestamp 1669390400
transform 1 0 32256 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_280
timestamp 1669390400
transform 1 0 32704 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_284
timestamp 1669390400
transform 1 0 33152 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_294
timestamp 1669390400
transform 1 0 34272 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_298
timestamp 1669390400
transform 1 0 34720 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_302
timestamp 1669390400
transform 1 0 35168 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_311
timestamp 1669390400
transform 1 0 36176 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_315
timestamp 1669390400
transform 1 0 36624 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_321
timestamp 1669390400
transform 1 0 37296 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_324
timestamp 1669390400
transform 1 0 37632 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_328
timestamp 1669390400
transform 1 0 38080 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_332
timestamp 1669390400
transform 1 0 38528 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_336
timestamp 1669390400
transform 1 0 38976 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_340
timestamp 1669390400
transform 1 0 39424 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_346
timestamp 1669390400
transform 1 0 40096 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_350
timestamp 1669390400
transform 1 0 40544 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_362
timestamp 1669390400
transform 1 0 41888 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_366
timestamp 1669390400
transform 1 0 42336 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_376
timestamp 1669390400
transform 1 0 43456 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_382
timestamp 1669390400
transform 1 0 44128 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_386
timestamp 1669390400
transform 1 0 44576 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_392
timestamp 1669390400
transform 1 0 45248 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_395
timestamp 1669390400
transform 1 0 45584 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_399
timestamp 1669390400
transform 1 0 46032 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_406
timestamp 1669390400
transform 1 0 46816 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_413
timestamp 1669390400
transform 1 0 47600 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_417
timestamp 1669390400
transform 1 0 48048 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_433
timestamp 1669390400
transform 1 0 49840 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_443
timestamp 1669390400
transform 1 0 50960 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_447
timestamp 1669390400
transform 1 0 51408 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_455
timestamp 1669390400
transform 1 0 52304 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_459
timestamp 1669390400
transform 1 0 52752 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_463
timestamp 1669390400
transform 1 0 53200 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_472
timestamp 1669390400
transform 1 0 54208 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_482
timestamp 1669390400
transform 1 0 55328 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_490
timestamp 1669390400
transform 1 0 56224 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_506
timestamp 1669390400
transform 1 0 58016 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_510
timestamp 1669390400
transform 1 0 58464 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_512
timestamp 1669390400
transform 1 0 58688 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_2
timestamp 1669390400
transform 1 0 1568 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_4
timestamp 1669390400
transform 1 0 1792 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_7
timestamp 1669390400
transform 1 0 2128 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_11
timestamp 1669390400
transform 1 0 2576 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_24
timestamp 1669390400
transform 1 0 4032 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_32
timestamp 1669390400
transform 1 0 4928 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_36
timestamp 1669390400
transform 1 0 5376 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_40
timestamp 1669390400
transform 1 0 5824 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_44
timestamp 1669390400
transform 1 0 6272 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_48
timestamp 1669390400
transform 1 0 6720 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_67
timestamp 1669390400
transform 1 0 8848 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_73
timestamp 1669390400
transform 1 0 9520 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_84
timestamp 1669390400
transform 1 0 10752 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_91
timestamp 1669390400
transform 1 0 11536 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_95
timestamp 1669390400
transform 1 0 11984 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_98
timestamp 1669390400
transform 1 0 12320 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_112
timestamp 1669390400
transform 1 0 13888 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_114
timestamp 1669390400
transform 1 0 14112 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_130
timestamp 1669390400
transform 1 0 15904 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_140
timestamp 1669390400
transform 1 0 17024 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_144
timestamp 1669390400
transform 1 0 17472 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_156
timestamp 1669390400
transform 1 0 18816 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_160
timestamp 1669390400
transform 1 0 19264 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_163
timestamp 1669390400
transform 1 0 19600 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_167
timestamp 1669390400
transform 1 0 20048 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_180
timestamp 1669390400
transform 1 0 21504 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_190
timestamp 1669390400
transform 1 0 22624 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_196
timestamp 1669390400
transform 1 0 23296 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_200
timestamp 1669390400
transform 1 0 23744 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_204
timestamp 1669390400
transform 1 0 24192 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_208
timestamp 1669390400
transform 1 0 24640 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_212
timestamp 1669390400
transform 1 0 25088 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_215
timestamp 1669390400
transform 1 0 25424 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_221
timestamp 1669390400
transform 1 0 26096 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_225
timestamp 1669390400
transform 1 0 26544 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_240
timestamp 1669390400
transform 1 0 28224 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_244
timestamp 1669390400
transform 1 0 28672 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_255
timestamp 1669390400
transform 1 0 29904 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_259
timestamp 1669390400
transform 1 0 30352 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_263
timestamp 1669390400
transform 1 0 30800 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_279
timestamp 1669390400
transform 1 0 32592 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_283
timestamp 1669390400
transform 1 0 33040 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_286
timestamp 1669390400
transform 1 0 33376 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_289
timestamp 1669390400
transform 1 0 33712 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_291
timestamp 1669390400
transform 1 0 33936 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_301
timestamp 1669390400
transform 1 0 35056 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_305
timestamp 1669390400
transform 1 0 35504 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_330
timestamp 1669390400
transform 1 0 38304 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_337
timestamp 1669390400
transform 1 0 39088 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_339
timestamp 1669390400
transform 1 0 39312 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_353
timestamp 1669390400
transform 1 0 40880 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_357
timestamp 1669390400
transform 1 0 41328 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_360
timestamp 1669390400
transform 1 0 41664 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_364
timestamp 1669390400
transform 1 0 42112 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_378
timestamp 1669390400
transform 1 0 43680 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_392
timestamp 1669390400
transform 1 0 45248 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_396
timestamp 1669390400
transform 1 0 45696 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_421
timestamp 1669390400
transform 1 0 48496 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_425
timestamp 1669390400
transform 1 0 48944 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_43_428
timestamp 1669390400
transform 1 0 49280 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_460
timestamp 1669390400
transform 1 0 52864 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_468
timestamp 1669390400
transform 1 0 53760 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_472
timestamp 1669390400
transform 1 0 54208 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_475
timestamp 1669390400
transform 1 0 54544 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_479
timestamp 1669390400
transform 1 0 54992 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_487
timestamp 1669390400
transform 1 0 55888 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_489
timestamp 1669390400
transform 1 0 56112 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_492
timestamp 1669390400
transform 1 0 56448 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_496
timestamp 1669390400
transform 1 0 56896 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_499
timestamp 1669390400
transform 1 0 57232 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_506
timestamp 1669390400
transform 1 0 58016 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_510
timestamp 1669390400
transform 1 0 58464 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_512
timestamp 1669390400
transform 1 0 58688 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_2
timestamp 1669390400
transform 1 0 1568 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_6
timestamp 1669390400
transform 1 0 2016 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_10
timestamp 1669390400
transform 1 0 2464 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_20
timestamp 1669390400
transform 1 0 3584 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_30
timestamp 1669390400
transform 1 0 4704 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_34
timestamp 1669390400
transform 1 0 5152 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_37
timestamp 1669390400
transform 1 0 5488 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_61
timestamp 1669390400
transform 1 0 8176 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_73
timestamp 1669390400
transform 1 0 9520 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_77
timestamp 1669390400
transform 1 0 9968 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_81
timestamp 1669390400
transform 1 0 10416 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_85
timestamp 1669390400
transform 1 0 10864 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_89
timestamp 1669390400
transform 1 0 11312 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_93
timestamp 1669390400
transform 1 0 11760 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_97
timestamp 1669390400
transform 1 0 12208 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_101
timestamp 1669390400
transform 1 0 12656 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_105
timestamp 1669390400
transform 1 0 13104 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_108
timestamp 1669390400
transform 1 0 13440 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_127
timestamp 1669390400
transform 1 0 15568 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_135
timestamp 1669390400
transform 1 0 16464 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_139
timestamp 1669390400
transform 1 0 16912 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_143
timestamp 1669390400
transform 1 0 17360 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_147
timestamp 1669390400
transform 1 0 17808 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_151
timestamp 1669390400
transform 1 0 18256 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_155
timestamp 1669390400
transform 1 0 18704 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_159
timestamp 1669390400
transform 1 0 19152 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_176
timestamp 1669390400
transform 1 0 21056 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_179
timestamp 1669390400
transform 1 0 21392 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_199
timestamp 1669390400
transform 1 0 23632 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_219
timestamp 1669390400
transform 1 0 25872 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_233
timestamp 1669390400
transform 1 0 27440 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_240
timestamp 1669390400
transform 1 0 28224 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_244
timestamp 1669390400
transform 1 0 28672 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_247
timestamp 1669390400
transform 1 0 29008 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_250
timestamp 1669390400
transform 1 0 29344 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_253
timestamp 1669390400
transform 1 0 29680 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_257
timestamp 1669390400
transform 1 0 30128 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_277
timestamp 1669390400
transform 1 0 32368 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_281
timestamp 1669390400
transform 1 0 32816 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_283
timestamp 1669390400
transform 1 0 33040 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_289
timestamp 1669390400
transform 1 0 33712 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_299
timestamp 1669390400
transform 1 0 34832 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_309
timestamp 1669390400
transform 1 0 35952 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_313
timestamp 1669390400
transform 1 0 36400 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_317
timestamp 1669390400
transform 1 0 36848 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_321
timestamp 1669390400
transform 1 0 37296 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_324
timestamp 1669390400
transform 1 0 37632 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_338
timestamp 1669390400
transform 1 0 39200 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_340
timestamp 1669390400
transform 1 0 39424 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_349
timestamp 1669390400
transform 1 0 40432 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_353
timestamp 1669390400
transform 1 0 40880 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_357
timestamp 1669390400
transform 1 0 41328 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_361
timestamp 1669390400
transform 1 0 41776 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_365
timestamp 1669390400
transform 1 0 42224 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_373
timestamp 1669390400
transform 1 0 43120 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_385
timestamp 1669390400
transform 1 0 44464 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_389
timestamp 1669390400
transform 1 0 44912 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_392
timestamp 1669390400
transform 1 0 45248 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_394
timestamp 1669390400
transform 1 0 45472 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_397
timestamp 1669390400
transform 1 0 45808 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_401
timestamp 1669390400
transform 1 0 46256 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_411
timestamp 1669390400
transform 1 0 47376 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_427
timestamp 1669390400
transform 1 0 49168 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_431
timestamp 1669390400
transform 1 0 49616 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_446
timestamp 1669390400
transform 1 0 51296 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_453
timestamp 1669390400
transform 1 0 52080 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_463
timestamp 1669390400
transform 1 0 53200 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_472
timestamp 1669390400
transform 1 0 54208 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_476
timestamp 1669390400
transform 1 0 54656 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_496
timestamp 1669390400
transform 1 0 56896 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_511
timestamp 1669390400
transform 1 0 58576 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_2
timestamp 1669390400
transform 1 0 1568 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_4
timestamp 1669390400
transform 1 0 1792 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_13
timestamp 1669390400
transform 1 0 2800 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_25
timestamp 1669390400
transform 1 0 4144 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_27
timestamp 1669390400
transform 1 0 4368 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_36
timestamp 1669390400
transform 1 0 5376 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_40
timestamp 1669390400
transform 1 0 5824 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_50
timestamp 1669390400
transform 1 0 6944 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_63
timestamp 1669390400
transform 1 0 8400 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_67
timestamp 1669390400
transform 1 0 8848 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_70
timestamp 1669390400
transform 1 0 9184 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_73
timestamp 1669390400
transform 1 0 9520 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_77
timestamp 1669390400
transform 1 0 9968 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_87
timestamp 1669390400
transform 1 0 11088 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_91
timestamp 1669390400
transform 1 0 11536 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_104
timestamp 1669390400
transform 1 0 12992 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_108
timestamp 1669390400
transform 1 0 13440 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_112
timestamp 1669390400
transform 1 0 13888 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_122
timestamp 1669390400
transform 1 0 15008 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_129
timestamp 1669390400
transform 1 0 15792 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_133
timestamp 1669390400
transform 1 0 16240 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_141
timestamp 1669390400
transform 1 0 17136 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_144
timestamp 1669390400
transform 1 0 17472 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_153
timestamp 1669390400
transform 1 0 18480 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_157
timestamp 1669390400
transform 1 0 18928 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_168
timestamp 1669390400
transform 1 0 20160 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_187
timestamp 1669390400
transform 1 0 22288 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_189
timestamp 1669390400
transform 1 0 22512 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_192
timestamp 1669390400
transform 1 0 22848 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_196
timestamp 1669390400
transform 1 0 23296 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_200
timestamp 1669390400
transform 1 0 23744 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_204
timestamp 1669390400
transform 1 0 24192 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_208
timestamp 1669390400
transform 1 0 24640 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_212
timestamp 1669390400
transform 1 0 25088 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_215
timestamp 1669390400
transform 1 0 25424 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_238
timestamp 1669390400
transform 1 0 28000 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_242
timestamp 1669390400
transform 1 0 28448 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_245
timestamp 1669390400
transform 1 0 28784 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_260
timestamp 1669390400
transform 1 0 30464 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_264
timestamp 1669390400
transform 1 0 30912 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_276
timestamp 1669390400
transform 1 0 32256 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_278
timestamp 1669390400
transform 1 0 32480 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_281
timestamp 1669390400
transform 1 0 32816 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_283
timestamp 1669390400
transform 1 0 33040 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_286
timestamp 1669390400
transform 1 0 33376 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_295
timestamp 1669390400
transform 1 0 34384 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_313
timestamp 1669390400
transform 1 0 36400 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_317
timestamp 1669390400
transform 1 0 36848 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_321
timestamp 1669390400
transform 1 0 37296 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_325
timestamp 1669390400
transform 1 0 37744 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_333
timestamp 1669390400
transform 1 0 38640 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_337
timestamp 1669390400
transform 1 0 39088 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_340
timestamp 1669390400
transform 1 0 39424 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_354
timestamp 1669390400
transform 1 0 40992 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_357
timestamp 1669390400
transform 1 0 41328 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_361
timestamp 1669390400
transform 1 0 41776 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_365
timestamp 1669390400
transform 1 0 42224 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_369
timestamp 1669390400
transform 1 0 42672 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_373
timestamp 1669390400
transform 1 0 43120 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_391
timestamp 1669390400
transform 1 0 45136 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_395
timestamp 1669390400
transform 1 0 45584 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_399
timestamp 1669390400
transform 1 0 46032 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_403
timestamp 1669390400
transform 1 0 46480 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_407
timestamp 1669390400
transform 1 0 46928 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_411
timestamp 1669390400
transform 1 0 47376 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_425
timestamp 1669390400
transform 1 0 48944 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_428
timestamp 1669390400
transform 1 0 49280 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_441
timestamp 1669390400
transform 1 0 50736 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_456
timestamp 1669390400
transform 1 0 52416 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_460
timestamp 1669390400
transform 1 0 52864 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_486
timestamp 1669390400
transform 1 0 55776 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_496
timestamp 1669390400
transform 1 0 56896 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_499
timestamp 1669390400
transform 1 0 57232 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_512
timestamp 1669390400
transform 1 0 58688 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_2
timestamp 1669390400
transform 1 0 1568 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_4
timestamp 1669390400
transform 1 0 1792 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_7
timestamp 1669390400
transform 1 0 2128 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_17
timestamp 1669390400
transform 1 0 3248 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_19
timestamp 1669390400
transform 1 0 3472 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_22
timestamp 1669390400
transform 1 0 3808 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_26
timestamp 1669390400
transform 1 0 4256 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_30
timestamp 1669390400
transform 1 0 4704 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_34
timestamp 1669390400
transform 1 0 5152 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_37
timestamp 1669390400
transform 1 0 5488 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_40
timestamp 1669390400
transform 1 0 5824 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_47
timestamp 1669390400
transform 1 0 6608 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_51
timestamp 1669390400
transform 1 0 7056 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_60
timestamp 1669390400
transform 1 0 8064 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_64
timestamp 1669390400
transform 1 0 8512 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_68
timestamp 1669390400
transform 1 0 8960 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_72
timestamp 1669390400
transform 1 0 9408 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_86
timestamp 1669390400
transform 1 0 10976 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_88
timestamp 1669390400
transform 1 0 11200 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_97
timestamp 1669390400
transform 1 0 12208 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_101
timestamp 1669390400
transform 1 0 12656 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_105
timestamp 1669390400
transform 1 0 13104 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_108
timestamp 1669390400
transform 1 0 13440 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_111
timestamp 1669390400
transform 1 0 13776 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_115
timestamp 1669390400
transform 1 0 14224 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_127
timestamp 1669390400
transform 1 0 15568 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_131
timestamp 1669390400
transform 1 0 16016 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_134
timestamp 1669390400
transform 1 0 16352 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_148
timestamp 1669390400
transform 1 0 17920 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_159
timestamp 1669390400
transform 1 0 19152 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_169
timestamp 1669390400
transform 1 0 20272 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_173
timestamp 1669390400
transform 1 0 20720 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_176
timestamp 1669390400
transform 1 0 21056 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_179
timestamp 1669390400
transform 1 0 21392 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_188
timestamp 1669390400
transform 1 0 22400 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_194
timestamp 1669390400
transform 1 0 23072 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_214
timestamp 1669390400
transform 1 0 25312 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_216
timestamp 1669390400
transform 1 0 25536 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_219
timestamp 1669390400
transform 1 0 25872 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_223
timestamp 1669390400
transform 1 0 26320 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_247
timestamp 1669390400
transform 1 0 29008 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_250
timestamp 1669390400
transform 1 0 29344 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_305
timestamp 1669390400
transform 1 0 35504 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_315
timestamp 1669390400
transform 1 0 36624 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_321
timestamp 1669390400
transform 1 0 37296 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_329
timestamp 1669390400
transform 1 0 38192 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_331
timestamp 1669390400
transform 1 0 38416 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_334
timestamp 1669390400
transform 1 0 38752 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_342
timestamp 1669390400
transform 1 0 39648 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_346
timestamp 1669390400
transform 1 0 40096 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_348
timestamp 1669390400
transform 1 0 40320 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_351
timestamp 1669390400
transform 1 0 40656 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_365
timestamp 1669390400
transform 1 0 42224 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_375
timestamp 1669390400
transform 1 0 43344 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_389
timestamp 1669390400
transform 1 0 44912 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_392
timestamp 1669390400
transform 1 0 45248 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_401
timestamp 1669390400
transform 1 0 46256 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_405
timestamp 1669390400
transform 1 0 46704 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_425
timestamp 1669390400
transform 1 0 48944 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_438
timestamp 1669390400
transform 1 0 50400 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_448
timestamp 1669390400
transform 1 0 51520 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_456
timestamp 1669390400
transform 1 0 52416 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_460
timestamp 1669390400
transform 1 0 52864 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_463
timestamp 1669390400
transform 1 0 53200 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_471
timestamp 1669390400
transform 1 0 54096 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_478
timestamp 1669390400
transform 1 0 54880 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_486
timestamp 1669390400
transform 1 0 55776 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_490
timestamp 1669390400
transform 1 0 56224 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_492
timestamp 1669390400
transform 1 0 56448 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_495
timestamp 1669390400
transform 1 0 56784 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_510
timestamp 1669390400
transform 1 0 58464 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_512
timestamp 1669390400
transform 1 0 58688 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_2
timestamp 1669390400
transform 1 0 1568 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_11
timestamp 1669390400
transform 1 0 2576 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_21
timestamp 1669390400
transform 1 0 3696 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_27
timestamp 1669390400
transform 1 0 4368 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_31
timestamp 1669390400
transform 1 0 4816 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_35
timestamp 1669390400
transform 1 0 5264 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_42
timestamp 1669390400
transform 1 0 6048 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_44
timestamp 1669390400
transform 1 0 6272 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_47
timestamp 1669390400
transform 1 0 6608 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_60
timestamp 1669390400
transform 1 0 8064 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_70
timestamp 1669390400
transform 1 0 9184 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_73
timestamp 1669390400
transform 1 0 9520 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_76
timestamp 1669390400
transform 1 0 9856 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_84
timestamp 1669390400
transform 1 0 10752 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_98
timestamp 1669390400
transform 1 0 12320 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_102
timestamp 1669390400
transform 1 0 12768 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_106
timestamp 1669390400
transform 1 0 13216 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_113
timestamp 1669390400
transform 1 0 14000 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_120
timestamp 1669390400
transform 1 0 14784 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_127
timestamp 1669390400
transform 1 0 15568 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_131
timestamp 1669390400
transform 1 0 16016 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_141
timestamp 1669390400
transform 1 0 17136 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_144
timestamp 1669390400
transform 1 0 17472 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_147
timestamp 1669390400
transform 1 0 17808 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_157
timestamp 1669390400
transform 1 0 18928 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_161
timestamp 1669390400
transform 1 0 19376 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_165
timestamp 1669390400
transform 1 0 19824 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_169
timestamp 1669390400
transform 1 0 20272 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_181
timestamp 1669390400
transform 1 0 21616 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_185
timestamp 1669390400
transform 1 0 22064 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_188
timestamp 1669390400
transform 1 0 22400 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_192
timestamp 1669390400
transform 1 0 22848 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_212
timestamp 1669390400
transform 1 0 25088 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_215
timestamp 1669390400
transform 1 0 25424 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_218
timestamp 1669390400
transform 1 0 25760 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_222
timestamp 1669390400
transform 1 0 26208 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_232
timestamp 1669390400
transform 1 0 27328 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_239
timestamp 1669390400
transform 1 0 28112 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_245
timestamp 1669390400
transform 1 0 28784 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_249
timestamp 1669390400
transform 1 0 29232 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_260
timestamp 1669390400
transform 1 0 30464 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_262
timestamp 1669390400
transform 1 0 30688 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_265
timestamp 1669390400
transform 1 0 31024 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_273
timestamp 1669390400
transform 1 0 31920 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_283
timestamp 1669390400
transform 1 0 33040 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_286
timestamp 1669390400
transform 1 0 33376 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_289
timestamp 1669390400
transform 1 0 33712 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_303
timestamp 1669390400
transform 1 0 35280 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_307
timestamp 1669390400
transform 1 0 35728 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_311
timestamp 1669390400
transform 1 0 36176 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_315
timestamp 1669390400
transform 1 0 36624 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_319
timestamp 1669390400
transform 1 0 37072 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_323
timestamp 1669390400
transform 1 0 37520 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_327
timestamp 1669390400
transform 1 0 37968 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_329
timestamp 1669390400
transform 1 0 38192 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_332
timestamp 1669390400
transform 1 0 38528 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_353
timestamp 1669390400
transform 1 0 40880 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_357
timestamp 1669390400
transform 1 0 41328 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_376
timestamp 1669390400
transform 1 0 43456 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_390
timestamp 1669390400
transform 1 0 45024 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_402
timestamp 1669390400
transform 1 0 46368 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_404
timestamp 1669390400
transform 1 0 46592 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_415
timestamp 1669390400
transform 1 0 47824 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_422
timestamp 1669390400
transform 1 0 48608 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_428
timestamp 1669390400
transform 1 0 49280 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_432
timestamp 1669390400
transform 1 0 49728 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_436
timestamp 1669390400
transform 1 0 50176 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_438
timestamp 1669390400
transform 1 0 50400 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_444
timestamp 1669390400
transform 1 0 51072 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_460
timestamp 1669390400
transform 1 0 52864 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_464
timestamp 1669390400
transform 1 0 53312 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_468
timestamp 1669390400
transform 1 0 53760 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_472
timestamp 1669390400
transform 1 0 54208 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_476
timestamp 1669390400
transform 1 0 54656 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_492
timestamp 1669390400
transform 1 0 56448 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_496
timestamp 1669390400
transform 1 0 56896 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_499
timestamp 1669390400
transform 1 0 57232 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_506
timestamp 1669390400
transform 1 0 58016 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_510
timestamp 1669390400
transform 1 0 58464 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_512
timestamp 1669390400
transform 1 0 58688 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_2
timestamp 1669390400
transform 1 0 1568 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_8
timestamp 1669390400
transform 1 0 2240 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_12
timestamp 1669390400
transform 1 0 2688 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_25
timestamp 1669390400
transform 1 0 4144 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_27
timestamp 1669390400
transform 1 0 4368 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_30
timestamp 1669390400
transform 1 0 4704 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_34
timestamp 1669390400
transform 1 0 5152 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_37
timestamp 1669390400
transform 1 0 5488 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_57
timestamp 1669390400
transform 1 0 7728 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_61
timestamp 1669390400
transform 1 0 8176 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_64
timestamp 1669390400
transform 1 0 8512 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_78
timestamp 1669390400
transform 1 0 10080 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_82
timestamp 1669390400
transform 1 0 10528 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_85
timestamp 1669390400
transform 1 0 10864 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_89
timestamp 1669390400
transform 1 0 11312 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_93
timestamp 1669390400
transform 1 0 11760 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_97
timestamp 1669390400
transform 1 0 12208 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_101
timestamp 1669390400
transform 1 0 12656 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_105
timestamp 1669390400
transform 1 0 13104 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_108
timestamp 1669390400
transform 1 0 13440 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_122
timestamp 1669390400
transform 1 0 15008 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_128
timestamp 1669390400
transform 1 0 15680 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_132
timestamp 1669390400
transform 1 0 16128 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_136
timestamp 1669390400
transform 1 0 16576 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_140
timestamp 1669390400
transform 1 0 17024 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_144
timestamp 1669390400
transform 1 0 17472 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_148
timestamp 1669390400
transform 1 0 17920 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_152
timestamp 1669390400
transform 1 0 18368 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_156
timestamp 1669390400
transform 1 0 18816 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_166
timestamp 1669390400
transform 1 0 19936 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_170
timestamp 1669390400
transform 1 0 20384 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_176
timestamp 1669390400
transform 1 0 21056 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_179
timestamp 1669390400
transform 1 0 21392 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_182
timestamp 1669390400
transform 1 0 21728 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_186
timestamp 1669390400
transform 1 0 22176 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_189
timestamp 1669390400
transform 1 0 22512 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_193
timestamp 1669390400
transform 1 0 22960 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_197
timestamp 1669390400
transform 1 0 23408 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_201
timestamp 1669390400
transform 1 0 23856 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_215
timestamp 1669390400
transform 1 0 25424 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_219
timestamp 1669390400
transform 1 0 25872 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_233
timestamp 1669390400
transform 1 0 27440 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_247
timestamp 1669390400
transform 1 0 29008 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_250
timestamp 1669390400
transform 1 0 29344 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_278
timestamp 1669390400
transform 1 0 32480 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_282
timestamp 1669390400
transform 1 0 32928 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_299
timestamp 1669390400
transform 1 0 34832 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_303
timestamp 1669390400
transform 1 0 35280 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_307
timestamp 1669390400
transform 1 0 35728 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_318
timestamp 1669390400
transform 1 0 36960 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_321
timestamp 1669390400
transform 1 0 37296 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_334
timestamp 1669390400
transform 1 0 38752 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_338
timestamp 1669390400
transform 1 0 39200 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_347
timestamp 1669390400
transform 1 0 40208 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_354
timestamp 1669390400
transform 1 0 40992 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_358
timestamp 1669390400
transform 1 0 41440 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_362
timestamp 1669390400
transform 1 0 41888 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_366
timestamp 1669390400
transform 1 0 42336 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_370
timestamp 1669390400
transform 1 0 42784 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_374
timestamp 1669390400
transform 1 0 43232 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_381
timestamp 1669390400
transform 1 0 44016 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_388
timestamp 1669390400
transform 1 0 44800 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_392
timestamp 1669390400
transform 1 0 45248 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_395
timestamp 1669390400
transform 1 0 45584 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_415
timestamp 1669390400
transform 1 0 47824 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_432
timestamp 1669390400
transform 1 0 49728 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_439
timestamp 1669390400
transform 1 0 50512 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_443
timestamp 1669390400
transform 1 0 50960 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_447
timestamp 1669390400
transform 1 0 51408 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_453
timestamp 1669390400
transform 1 0 52080 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_457
timestamp 1669390400
transform 1 0 52528 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_460
timestamp 1669390400
transform 1 0 52864 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_463
timestamp 1669390400
transform 1 0 53200 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_470
timestamp 1669390400
transform 1 0 53984 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_480
timestamp 1669390400
transform 1 0 55104 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_484
timestamp 1669390400
transform 1 0 55552 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_488
timestamp 1669390400
transform 1 0 56000 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_492
timestamp 1669390400
transform 1 0 56448 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_495
timestamp 1669390400
transform 1 0 56784 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_505
timestamp 1669390400
transform 1 0 57904 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_2
timestamp 1669390400
transform 1 0 1568 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_4
timestamp 1669390400
transform 1 0 1792 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_7
timestamp 1669390400
transform 1 0 2128 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_17
timestamp 1669390400
transform 1 0 3248 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_27
timestamp 1669390400
transform 1 0 4368 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_31
timestamp 1669390400
transform 1 0 4816 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_34
timestamp 1669390400
transform 1 0 5152 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_38
timestamp 1669390400
transform 1 0 5600 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_42
timestamp 1669390400
transform 1 0 6048 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_61
timestamp 1669390400
transform 1 0 8176 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_69
timestamp 1669390400
transform 1 0 9072 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_73
timestamp 1669390400
transform 1 0 9520 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_76
timestamp 1669390400
transform 1 0 9856 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_80
timestamp 1669390400
transform 1 0 10304 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_90
timestamp 1669390400
transform 1 0 11424 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_94
timestamp 1669390400
transform 1 0 11872 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_97
timestamp 1669390400
transform 1 0 12208 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_101
timestamp 1669390400
transform 1 0 12656 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_111
timestamp 1669390400
transform 1 0 13776 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_125
timestamp 1669390400
transform 1 0 15344 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_129
timestamp 1669390400
transform 1 0 15792 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_133
timestamp 1669390400
transform 1 0 16240 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_137
timestamp 1669390400
transform 1 0 16688 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_141
timestamp 1669390400
transform 1 0 17136 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_144
timestamp 1669390400
transform 1 0 17472 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_151
timestamp 1669390400
transform 1 0 18256 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_157
timestamp 1669390400
transform 1 0 18928 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_168
timestamp 1669390400
transform 1 0 20160 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_178
timestamp 1669390400
transform 1 0 21280 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_190
timestamp 1669390400
transform 1 0 22624 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_194
timestamp 1669390400
transform 1 0 23072 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_196
timestamp 1669390400
transform 1 0 23296 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_212
timestamp 1669390400
transform 1 0 25088 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_215
timestamp 1669390400
transform 1 0 25424 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_217
timestamp 1669390400
transform 1 0 25648 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_220
timestamp 1669390400
transform 1 0 25984 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_238
timestamp 1669390400
transform 1 0 28000 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_255
timestamp 1669390400
transform 1 0 29904 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_259
timestamp 1669390400
transform 1 0 30352 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_268
timestamp 1669390400
transform 1 0 31360 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_270
timestamp 1669390400
transform 1 0 31584 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_273
timestamp 1669390400
transform 1 0 31920 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_283
timestamp 1669390400
transform 1 0 33040 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_286
timestamp 1669390400
transform 1 0 33376 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_288
timestamp 1669390400
transform 1 0 33600 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_299
timestamp 1669390400
transform 1 0 34832 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_303
timestamp 1669390400
transform 1 0 35280 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_316
timestamp 1669390400
transform 1 0 36736 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_327
timestamp 1669390400
transform 1 0 37968 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_334
timestamp 1669390400
transform 1 0 38752 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_336
timestamp 1669390400
transform 1 0 38976 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_350
timestamp 1669390400
transform 1 0 40544 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_354
timestamp 1669390400
transform 1 0 40992 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_357
timestamp 1669390400
transform 1 0 41328 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_360
timestamp 1669390400
transform 1 0 41664 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_362
timestamp 1669390400
transform 1 0 41888 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_369
timestamp 1669390400
transform 1 0 42672 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_377
timestamp 1669390400
transform 1 0 43568 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_381
timestamp 1669390400
transform 1 0 44016 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_390
timestamp 1669390400
transform 1 0 45024 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_394
timestamp 1669390400
transform 1 0 45472 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_398
timestamp 1669390400
transform 1 0 45920 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_400
timestamp 1669390400
transform 1 0 46144 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_411
timestamp 1669390400
transform 1 0 47376 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_425
timestamp 1669390400
transform 1 0 48944 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_428
timestamp 1669390400
transform 1 0 49280 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_453
timestamp 1669390400
transform 1 0 52080 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_466
timestamp 1669390400
transform 1 0 53536 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_478
timestamp 1669390400
transform 1 0 54880 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_495
timestamp 1669390400
transform 1 0 56784 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_499
timestamp 1669390400
transform 1 0 57232 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_512
timestamp 1669390400
transform 1 0 58688 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_2
timestamp 1669390400
transform 1 0 1568 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_8
timestamp 1669390400
transform 1 0 2240 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_12
timestamp 1669390400
transform 1 0 2688 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_16
timestamp 1669390400
transform 1 0 3136 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_25
timestamp 1669390400
transform 1 0 4144 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_27
timestamp 1669390400
transform 1 0 4368 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_30
timestamp 1669390400
transform 1 0 4704 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_34
timestamp 1669390400
transform 1 0 5152 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_37
timestamp 1669390400
transform 1 0 5488 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_51
timestamp 1669390400
transform 1 0 7056 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_55
timestamp 1669390400
transform 1 0 7504 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_61
timestamp 1669390400
transform 1 0 8176 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_72
timestamp 1669390400
transform 1 0 9408 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_78
timestamp 1669390400
transform 1 0 10080 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_82
timestamp 1669390400
transform 1 0 10528 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_99
timestamp 1669390400
transform 1 0 12432 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_105
timestamp 1669390400
transform 1 0 13104 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_108
timestamp 1669390400
transform 1 0 13440 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_118
timestamp 1669390400
transform 1 0 14560 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_122
timestamp 1669390400
transform 1 0 15008 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_125
timestamp 1669390400
transform 1 0 15344 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_137
timestamp 1669390400
transform 1 0 16688 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_149
timestamp 1669390400
transform 1 0 18032 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_157
timestamp 1669390400
transform 1 0 18928 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_161
timestamp 1669390400
transform 1 0 19376 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_164
timestamp 1669390400
transform 1 0 19712 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_168
timestamp 1669390400
transform 1 0 20160 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_172
timestamp 1669390400
transform 1 0 20608 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_176
timestamp 1669390400
transform 1 0 21056 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_179
timestamp 1669390400
transform 1 0 21392 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_190
timestamp 1669390400
transform 1 0 22624 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_192
timestamp 1669390400
transform 1 0 22848 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_195
timestamp 1669390400
transform 1 0 23184 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_215
timestamp 1669390400
transform 1 0 25424 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_229
timestamp 1669390400
transform 1 0 26992 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_235
timestamp 1669390400
transform 1 0 27664 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_239
timestamp 1669390400
transform 1 0 28112 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_243
timestamp 1669390400
transform 1 0 28560 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_247
timestamp 1669390400
transform 1 0 29008 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_250
timestamp 1669390400
transform 1 0 29344 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_252
timestamp 1669390400
transform 1 0 29568 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_258
timestamp 1669390400
transform 1 0 30240 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_262
timestamp 1669390400
transform 1 0 30688 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_265
timestamp 1669390400
transform 1 0 31024 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_318
timestamp 1669390400
transform 1 0 36960 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_321
timestamp 1669390400
transform 1 0 37296 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_323
timestamp 1669390400
transform 1 0 37520 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_329
timestamp 1669390400
transform 1 0 38192 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_345
timestamp 1669390400
transform 1 0 39984 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_354
timestamp 1669390400
transform 1 0 40992 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_358
timestamp 1669390400
transform 1 0 41440 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_360
timestamp 1669390400
transform 1 0 41664 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_363
timestamp 1669390400
transform 1 0 42000 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_367
timestamp 1669390400
transform 1 0 42448 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_371
timestamp 1669390400
transform 1 0 42896 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_377
timestamp 1669390400
transform 1 0 43568 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_385
timestamp 1669390400
transform 1 0 44464 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_389
timestamp 1669390400
transform 1 0 44912 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_392
timestamp 1669390400
transform 1 0 45248 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_401
timestamp 1669390400
transform 1 0 46256 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_405
timestamp 1669390400
transform 1 0 46704 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_417
timestamp 1669390400
transform 1 0 48048 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_421
timestamp 1669390400
transform 1 0 48496 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_430
timestamp 1669390400
transform 1 0 49504 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_50_434
timestamp 1669390400
transform 1 0 49952 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_450
timestamp 1669390400
transform 1 0 51744 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_452
timestamp 1669390400
transform 1 0 51968 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_455
timestamp 1669390400
transform 1 0 52304 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_459
timestamp 1669390400
transform 1 0 52752 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_463
timestamp 1669390400
transform 1 0 53200 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_472
timestamp 1669390400
transform 1 0 54208 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_476
timestamp 1669390400
transform 1 0 54656 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_485
timestamp 1669390400
transform 1 0 55664 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_492
timestamp 1669390400
transform 1 0 56448 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_496
timestamp 1669390400
transform 1 0 56896 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_500
timestamp 1669390400
transform 1 0 57344 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_504
timestamp 1669390400
transform 1 0 57792 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_512
timestamp 1669390400
transform 1 0 58688 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_2
timestamp 1669390400
transform 1 0 1568 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_12
timestamp 1669390400
transform 1 0 2688 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_29
timestamp 1669390400
transform 1 0 4592 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_31
timestamp 1669390400
transform 1 0 4816 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_40
timestamp 1669390400
transform 1 0 5824 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_46
timestamp 1669390400
transform 1 0 6496 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_50
timestamp 1669390400
transform 1 0 6944 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_54
timestamp 1669390400
transform 1 0 7392 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_58
timestamp 1669390400
transform 1 0 7840 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_62
timestamp 1669390400
transform 1 0 8288 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_66
timestamp 1669390400
transform 1 0 8736 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_70
timestamp 1669390400
transform 1 0 9184 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_73
timestamp 1669390400
transform 1 0 9520 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_85
timestamp 1669390400
transform 1 0 10864 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_89
timestamp 1669390400
transform 1 0 11312 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_92
timestamp 1669390400
transform 1 0 11648 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_106
timestamp 1669390400
transform 1 0 13216 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_110
timestamp 1669390400
transform 1 0 13664 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_114
timestamp 1669390400
transform 1 0 14112 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_124
timestamp 1669390400
transform 1 0 15232 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_128
timestamp 1669390400
transform 1 0 15680 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_140
timestamp 1669390400
transform 1 0 17024 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_144
timestamp 1669390400
transform 1 0 17472 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_151
timestamp 1669390400
transform 1 0 18256 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_165
timestamp 1669390400
transform 1 0 19824 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_186
timestamp 1669390400
transform 1 0 22176 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_192
timestamp 1669390400
transform 1 0 22848 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_196
timestamp 1669390400
transform 1 0 23296 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_200
timestamp 1669390400
transform 1 0 23744 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_204
timestamp 1669390400
transform 1 0 24192 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_208
timestamp 1669390400
transform 1 0 24640 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_212
timestamp 1669390400
transform 1 0 25088 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_215
timestamp 1669390400
transform 1 0 25424 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_221
timestamp 1669390400
transform 1 0 26096 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_225
timestamp 1669390400
transform 1 0 26544 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_229
timestamp 1669390400
transform 1 0 26992 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_233
timestamp 1669390400
transform 1 0 27440 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_244
timestamp 1669390400
transform 1 0 28672 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_250
timestamp 1669390400
transform 1 0 29344 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_254
timestamp 1669390400
transform 1 0 29792 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_260
timestamp 1669390400
transform 1 0 30464 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_272
timestamp 1669390400
transform 1 0 31808 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_276
timestamp 1669390400
transform 1 0 32256 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_283
timestamp 1669390400
transform 1 0 33040 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_286
timestamp 1669390400
transform 1 0 33376 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_289
timestamp 1669390400
transform 1 0 33712 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_291
timestamp 1669390400
transform 1 0 33936 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_307
timestamp 1669390400
transform 1 0 35728 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_311
timestamp 1669390400
transform 1 0 36176 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_315
timestamp 1669390400
transform 1 0 36624 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_319
timestamp 1669390400
transform 1 0 37072 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_323
timestamp 1669390400
transform 1 0 37520 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_327
timestamp 1669390400
transform 1 0 37968 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_331
timestamp 1669390400
transform 1 0 38416 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_335
timestamp 1669390400
transform 1 0 38864 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_339
timestamp 1669390400
transform 1 0 39312 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_343
timestamp 1669390400
transform 1 0 39760 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_354
timestamp 1669390400
transform 1 0 40992 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_357
timestamp 1669390400
transform 1 0 41328 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_360
timestamp 1669390400
transform 1 0 41664 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_375
timestamp 1669390400
transform 1 0 43344 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_383
timestamp 1669390400
transform 1 0 44240 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_387
timestamp 1669390400
transform 1 0 44688 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_391
timestamp 1669390400
transform 1 0 45136 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_395
timestamp 1669390400
transform 1 0 45584 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_401
timestamp 1669390400
transform 1 0 46256 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_405
timestamp 1669390400
transform 1 0 46704 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_409
timestamp 1669390400
transform 1 0 47152 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_413
timestamp 1669390400
transform 1 0 47600 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_417
timestamp 1669390400
transform 1 0 48048 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_421
timestamp 1669390400
transform 1 0 48496 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_425
timestamp 1669390400
transform 1 0 48944 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_51_428
timestamp 1669390400
transform 1 0 49280 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_460
timestamp 1669390400
transform 1 0 52864 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_468
timestamp 1669390400
transform 1 0 53760 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_483
timestamp 1669390400
transform 1 0 55440 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_496
timestamp 1669390400
transform 1 0 56896 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_499
timestamp 1669390400
transform 1 0 57232 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_512
timestamp 1669390400
transform 1 0 58688 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_2
timestamp 1669390400
transform 1 0 1568 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_18
timestamp 1669390400
transform 1 0 3360 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_29
timestamp 1669390400
transform 1 0 4592 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_31
timestamp 1669390400
transform 1 0 4816 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_34
timestamp 1669390400
transform 1 0 5152 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_37
timestamp 1669390400
transform 1 0 5488 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_50
timestamp 1669390400
transform 1 0 6944 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_56
timestamp 1669390400
transform 1 0 7616 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_60
timestamp 1669390400
transform 1 0 8064 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_75
timestamp 1669390400
transform 1 0 9744 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_90
timestamp 1669390400
transform 1 0 11424 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_102
timestamp 1669390400
transform 1 0 12768 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_108
timestamp 1669390400
transform 1 0 13440 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_110
timestamp 1669390400
transform 1 0 13664 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_113
timestamp 1669390400
transform 1 0 14000 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_124
timestamp 1669390400
transform 1 0 15232 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_136
timestamp 1669390400
transform 1 0 16576 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_140
timestamp 1669390400
transform 1 0 17024 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_144
timestamp 1669390400
transform 1 0 17472 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_154
timestamp 1669390400
transform 1 0 18592 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_164
timestamp 1669390400
transform 1 0 19712 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_176
timestamp 1669390400
transform 1 0 21056 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_179
timestamp 1669390400
transform 1 0 21392 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_190
timestamp 1669390400
transform 1 0 22624 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_192
timestamp 1669390400
transform 1 0 22848 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_195
timestamp 1669390400
transform 1 0 23184 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_199
timestamp 1669390400
transform 1 0 23632 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_203
timestamp 1669390400
transform 1 0 24080 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_213
timestamp 1669390400
transform 1 0 25200 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_217
timestamp 1669390400
transform 1 0 25648 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_220
timestamp 1669390400
transform 1 0 25984 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_230
timestamp 1669390400
transform 1 0 27104 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_242
timestamp 1669390400
transform 1 0 28448 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_244
timestamp 1669390400
transform 1 0 28672 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_247
timestamp 1669390400
transform 1 0 29008 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_250
timestamp 1669390400
transform 1 0 29344 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_253
timestamp 1669390400
transform 1 0 29680 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_261
timestamp 1669390400
transform 1 0 30576 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_265
timestamp 1669390400
transform 1 0 31024 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_318
timestamp 1669390400
transform 1 0 36960 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_321
timestamp 1669390400
transform 1 0 37296 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_336
timestamp 1669390400
transform 1 0 38976 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_340
timestamp 1669390400
transform 1 0 39424 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_349
timestamp 1669390400
transform 1 0 40432 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_353
timestamp 1669390400
transform 1 0 40880 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_360
timestamp 1669390400
transform 1 0 41664 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_364
timestamp 1669390400
transform 1 0 42112 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_378
timestamp 1669390400
transform 1 0 43680 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_380
timestamp 1669390400
transform 1 0 43904 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_389
timestamp 1669390400
transform 1 0 44912 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_392
timestamp 1669390400
transform 1 0 45248 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_406
timestamp 1669390400
transform 1 0 46816 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_414
timestamp 1669390400
transform 1 0 47712 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_428
timestamp 1669390400
transform 1 0 49280 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_438
timestamp 1669390400
transform 1 0 50400 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_454
timestamp 1669390400
transform 1 0 52192 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_458
timestamp 1669390400
transform 1 0 52640 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_460
timestamp 1669390400
transform 1 0 52864 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_463
timestamp 1669390400
transform 1 0 53200 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_479
timestamp 1669390400
transform 1 0 54992 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_487
timestamp 1669390400
transform 1 0 55888 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_501
timestamp 1669390400
transform 1 0 57456 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_505
timestamp 1669390400
transform 1 0 57904 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_2
timestamp 1669390400
transform 1 0 1568 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_12
timestamp 1669390400
transform 1 0 2688 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_22
timestamp 1669390400
transform 1 0 3808 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_30
timestamp 1669390400
transform 1 0 4704 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_37
timestamp 1669390400
transform 1 0 5488 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_41
timestamp 1669390400
transform 1 0 5936 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_44
timestamp 1669390400
transform 1 0 6272 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_57
timestamp 1669390400
transform 1 0 7728 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_67
timestamp 1669390400
transform 1 0 8848 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_73
timestamp 1669390400
transform 1 0 9520 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_76
timestamp 1669390400
transform 1 0 9856 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_80
timestamp 1669390400
transform 1 0 10304 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_95
timestamp 1669390400
transform 1 0 11984 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_123
timestamp 1669390400
transform 1 0 15120 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_129
timestamp 1669390400
transform 1 0 15792 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_133
timestamp 1669390400
transform 1 0 16240 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_137
timestamp 1669390400
transform 1 0 16688 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_141
timestamp 1669390400
transform 1 0 17136 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_144
timestamp 1669390400
transform 1 0 17472 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_154
timestamp 1669390400
transform 1 0 18592 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_158
timestamp 1669390400
transform 1 0 19040 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_162
timestamp 1669390400
transform 1 0 19488 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_187
timestamp 1669390400
transform 1 0 22288 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_193
timestamp 1669390400
transform 1 0 22960 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_197
timestamp 1669390400
transform 1 0 23408 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_208
timestamp 1669390400
transform 1 0 24640 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_212
timestamp 1669390400
transform 1 0 25088 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_215
timestamp 1669390400
transform 1 0 25424 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_222
timestamp 1669390400
transform 1 0 26208 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_226
timestamp 1669390400
transform 1 0 26656 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_239
timestamp 1669390400
transform 1 0 28112 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_241
timestamp 1669390400
transform 1 0 28336 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_254
timestamp 1669390400
transform 1 0 29792 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_265
timestamp 1669390400
transform 1 0 31024 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_275
timestamp 1669390400
transform 1 0 32144 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_279
timestamp 1669390400
transform 1 0 32592 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_283
timestamp 1669390400
transform 1 0 33040 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_286
timestamp 1669390400
transform 1 0 33376 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_289
timestamp 1669390400
transform 1 0 33712 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_293
timestamp 1669390400
transform 1 0 34160 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_303
timestamp 1669390400
transform 1 0 35280 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_317
timestamp 1669390400
transform 1 0 36848 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_321
timestamp 1669390400
transform 1 0 37296 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_325
timestamp 1669390400
transform 1 0 37744 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_332
timestamp 1669390400
transform 1 0 38528 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_336
timestamp 1669390400
transform 1 0 38976 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_340
timestamp 1669390400
transform 1 0 39424 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_346
timestamp 1669390400
transform 1 0 40096 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_350
timestamp 1669390400
transform 1 0 40544 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_354
timestamp 1669390400
transform 1 0 40992 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_357
timestamp 1669390400
transform 1 0 41328 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_360
timestamp 1669390400
transform 1 0 41664 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_364
timestamp 1669390400
transform 1 0 42112 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_373
timestamp 1669390400
transform 1 0 43120 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_379
timestamp 1669390400
transform 1 0 43792 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_386
timestamp 1669390400
transform 1 0 44576 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_394
timestamp 1669390400
transform 1 0 45472 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_398
timestamp 1669390400
transform 1 0 45920 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_414
timestamp 1669390400
transform 1 0 47712 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_416
timestamp 1669390400
transform 1 0 47936 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_425
timestamp 1669390400
transform 1 0 48944 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_428
timestamp 1669390400
transform 1 0 49280 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_441
timestamp 1669390400
transform 1 0 50736 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_462
timestamp 1669390400
transform 1 0 53088 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_472
timestamp 1669390400
transform 1 0 54208 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_488
timestamp 1669390400
transform 1 0 56000 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_495
timestamp 1669390400
transform 1 0 56784 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_499
timestamp 1669390400
transform 1 0 57232 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_508
timestamp 1669390400
transform 1 0 58240 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_512
timestamp 1669390400
transform 1 0 58688 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_2
timestamp 1669390400
transform 1 0 1568 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_6
timestamp 1669390400
transform 1 0 2016 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_23
timestamp 1669390400
transform 1 0 3920 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_25
timestamp 1669390400
transform 1 0 4144 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_31
timestamp 1669390400
transform 1 0 4816 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_37
timestamp 1669390400
transform 1 0 5488 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_39
timestamp 1669390400
transform 1 0 5712 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_42
timestamp 1669390400
transform 1 0 6048 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_53
timestamp 1669390400
transform 1 0 7280 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_63
timestamp 1669390400
transform 1 0 8400 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_70
timestamp 1669390400
transform 1 0 9184 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_74
timestamp 1669390400
transform 1 0 9632 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_77
timestamp 1669390400
transform 1 0 9968 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_105
timestamp 1669390400
transform 1 0 13104 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_108
timestamp 1669390400
transform 1 0 13440 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_110
timestamp 1669390400
transform 1 0 13664 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_116
timestamp 1669390400
transform 1 0 14336 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_133
timestamp 1669390400
transform 1 0 16240 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_135
timestamp 1669390400
transform 1 0 16464 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_176
timestamp 1669390400
transform 1 0 21056 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_179
timestamp 1669390400
transform 1 0 21392 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_182
timestamp 1669390400
transform 1 0 21728 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_184
timestamp 1669390400
transform 1 0 21952 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_187
timestamp 1669390400
transform 1 0 22288 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_199
timestamp 1669390400
transform 1 0 23632 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_211
timestamp 1669390400
transform 1 0 24976 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_221
timestamp 1669390400
transform 1 0 26096 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_225
timestamp 1669390400
transform 1 0 26544 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_234
timestamp 1669390400
transform 1 0 27552 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_236
timestamp 1669390400
transform 1 0 27776 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_239
timestamp 1669390400
transform 1 0 28112 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_243
timestamp 1669390400
transform 1 0 28560 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_247
timestamp 1669390400
transform 1 0 29008 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_250
timestamp 1669390400
transform 1 0 29344 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_257
timestamp 1669390400
transform 1 0 30128 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_264
timestamp 1669390400
transform 1 0 30912 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_268
timestamp 1669390400
transform 1 0 31360 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_272
timestamp 1669390400
transform 1 0 31808 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_274
timestamp 1669390400
transform 1 0 32032 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_277
timestamp 1669390400
transform 1 0 32368 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_289
timestamp 1669390400
transform 1 0 33712 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_299
timestamp 1669390400
transform 1 0 34832 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_309
timestamp 1669390400
transform 1 0 35952 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_313
timestamp 1669390400
transform 1 0 36400 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_317
timestamp 1669390400
transform 1 0 36848 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_321
timestamp 1669390400
transform 1 0 37296 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_335
timestamp 1669390400
transform 1 0 38864 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_337
timestamp 1669390400
transform 1 0 39088 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_344
timestamp 1669390400
transform 1 0 39872 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_348
timestamp 1669390400
transform 1 0 40320 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_352
timestamp 1669390400
transform 1 0 40768 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_354
timestamp 1669390400
transform 1 0 40992 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_367
timestamp 1669390400
transform 1 0 42448 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_375
timestamp 1669390400
transform 1 0 43344 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_379
timestamp 1669390400
transform 1 0 43792 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_381
timestamp 1669390400
transform 1 0 44016 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_384
timestamp 1669390400
transform 1 0 44352 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_388
timestamp 1669390400
transform 1 0 44800 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_392
timestamp 1669390400
transform 1 0 45248 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_401
timestamp 1669390400
transform 1 0 46256 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_408
timestamp 1669390400
transform 1 0 47040 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_416
timestamp 1669390400
transform 1 0 47936 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_420
timestamp 1669390400
transform 1 0 48384 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_433
timestamp 1669390400
transform 1 0 49840 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_441
timestamp 1669390400
transform 1 0 50736 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_453
timestamp 1669390400
transform 1 0 52080 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_463
timestamp 1669390400
transform 1 0 53200 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_476
timestamp 1669390400
transform 1 0 54656 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_480
timestamp 1669390400
transform 1 0 55104 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_482
timestamp 1669390400
transform 1 0 55328 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_491
timestamp 1669390400
transform 1 0 56336 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_495
timestamp 1669390400
transform 1 0 56784 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_499
timestamp 1669390400
transform 1 0 57232 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_508
timestamp 1669390400
transform 1 0 58240 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_512
timestamp 1669390400
transform 1 0 58688 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_2
timestamp 1669390400
transform 1 0 1568 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_6
timestamp 1669390400
transform 1 0 2016 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_10
timestamp 1669390400
transform 1 0 2464 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_14
timestamp 1669390400
transform 1 0 2912 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_21
timestamp 1669390400
transform 1 0 3696 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_27
timestamp 1669390400
transform 1 0 4368 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_35
timestamp 1669390400
transform 1 0 5264 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_37
timestamp 1669390400
transform 1 0 5488 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_40
timestamp 1669390400
transform 1 0 5824 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_44
timestamp 1669390400
transform 1 0 6272 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_54
timestamp 1669390400
transform 1 0 7392 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_58
timestamp 1669390400
transform 1 0 7840 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_62
timestamp 1669390400
transform 1 0 8288 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_70
timestamp 1669390400
transform 1 0 9184 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_73
timestamp 1669390400
transform 1 0 9520 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_76
timestamp 1669390400
transform 1 0 9856 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_86
timestamp 1669390400
transform 1 0 10976 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_96
timestamp 1669390400
transform 1 0 12096 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_106
timestamp 1669390400
transform 1 0 13216 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_110
timestamp 1669390400
transform 1 0 13664 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_121
timestamp 1669390400
transform 1 0 14896 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_131
timestamp 1669390400
transform 1 0 16016 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_141
timestamp 1669390400
transform 1 0 17136 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_144
timestamp 1669390400
transform 1 0 17472 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_186
timestamp 1669390400
transform 1 0 22176 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_188
timestamp 1669390400
transform 1 0 22400 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_191
timestamp 1669390400
transform 1 0 22736 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_195
timestamp 1669390400
transform 1 0 23184 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_206
timestamp 1669390400
transform 1 0 24416 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_212
timestamp 1669390400
transform 1 0 25088 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_215
timestamp 1669390400
transform 1 0 25424 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_224
timestamp 1669390400
transform 1 0 26432 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_277
timestamp 1669390400
transform 1 0 32368 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_281
timestamp 1669390400
transform 1 0 32816 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_283
timestamp 1669390400
transform 1 0 33040 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_286
timestamp 1669390400
transform 1 0 33376 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_295
timestamp 1669390400
transform 1 0 34384 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_299
timestamp 1669390400
transform 1 0 34832 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_313
timestamp 1669390400
transform 1 0 36400 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_320
timestamp 1669390400
transform 1 0 37184 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_329
timestamp 1669390400
transform 1 0 38192 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_333
timestamp 1669390400
transform 1 0 38640 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_347
timestamp 1669390400
transform 1 0 40208 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_357
timestamp 1669390400
transform 1 0 41328 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_365
timestamp 1669390400
transform 1 0 42224 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_369
timestamp 1669390400
transform 1 0 42672 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_385
timestamp 1669390400
transform 1 0 44464 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_397
timestamp 1669390400
transform 1 0 45808 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_405
timestamp 1669390400
transform 1 0 46704 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_407
timestamp 1669390400
transform 1 0 46928 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_410
timestamp 1669390400
transform 1 0 47264 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_425
timestamp 1669390400
transform 1 0 48944 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_428
timestamp 1669390400
transform 1 0 49280 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_437
timestamp 1669390400
transform 1 0 50288 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_453
timestamp 1669390400
transform 1 0 52080 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_467
timestamp 1669390400
transform 1 0 53648 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_471
timestamp 1669390400
transform 1 0 54096 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_490
timestamp 1669390400
transform 1 0 56224 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_494
timestamp 1669390400
transform 1 0 56672 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_496
timestamp 1669390400
transform 1 0 56896 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_499
timestamp 1669390400
transform 1 0 57232 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_512
timestamp 1669390400
transform 1 0 58688 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_2
timestamp 1669390400
transform 1 0 1568 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_5
timestamp 1669390400
transform 1 0 1904 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_15
timestamp 1669390400
transform 1 0 3024 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_27
timestamp 1669390400
transform 1 0 4368 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_31
timestamp 1669390400
transform 1 0 4816 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_34
timestamp 1669390400
transform 1 0 5152 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_37
timestamp 1669390400
transform 1 0 5488 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_60
timestamp 1669390400
transform 1 0 8064 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_64
timestamp 1669390400
transform 1 0 8512 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_67
timestamp 1669390400
transform 1 0 8848 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_80
timestamp 1669390400
transform 1 0 10304 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_92
timestamp 1669390400
transform 1 0 11648 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_94
timestamp 1669390400
transform 1 0 11872 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_97
timestamp 1669390400
transform 1 0 12208 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_101
timestamp 1669390400
transform 1 0 12656 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_105
timestamp 1669390400
transform 1 0 13104 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_108
timestamp 1669390400
transform 1 0 13440 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_119
timestamp 1669390400
transform 1 0 14672 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_125
timestamp 1669390400
transform 1 0 15344 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_135
timestamp 1669390400
transform 1 0 16464 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_158
timestamp 1669390400
transform 1 0 19040 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_162
timestamp 1669390400
transform 1 0 19488 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_174
timestamp 1669390400
transform 1 0 20832 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_176
timestamp 1669390400
transform 1 0 21056 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_179
timestamp 1669390400
transform 1 0 21392 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_182
timestamp 1669390400
transform 1 0 21728 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_186
timestamp 1669390400
transform 1 0 22176 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_190
timestamp 1669390400
transform 1 0 22624 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_194
timestamp 1669390400
transform 1 0 23072 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_198
timestamp 1669390400
transform 1 0 23520 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_202
timestamp 1669390400
transform 1 0 23968 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_212
timestamp 1669390400
transform 1 0 25088 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_216
timestamp 1669390400
transform 1 0 25536 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_219
timestamp 1669390400
transform 1 0 25872 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_223
timestamp 1669390400
transform 1 0 26320 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_227
timestamp 1669390400
transform 1 0 26768 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_237
timestamp 1669390400
transform 1 0 27888 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_243
timestamp 1669390400
transform 1 0 28560 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_247
timestamp 1669390400
transform 1 0 29008 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_250
timestamp 1669390400
transform 1 0 29344 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_252
timestamp 1669390400
transform 1 0 29568 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_255
timestamp 1669390400
transform 1 0 29904 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_308
timestamp 1669390400
transform 1 0 35840 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_316
timestamp 1669390400
transform 1 0 36736 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_318
timestamp 1669390400
transform 1 0 36960 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_321
timestamp 1669390400
transform 1 0 37296 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_324
timestamp 1669390400
transform 1 0 37632 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_328
timestamp 1669390400
transform 1 0 38080 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_338
timestamp 1669390400
transform 1 0 39200 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_342
timestamp 1669390400
transform 1 0 39648 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_346
timestamp 1669390400
transform 1 0 40096 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_355
timestamp 1669390400
transform 1 0 41104 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_369
timestamp 1669390400
transform 1 0 42672 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_389
timestamp 1669390400
transform 1 0 44912 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_392
timestamp 1669390400
transform 1 0 45248 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_401
timestamp 1669390400
transform 1 0 46256 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_409
timestamp 1669390400
transform 1 0 47152 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_422
timestamp 1669390400
transform 1 0 48608 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_56_426
timestamp 1669390400
transform 1 0 49056 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_442
timestamp 1669390400
transform 1 0 50848 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_446
timestamp 1669390400
transform 1 0 51296 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_456
timestamp 1669390400
transform 1 0 52416 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_460
timestamp 1669390400
transform 1 0 52864 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_463
timestamp 1669390400
transform 1 0 53200 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_471
timestamp 1669390400
transform 1 0 54096 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_473
timestamp 1669390400
transform 1 0 54320 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_487
timestamp 1669390400
transform 1 0 55888 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_56_497
timestamp 1669390400
transform 1 0 57008 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_2
timestamp 1669390400
transform 1 0 1568 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_4
timestamp 1669390400
transform 1 0 1792 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_7
timestamp 1669390400
transform 1 0 2128 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_11
timestamp 1669390400
transform 1 0 2576 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_15
timestamp 1669390400
transform 1 0 3024 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_25
timestamp 1669390400
transform 1 0 4144 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_29
timestamp 1669390400
transform 1 0 4592 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_70
timestamp 1669390400
transform 1 0 9184 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_73
timestamp 1669390400
transform 1 0 9520 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_84
timestamp 1669390400
transform 1 0 10752 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_88
timestamp 1669390400
transform 1 0 11200 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_91
timestamp 1669390400
transform 1 0 11536 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_95
timestamp 1669390400
transform 1 0 11984 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_99
timestamp 1669390400
transform 1 0 12432 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_109
timestamp 1669390400
transform 1 0 13552 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_122
timestamp 1669390400
transform 1 0 15008 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_124
timestamp 1669390400
transform 1 0 15232 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_134
timestamp 1669390400
transform 1 0 16352 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_138
timestamp 1669390400
transform 1 0 16800 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_141
timestamp 1669390400
transform 1 0 17136 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_144
timestamp 1669390400
transform 1 0 17472 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_155
timestamp 1669390400
transform 1 0 18704 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_161
timestamp 1669390400
transform 1 0 19376 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_186
timestamp 1669390400
transform 1 0 22176 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_192
timestamp 1669390400
transform 1 0 22848 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_204
timestamp 1669390400
transform 1 0 24192 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_208
timestamp 1669390400
transform 1 0 24640 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_212
timestamp 1669390400
transform 1 0 25088 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_215
timestamp 1669390400
transform 1 0 25424 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_217
timestamp 1669390400
transform 1 0 25648 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_220
timestamp 1669390400
transform 1 0 25984 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_224
timestamp 1669390400
transform 1 0 26432 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_227
timestamp 1669390400
transform 1 0 26768 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_280
timestamp 1669390400
transform 1 0 32704 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_286
timestamp 1669390400
transform 1 0 33376 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_299
timestamp 1669390400
transform 1 0 34832 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_301
timestamp 1669390400
transform 1 0 35056 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_315
timestamp 1669390400
transform 1 0 36624 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_319
timestamp 1669390400
transform 1 0 37072 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_323
timestamp 1669390400
transform 1 0 37520 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_336
timestamp 1669390400
transform 1 0 38976 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_351
timestamp 1669390400
transform 1 0 40656 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_357
timestamp 1669390400
transform 1 0 41328 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_365
timestamp 1669390400
transform 1 0 42224 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_381
timestamp 1669390400
transform 1 0 44016 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_389
timestamp 1669390400
transform 1 0 44912 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_393
timestamp 1669390400
transform 1 0 45360 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_406
timestamp 1669390400
transform 1 0 46816 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_422
timestamp 1669390400
transform 1 0 48608 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_428
timestamp 1669390400
transform 1 0 49280 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_433
timestamp 1669390400
transform 1 0 49840 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_437
timestamp 1669390400
transform 1 0 50288 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_447
timestamp 1669390400
transform 1 0 51408 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_460
timestamp 1669390400
transform 1 0 52864 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_464
timestamp 1669390400
transform 1 0 53312 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_472
timestamp 1669390400
transform 1 0 54208 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_488
timestamp 1669390400
transform 1 0 56000 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_492
timestamp 1669390400
transform 1 0 56448 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_496
timestamp 1669390400
transform 1 0 56896 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_499
timestamp 1669390400
transform 1 0 57232 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_512
timestamp 1669390400
transform 1 0 58688 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_2
timestamp 1669390400
transform 1 0 1568 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_6
timestamp 1669390400
transform 1 0 2016 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_10
timestamp 1669390400
transform 1 0 2464 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_14
timestamp 1669390400
transform 1 0 2912 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_24
timestamp 1669390400
transform 1 0 4032 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_30
timestamp 1669390400
transform 1 0 4704 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_34
timestamp 1669390400
transform 1 0 5152 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_37
timestamp 1669390400
transform 1 0 5488 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_44
timestamp 1669390400
transform 1 0 6272 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_56
timestamp 1669390400
transform 1 0 7616 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_60
timestamp 1669390400
transform 1 0 8064 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_64
timestamp 1669390400
transform 1 0 8512 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_68
timestamp 1669390400
transform 1 0 8960 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_72
timestamp 1669390400
transform 1 0 9408 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_82
timestamp 1669390400
transform 1 0 10528 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_84
timestamp 1669390400
transform 1 0 10752 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_93
timestamp 1669390400
transform 1 0 11760 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_105
timestamp 1669390400
transform 1 0 13104 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_108
timestamp 1669390400
transform 1 0 13440 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_114
timestamp 1669390400
transform 1 0 14112 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_118
timestamp 1669390400
transform 1 0 14560 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_125
timestamp 1669390400
transform 1 0 15344 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_129
timestamp 1669390400
transform 1 0 15792 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_133
timestamp 1669390400
transform 1 0 16240 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_137
timestamp 1669390400
transform 1 0 16688 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_141
timestamp 1669390400
transform 1 0 17136 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_145
timestamp 1669390400
transform 1 0 17584 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_156
timestamp 1669390400
transform 1 0 18816 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_176
timestamp 1669390400
transform 1 0 21056 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_179
timestamp 1669390400
transform 1 0 21392 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_185
timestamp 1669390400
transform 1 0 22064 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_206
timestamp 1669390400
transform 1 0 24416 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_217
timestamp 1669390400
transform 1 0 25648 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_221
timestamp 1669390400
transform 1 0 26096 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_225
timestamp 1669390400
transform 1 0 26544 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_229
timestamp 1669390400
transform 1 0 26992 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_235
timestamp 1669390400
transform 1 0 27664 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_239
timestamp 1669390400
transform 1 0 28112 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_243
timestamp 1669390400
transform 1 0 28560 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_247
timestamp 1669390400
transform 1 0 29008 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_250
timestamp 1669390400
transform 1 0 29344 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_302
timestamp 1669390400
transform 1 0 35168 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_316
timestamp 1669390400
transform 1 0 36736 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_318
timestamp 1669390400
transform 1 0 36960 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_321
timestamp 1669390400
transform 1 0 37296 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_324
timestamp 1669390400
transform 1 0 37632 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_328
timestamp 1669390400
transform 1 0 38080 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_332
timestamp 1669390400
transform 1 0 38528 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_336
timestamp 1669390400
transform 1 0 38976 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_58_343
timestamp 1669390400
transform 1 0 39760 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_359
timestamp 1669390400
transform 1 0 41552 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_366
timestamp 1669390400
transform 1 0 42336 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_370
timestamp 1669390400
transform 1 0 42784 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_372
timestamp 1669390400
transform 1 0 43008 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_378
timestamp 1669390400
transform 1 0 43680 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_382
timestamp 1669390400
transform 1 0 44128 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_389
timestamp 1669390400
transform 1 0 44912 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_392
timestamp 1669390400
transform 1 0 45248 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_396
timestamp 1669390400
transform 1 0 45696 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_398
timestamp 1669390400
transform 1 0 45920 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_412
timestamp 1669390400
transform 1 0 47488 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_420
timestamp 1669390400
transform 1 0 48384 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_424
timestamp 1669390400
transform 1 0 48832 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_433
timestamp 1669390400
transform 1 0 49840 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_441
timestamp 1669390400
transform 1 0 50736 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_443
timestamp 1669390400
transform 1 0 50960 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_446
timestamp 1669390400
transform 1 0 51296 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_460
timestamp 1669390400
transform 1 0 52864 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_463
timestamp 1669390400
transform 1 0 53200 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_469
timestamp 1669390400
transform 1 0 53872 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_473
timestamp 1669390400
transform 1 0 54320 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_486
timestamp 1669390400
transform 1 0 55776 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_506
timestamp 1669390400
transform 1 0 58016 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_510
timestamp 1669390400
transform 1 0 58464 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_512
timestamp 1669390400
transform 1 0 58688 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_2
timestamp 1669390400
transform 1 0 1568 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_4
timestamp 1669390400
transform 1 0 1792 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_7
timestamp 1669390400
transform 1 0 2128 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_11
timestamp 1669390400
transform 1 0 2576 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_15
timestamp 1669390400
transform 1 0 3024 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_25
timestamp 1669390400
transform 1 0 4144 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_35
timestamp 1669390400
transform 1 0 5264 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_45
timestamp 1669390400
transform 1 0 6384 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_47
timestamp 1669390400
transform 1 0 6608 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_56
timestamp 1669390400
transform 1 0 7616 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_66
timestamp 1669390400
transform 1 0 8736 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_70
timestamp 1669390400
transform 1 0 9184 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_73
timestamp 1669390400
transform 1 0 9520 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_75
timestamp 1669390400
transform 1 0 9744 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_88
timestamp 1669390400
transform 1 0 11200 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_95
timestamp 1669390400
transform 1 0 11984 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_102
timestamp 1669390400
transform 1 0 12768 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_112
timestamp 1669390400
transform 1 0 13888 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_122
timestamp 1669390400
transform 1 0 15008 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_124
timestamp 1669390400
transform 1 0 15232 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_131
timestamp 1669390400
transform 1 0 16016 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_137
timestamp 1669390400
transform 1 0 16688 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_141
timestamp 1669390400
transform 1 0 17136 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_144
timestamp 1669390400
transform 1 0 17472 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_150
timestamp 1669390400
transform 1 0 18144 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_162
timestamp 1669390400
transform 1 0 19488 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_164
timestamp 1669390400
transform 1 0 19712 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_167
timestamp 1669390400
transform 1 0 20048 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_191
timestamp 1669390400
transform 1 0 22736 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_211
timestamp 1669390400
transform 1 0 24976 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_215
timestamp 1669390400
transform 1 0 25424 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_219
timestamp 1669390400
transform 1 0 25872 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_223
timestamp 1669390400
transform 1 0 26320 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_233
timestamp 1669390400
transform 1 0 27440 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_239
timestamp 1669390400
transform 1 0 28112 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_243
timestamp 1669390400
transform 1 0 28560 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_247
timestamp 1669390400
transform 1 0 29008 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_255
timestamp 1669390400
transform 1 0 29904 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_265
timestamp 1669390400
transform 1 0 31024 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_274
timestamp 1669390400
transform 1 0 32032 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_282
timestamp 1669390400
transform 1 0 32928 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_286
timestamp 1669390400
transform 1 0 33376 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_299
timestamp 1669390400
transform 1 0 34832 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_303
timestamp 1669390400
transform 1 0 35280 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_312
timestamp 1669390400
transform 1 0 36288 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_316
timestamp 1669390400
transform 1 0 36736 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_320
timestamp 1669390400
transform 1 0 37184 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_324
timestamp 1669390400
transform 1 0 37632 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_346
timestamp 1669390400
transform 1 0 40096 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_350
timestamp 1669390400
transform 1 0 40544 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_354
timestamp 1669390400
transform 1 0 40992 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_357
timestamp 1669390400
transform 1 0 41328 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_371
timestamp 1669390400
transform 1 0 42896 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_381
timestamp 1669390400
transform 1 0 44016 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_389
timestamp 1669390400
transform 1 0 44912 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_393
timestamp 1669390400
transform 1 0 45360 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_395
timestamp 1669390400
transform 1 0 45584 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_401
timestamp 1669390400
transform 1 0 46256 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_425
timestamp 1669390400
transform 1 0 48944 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_428
timestamp 1669390400
transform 1 0 49280 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_437
timestamp 1669390400
transform 1 0 50288 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_441
timestamp 1669390400
transform 1 0 50736 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_444
timestamp 1669390400
transform 1 0 51072 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_448
timestamp 1669390400
transform 1 0 51520 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_460
timestamp 1669390400
transform 1 0 52864 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_464
timestamp 1669390400
transform 1 0 53312 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_470
timestamp 1669390400
transform 1 0 53984 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_478
timestamp 1669390400
transform 1 0 54880 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_492
timestamp 1669390400
transform 1 0 56448 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_496
timestamp 1669390400
transform 1 0 56896 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_499
timestamp 1669390400
transform 1 0 57232 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_505
timestamp 1669390400
transform 1 0 57904 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_512
timestamp 1669390400
transform 1 0 58688 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_2
timestamp 1669390400
transform 1 0 1568 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_8
timestamp 1669390400
transform 1 0 2240 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_12
timestamp 1669390400
transform 1 0 2688 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_16
timestamp 1669390400
transform 1 0 3136 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_26
timestamp 1669390400
transform 1 0 4256 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_30
timestamp 1669390400
transform 1 0 4704 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_34
timestamp 1669390400
transform 1 0 5152 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_37
timestamp 1669390400
transform 1 0 5488 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_41
timestamp 1669390400
transform 1 0 5936 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_53
timestamp 1669390400
transform 1 0 7280 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_61
timestamp 1669390400
transform 1 0 8176 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_63
timestamp 1669390400
transform 1 0 8400 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_87
timestamp 1669390400
transform 1 0 11088 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_91
timestamp 1669390400
transform 1 0 11536 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_101
timestamp 1669390400
transform 1 0 12656 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_105
timestamp 1669390400
transform 1 0 13104 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_108
timestamp 1669390400
transform 1 0 13440 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_121
timestamp 1669390400
transform 1 0 14896 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_131
timestamp 1669390400
transform 1 0 16016 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_139
timestamp 1669390400
transform 1 0 16912 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_143
timestamp 1669390400
transform 1 0 17360 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_152
timestamp 1669390400
transform 1 0 18368 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_162
timestamp 1669390400
transform 1 0 19488 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_176
timestamp 1669390400
transform 1 0 21056 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_179
timestamp 1669390400
transform 1 0 21392 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_185
timestamp 1669390400
transform 1 0 22064 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_189
timestamp 1669390400
transform 1 0 22512 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_193
timestamp 1669390400
transform 1 0 22960 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_197
timestamp 1669390400
transform 1 0 23408 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_201
timestamp 1669390400
transform 1 0 23856 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_205
timestamp 1669390400
transform 1 0 24304 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_214
timestamp 1669390400
transform 1 0 25312 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_220
timestamp 1669390400
transform 1 0 25984 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_234
timestamp 1669390400
transform 1 0 27552 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_242
timestamp 1669390400
transform 1 0 28448 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_244
timestamp 1669390400
transform 1 0 28672 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_247
timestamp 1669390400
transform 1 0 29008 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_250
timestamp 1669390400
transform 1 0 29344 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_263
timestamp 1669390400
transform 1 0 30800 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_270
timestamp 1669390400
transform 1 0 31584 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_272
timestamp 1669390400
transform 1 0 31808 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_275
timestamp 1669390400
transform 1 0 32144 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_279
timestamp 1669390400
transform 1 0 32592 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_281
timestamp 1669390400
transform 1 0 32816 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_288
timestamp 1669390400
transform 1 0 33600 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_292
timestamp 1669390400
transform 1 0 34048 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_296
timestamp 1669390400
transform 1 0 34496 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_300
timestamp 1669390400
transform 1 0 34944 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_304
timestamp 1669390400
transform 1 0 35392 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_318
timestamp 1669390400
transform 1 0 36960 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_321
timestamp 1669390400
transform 1 0 37296 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_334
timestamp 1669390400
transform 1 0 38752 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_344
timestamp 1669390400
transform 1 0 39872 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_352
timestamp 1669390400
transform 1 0 40768 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_356
timestamp 1669390400
transform 1 0 41216 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_364
timestamp 1669390400
transform 1 0 42112 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_379
timestamp 1669390400
transform 1 0 43792 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_387
timestamp 1669390400
transform 1 0 44688 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_389
timestamp 1669390400
transform 1 0 44912 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_392
timestamp 1669390400
transform 1 0 45248 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_396
timestamp 1669390400
transform 1 0 45696 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_403
timestamp 1669390400
transform 1 0 46480 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_410
timestamp 1669390400
transform 1 0 47264 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_418
timestamp 1669390400
transform 1 0 48160 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_442
timestamp 1669390400
transform 1 0 50848 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_452
timestamp 1669390400
transform 1 0 51968 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_460
timestamp 1669390400
transform 1 0 52864 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_463
timestamp 1669390400
transform 1 0 53200 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_465
timestamp 1669390400
transform 1 0 53424 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_468
timestamp 1669390400
transform 1 0 53760 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_480
timestamp 1669390400
transform 1 0 55104 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_484
timestamp 1669390400
transform 1 0 55552 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_493
timestamp 1669390400
transform 1 0 56560 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_503
timestamp 1669390400
transform 1 0 57680 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_510
timestamp 1669390400
transform 1 0 58464 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_512
timestamp 1669390400
transform 1 0 58688 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_2
timestamp 1669390400
transform 1 0 1568 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_6
timestamp 1669390400
transform 1 0 2016 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_10
timestamp 1669390400
transform 1 0 2464 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_14
timestamp 1669390400
transform 1 0 2912 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_18
timestamp 1669390400
transform 1 0 3360 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_22
timestamp 1669390400
transform 1 0 3808 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_26
timestamp 1669390400
transform 1 0 4256 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_30
timestamp 1669390400
transform 1 0 4704 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_33
timestamp 1669390400
transform 1 0 5040 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_37
timestamp 1669390400
transform 1 0 5488 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_41
timestamp 1669390400
transform 1 0 5936 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_51
timestamp 1669390400
transform 1 0 7056 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_61
timestamp 1669390400
transform 1 0 8176 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_70
timestamp 1669390400
transform 1 0 9184 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_73
timestamp 1669390400
transform 1 0 9520 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_97
timestamp 1669390400
transform 1 0 12208 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_101
timestamp 1669390400
transform 1 0 12656 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_121
timestamp 1669390400
transform 1 0 14896 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_135
timestamp 1669390400
transform 1 0 16464 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_141
timestamp 1669390400
transform 1 0 17136 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_144
timestamp 1669390400
transform 1 0 17472 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_146
timestamp 1669390400
transform 1 0 17696 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_149
timestamp 1669390400
transform 1 0 18032 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_158
timestamp 1669390400
transform 1 0 19040 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_172
timestamp 1669390400
transform 1 0 20608 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_176
timestamp 1669390400
transform 1 0 21056 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_179
timestamp 1669390400
transform 1 0 21392 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_183
timestamp 1669390400
transform 1 0 21840 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_187
timestamp 1669390400
transform 1 0 22288 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_191
timestamp 1669390400
transform 1 0 22736 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_200
timestamp 1669390400
transform 1 0 23744 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_212
timestamp 1669390400
transform 1 0 25088 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_215
timestamp 1669390400
transform 1 0 25424 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_217
timestamp 1669390400
transform 1 0 25648 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_228
timestamp 1669390400
transform 1 0 26880 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_242
timestamp 1669390400
transform 1 0 28448 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_246
timestamp 1669390400
transform 1 0 28896 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_253
timestamp 1669390400
transform 1 0 29680 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_268
timestamp 1669390400
transform 1 0 31360 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_283
timestamp 1669390400
transform 1 0 33040 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_286
timestamp 1669390400
transform 1 0 33376 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_299
timestamp 1669390400
transform 1 0 34832 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_307
timestamp 1669390400
transform 1 0 35728 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_309
timestamp 1669390400
transform 1 0 35952 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_318
timestamp 1669390400
transform 1 0 36960 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_326
timestamp 1669390400
transform 1 0 37856 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_342
timestamp 1669390400
transform 1 0 39648 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_346
timestamp 1669390400
transform 1 0 40096 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_354
timestamp 1669390400
transform 1 0 40992 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_357
timestamp 1669390400
transform 1 0 41328 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_361
timestamp 1669390400
transform 1 0 41776 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_368
timestamp 1669390400
transform 1 0 42560 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_383
timestamp 1669390400
transform 1 0 44240 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_387
timestamp 1669390400
transform 1 0 44688 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_392
timestamp 1669390400
transform 1 0 45248 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_417
timestamp 1669390400
transform 1 0 48048 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_425
timestamp 1669390400
transform 1 0 48944 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_61_428
timestamp 1669390400
transform 1 0 49280 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_444
timestamp 1669390400
transform 1 0 51072 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_61_457
timestamp 1669390400
transform 1 0 52528 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_473
timestamp 1669390400
transform 1 0 54320 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_477
timestamp 1669390400
transform 1 0 54768 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_487
timestamp 1669390400
transform 1 0 55888 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_491
timestamp 1669390400
transform 1 0 56336 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_495
timestamp 1669390400
transform 1 0 56784 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_499
timestamp 1669390400
transform 1 0 57232 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_503
timestamp 1669390400
transform 1 0 57680 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_507
timestamp 1669390400
transform 1 0 58128 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_511
timestamp 1669390400
transform 1 0 58576 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_2
timestamp 1669390400
transform 1 0 1568 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_5
timestamp 1669390400
transform 1 0 1904 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_9
timestamp 1669390400
transform 1 0 2352 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_13
timestamp 1669390400
transform 1 0 2800 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_17
timestamp 1669390400
transform 1 0 3248 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_21
timestamp 1669390400
transform 1 0 3696 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_24
timestamp 1669390400
transform 1 0 4032 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_28
timestamp 1669390400
transform 1 0 4480 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_32
timestamp 1669390400
transform 1 0 4928 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_34
timestamp 1669390400
transform 1 0 5152 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_37
timestamp 1669390400
transform 1 0 5488 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_40
timestamp 1669390400
transform 1 0 5824 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_44
timestamp 1669390400
transform 1 0 6272 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_48
timestamp 1669390400
transform 1 0 6720 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_52
timestamp 1669390400
transform 1 0 7168 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_58
timestamp 1669390400
transform 1 0 7840 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_62
timestamp 1669390400
transform 1 0 8288 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_66
timestamp 1669390400
transform 1 0 8736 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_70
timestamp 1669390400
transform 1 0 9184 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_74
timestamp 1669390400
transform 1 0 9632 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_76
timestamp 1669390400
transform 1 0 9856 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_94
timestamp 1669390400
transform 1 0 11872 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_98
timestamp 1669390400
transform 1 0 12320 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_101
timestamp 1669390400
transform 1 0 12656 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_105
timestamp 1669390400
transform 1 0 13104 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_108
timestamp 1669390400
transform 1 0 13440 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_110
timestamp 1669390400
transform 1 0 13664 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_113
timestamp 1669390400
transform 1 0 14000 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_117
timestamp 1669390400
transform 1 0 14448 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_124
timestamp 1669390400
transform 1 0 15232 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_144
timestamp 1669390400
transform 1 0 17472 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_164
timestamp 1669390400
transform 1 0 19712 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_168
timestamp 1669390400
transform 1 0 20160 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_172
timestamp 1669390400
transform 1 0 20608 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_176
timestamp 1669390400
transform 1 0 21056 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_179
timestamp 1669390400
transform 1 0 21392 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_182
timestamp 1669390400
transform 1 0 21728 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_186
timestamp 1669390400
transform 1 0 22176 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_198
timestamp 1669390400
transform 1 0 23520 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_208
timestamp 1669390400
transform 1 0 24640 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_216
timestamp 1669390400
transform 1 0 25536 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_218
timestamp 1669390400
transform 1 0 25760 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_221
timestamp 1669390400
transform 1 0 26096 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_225
timestamp 1669390400
transform 1 0 26544 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_235
timestamp 1669390400
transform 1 0 27664 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_239
timestamp 1669390400
transform 1 0 28112 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_243
timestamp 1669390400
transform 1 0 28560 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_247
timestamp 1669390400
transform 1 0 29008 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_250
timestamp 1669390400
transform 1 0 29344 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_263
timestamp 1669390400
transform 1 0 30800 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_267
timestamp 1669390400
transform 1 0 31248 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_271
timestamp 1669390400
transform 1 0 31696 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_273
timestamp 1669390400
transform 1 0 31920 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_276
timestamp 1669390400
transform 1 0 32256 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_303
timestamp 1669390400
transform 1 0 35280 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_321
timestamp 1669390400
transform 1 0 37296 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_337
timestamp 1669390400
transform 1 0 39088 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_339
timestamp 1669390400
transform 1 0 39312 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_353
timestamp 1669390400
transform 1 0 40880 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_357
timestamp 1669390400
transform 1 0 41328 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_389
timestamp 1669390400
transform 1 0 44912 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_392
timestamp 1669390400
transform 1 0 45248 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_396
timestamp 1669390400
transform 1 0 45696 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_405
timestamp 1669390400
transform 1 0 46704 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_437
timestamp 1669390400
transform 1 0 50288 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_453
timestamp 1669390400
transform 1 0 52080 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_460
timestamp 1669390400
transform 1 0 52864 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_463
timestamp 1669390400
transform 1 0 53200 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_476
timestamp 1669390400
transform 1 0 54656 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_508
timestamp 1669390400
transform 1 0 58240 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_512
timestamp 1669390400
transform 1 0 58688 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_2
timestamp 1669390400
transform 1 0 1568 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_5
timestamp 1669390400
transform 1 0 1904 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_9
timestamp 1669390400
transform 1 0 2352 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_13
timestamp 1669390400
transform 1 0 2800 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_17
timestamp 1669390400
transform 1 0 3248 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_21
timestamp 1669390400
transform 1 0 3696 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_23
timestamp 1669390400
transform 1 0 3920 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_26
timestamp 1669390400
transform 1 0 4256 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_30
timestamp 1669390400
transform 1 0 4704 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_34
timestamp 1669390400
transform 1 0 5152 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_38
timestamp 1669390400
transform 1 0 5600 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_42
timestamp 1669390400
transform 1 0 6048 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_46
timestamp 1669390400
transform 1 0 6496 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_50
timestamp 1669390400
transform 1 0 6944 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_54
timestamp 1669390400
transform 1 0 7392 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_58
timestamp 1669390400
transform 1 0 7840 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_62
timestamp 1669390400
transform 1 0 8288 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_66
timestamp 1669390400
transform 1 0 8736 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_70
timestamp 1669390400
transform 1 0 9184 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_73
timestamp 1669390400
transform 1 0 9520 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_75
timestamp 1669390400
transform 1 0 9744 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_78
timestamp 1669390400
transform 1 0 10080 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_82
timestamp 1669390400
transform 1 0 10528 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_84
timestamp 1669390400
transform 1 0 10752 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_87
timestamp 1669390400
transform 1 0 11088 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_91
timestamp 1669390400
transform 1 0 11536 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_95
timestamp 1669390400
transform 1 0 11984 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_99
timestamp 1669390400
transform 1 0 12432 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_103
timestamp 1669390400
transform 1 0 12880 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_107
timestamp 1669390400
transform 1 0 13328 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_111
timestamp 1669390400
transform 1 0 13776 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_114
timestamp 1669390400
transform 1 0 14112 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_118
timestamp 1669390400
transform 1 0 14560 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_122
timestamp 1669390400
transform 1 0 15008 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_126
timestamp 1669390400
transform 1 0 15456 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_130
timestamp 1669390400
transform 1 0 15904 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_133
timestamp 1669390400
transform 1 0 16240 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_137
timestamp 1669390400
transform 1 0 16688 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_141
timestamp 1669390400
transform 1 0 17136 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_144
timestamp 1669390400
transform 1 0 17472 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_154
timestamp 1669390400
transform 1 0 18592 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_156
timestamp 1669390400
transform 1 0 18816 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_159
timestamp 1669390400
transform 1 0 19152 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_163
timestamp 1669390400
transform 1 0 19600 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_167
timestamp 1669390400
transform 1 0 20048 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_175
timestamp 1669390400
transform 1 0 20944 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_181
timestamp 1669390400
transform 1 0 21616 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_192
timestamp 1669390400
transform 1 0 22848 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_204
timestamp 1669390400
transform 1 0 24192 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_212
timestamp 1669390400
transform 1 0 25088 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_215
timestamp 1669390400
transform 1 0 25424 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_219
timestamp 1669390400
transform 1 0 25872 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_231
timestamp 1669390400
transform 1 0 27216 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_235
timestamp 1669390400
transform 1 0 27664 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_239
timestamp 1669390400
transform 1 0 28112 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_243
timestamp 1669390400
transform 1 0 28560 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_249
timestamp 1669390400
transform 1 0 29232 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_260
timestamp 1669390400
transform 1 0 30464 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_276
timestamp 1669390400
transform 1 0 32256 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_286
timestamp 1669390400
transform 1 0 33376 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_292
timestamp 1669390400
transform 1 0 34048 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_332
timestamp 1669390400
transform 1 0 38528 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_336
timestamp 1669390400
transform 1 0 38976 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_346
timestamp 1669390400
transform 1 0 40096 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_350
timestamp 1669390400
transform 1 0 40544 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_354
timestamp 1669390400
transform 1 0 40992 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_357
timestamp 1669390400
transform 1 0 41328 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_365
timestamp 1669390400
transform 1 0 42224 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_367
timestamp 1669390400
transform 1 0 42448 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_63_376
timestamp 1669390400
transform 1 0 43456 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_408
timestamp 1669390400
transform 1 0 47040 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_412
timestamp 1669390400
transform 1 0 47488 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_416
timestamp 1669390400
transform 1 0 47936 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_424
timestamp 1669390400
transform 1 0 48832 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_428
timestamp 1669390400
transform 1 0 49280 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_442
timestamp 1669390400
transform 1 0 50848 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_458
timestamp 1669390400
transform 1 0 52640 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_460
timestamp 1669390400
transform 1 0 52864 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_473
timestamp 1669390400
transform 1 0 54320 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_489
timestamp 1669390400
transform 1 0 56112 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_499
timestamp 1669390400
transform 1 0 57232 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_507
timestamp 1669390400
transform 1 0 58128 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_511
timestamp 1669390400
transform 1 0 58576 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_2
timestamp 1669390400
transform 1 0 1568 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_4
timestamp 1669390400
transform 1 0 1792 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_7
timestamp 1669390400
transform 1 0 2128 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_11
timestamp 1669390400
transform 1 0 2576 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_15
timestamp 1669390400
transform 1 0 3024 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_19
timestamp 1669390400
transform 1 0 3472 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_23
timestamp 1669390400
transform 1 0 3920 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_27
timestamp 1669390400
transform 1 0 4368 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_31
timestamp 1669390400
transform 1 0 4816 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_34
timestamp 1669390400
transform 1 0 5152 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_37
timestamp 1669390400
transform 1 0 5488 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_40
timestamp 1669390400
transform 1 0 5824 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_44
timestamp 1669390400
transform 1 0 6272 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_48
timestamp 1669390400
transform 1 0 6720 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_52
timestamp 1669390400
transform 1 0 7168 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_56
timestamp 1669390400
transform 1 0 7616 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_60
timestamp 1669390400
transform 1 0 8064 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_64
timestamp 1669390400
transform 1 0 8512 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_68
timestamp 1669390400
transform 1 0 8960 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_72
timestamp 1669390400
transform 1 0 9408 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_76
timestamp 1669390400
transform 1 0 9856 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_80
timestamp 1669390400
transform 1 0 10304 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_84
timestamp 1669390400
transform 1 0 10752 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_87
timestamp 1669390400
transform 1 0 11088 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_91
timestamp 1669390400
transform 1 0 11536 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_105
timestamp 1669390400
transform 1 0 13104 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_108
timestamp 1669390400
transform 1 0 13440 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_115
timestamp 1669390400
transform 1 0 14224 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_122
timestamp 1669390400
transform 1 0 15008 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_126
timestamp 1669390400
transform 1 0 15456 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_139
timestamp 1669390400
transform 1 0 16912 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_143
timestamp 1669390400
transform 1 0 17360 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_147
timestamp 1669390400
transform 1 0 17808 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_151
timestamp 1669390400
transform 1 0 18256 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_155
timestamp 1669390400
transform 1 0 18704 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_167
timestamp 1669390400
transform 1 0 20048 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_175
timestamp 1669390400
transform 1 0 20944 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_179
timestamp 1669390400
transform 1 0 21392 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_185
timestamp 1669390400
transform 1 0 22064 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_196
timestamp 1669390400
transform 1 0 23296 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_207
timestamp 1669390400
transform 1 0 24528 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_211
timestamp 1669390400
transform 1 0 24976 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_215
timestamp 1669390400
transform 1 0 25424 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_219
timestamp 1669390400
transform 1 0 25872 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_221
timestamp 1669390400
transform 1 0 26096 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_224
timestamp 1669390400
transform 1 0 26432 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_228
timestamp 1669390400
transform 1 0 26880 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_235
timestamp 1669390400
transform 1 0 27664 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_239
timestamp 1669390400
transform 1 0 28112 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_247
timestamp 1669390400
transform 1 0 29008 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_250
timestamp 1669390400
transform 1 0 29344 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_64_259
timestamp 1669390400
transform 1 0 30352 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_275
timestamp 1669390400
transform 1 0 32144 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_283
timestamp 1669390400
transform 1 0 33040 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_289
timestamp 1669390400
transform 1 0 33712 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_297
timestamp 1669390400
transform 1 0 34608 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_299
timestamp 1669390400
transform 1 0 34832 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_305
timestamp 1669390400
transform 1 0 35504 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_315
timestamp 1669390400
transform 1 0 36624 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_64_321
timestamp 1669390400
transform 1 0 37296 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_337
timestamp 1669390400
transform 1 0 39088 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_351
timestamp 1669390400
transform 1 0 40656 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_364
timestamp 1669390400
transform 1 0 42112 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_389
timestamp 1669390400
transform 1 0 44912 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_392
timestamp 1669390400
transform 1 0 45248 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_408
timestamp 1669390400
transform 1 0 47040 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_412
timestamp 1669390400
transform 1 0 47488 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_414
timestamp 1669390400
transform 1 0 47712 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_422
timestamp 1669390400
transform 1 0 48608 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_424
timestamp 1669390400
transform 1 0 48832 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_430
timestamp 1669390400
transform 1 0 49504 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_438
timestamp 1669390400
transform 1 0 50400 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_442
timestamp 1669390400
transform 1 0 50848 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_456
timestamp 1669390400
transform 1 0 52416 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_460
timestamp 1669390400
transform 1 0 52864 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_463
timestamp 1669390400
transform 1 0 53200 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_476
timestamp 1669390400
transform 1 0 54656 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_508
timestamp 1669390400
transform 1 0 58240 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_512
timestamp 1669390400
transform 1 0 58688 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_2
timestamp 1669390400
transform 1 0 1568 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_5
timestamp 1669390400
transform 1 0 1904 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_9
timestamp 1669390400
transform 1 0 2352 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_13
timestamp 1669390400
transform 1 0 2800 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_17
timestamp 1669390400
transform 1 0 3248 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_21
timestamp 1669390400
transform 1 0 3696 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_25
timestamp 1669390400
transform 1 0 4144 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_29
timestamp 1669390400
transform 1 0 4592 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_33
timestamp 1669390400
transform 1 0 5040 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_37
timestamp 1669390400
transform 1 0 5488 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_41
timestamp 1669390400
transform 1 0 5936 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_43
timestamp 1669390400
transform 1 0 6160 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_46
timestamp 1669390400
transform 1 0 6496 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_50
timestamp 1669390400
transform 1 0 6944 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_54
timestamp 1669390400
transform 1 0 7392 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_58
timestamp 1669390400
transform 1 0 7840 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_62
timestamp 1669390400
transform 1 0 8288 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_66
timestamp 1669390400
transform 1 0 8736 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_70
timestamp 1669390400
transform 1 0 9184 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_73
timestamp 1669390400
transform 1 0 9520 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_76
timestamp 1669390400
transform 1 0 9856 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_80
timestamp 1669390400
transform 1 0 10304 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_84
timestamp 1669390400
transform 1 0 10752 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_88
timestamp 1669390400
transform 1 0 11200 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_92
timestamp 1669390400
transform 1 0 11648 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_96
timestamp 1669390400
transform 1 0 12096 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_100
timestamp 1669390400
transform 1 0 12544 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_108
timestamp 1669390400
transform 1 0 13440 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_116
timestamp 1669390400
transform 1 0 14336 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_141
timestamp 1669390400
transform 1 0 17136 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_144
timestamp 1669390400
transform 1 0 17472 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_147
timestamp 1669390400
transform 1 0 17808 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_151
timestamp 1669390400
transform 1 0 18256 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_155
timestamp 1669390400
transform 1 0 18704 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_169
timestamp 1669390400
transform 1 0 20272 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_173
timestamp 1669390400
transform 1 0 20720 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_175
timestamp 1669390400
transform 1 0 20944 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_178
timestamp 1669390400
transform 1 0 21280 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_182
timestamp 1669390400
transform 1 0 21728 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_185
timestamp 1669390400
transform 1 0 22064 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_189
timestamp 1669390400
transform 1 0 22512 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_193
timestamp 1669390400
transform 1 0 22960 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_197
timestamp 1669390400
transform 1 0 23408 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_201
timestamp 1669390400
transform 1 0 23856 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_204
timestamp 1669390400
transform 1 0 24192 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_208
timestamp 1669390400
transform 1 0 24640 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_212
timestamp 1669390400
transform 1 0 25088 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_215
timestamp 1669390400
transform 1 0 25424 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_218
timestamp 1669390400
transform 1 0 25760 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_220
timestamp 1669390400
transform 1 0 25984 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_223
timestamp 1669390400
transform 1 0 26320 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_235
timestamp 1669390400
transform 1 0 27664 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_249
timestamp 1669390400
transform 1 0 29232 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_265
timestamp 1669390400
transform 1 0 31024 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_269
timestamp 1669390400
transform 1 0 31472 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_283
timestamp 1669390400
transform 1 0 33040 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_286
timestamp 1669390400
transform 1 0 33376 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_291
timestamp 1669390400
transform 1 0 33936 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_299
timestamp 1669390400
transform 1 0 34832 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_301
timestamp 1669390400
transform 1 0 35056 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_308
timestamp 1669390400
transform 1 0 35840 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_65_316
timestamp 1669390400
transform 1 0 36736 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_332
timestamp 1669390400
transform 1 0 38528 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_336
timestamp 1669390400
transform 1 0 38976 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_344
timestamp 1669390400
transform 1 0 39872 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_352
timestamp 1669390400
transform 1 0 40768 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_354
timestamp 1669390400
transform 1 0 40992 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_357
timestamp 1669390400
transform 1 0 41328 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_364
timestamp 1669390400
transform 1 0 42112 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_368
timestamp 1669390400
transform 1 0 42560 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_65_375
timestamp 1669390400
transform 1 0 43344 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_391
timestamp 1669390400
transform 1 0 45136 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_395
timestamp 1669390400
transform 1 0 45584 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_397
timestamp 1669390400
transform 1 0 45808 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_403
timestamp 1669390400
transform 1 0 46480 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_407
timestamp 1669390400
transform 1 0 46928 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_414
timestamp 1669390400
transform 1 0 47712 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_425
timestamp 1669390400
transform 1 0 48944 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_428
timestamp 1669390400
transform 1 0 49280 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_441
timestamp 1669390400
transform 1 0 50736 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_451
timestamp 1669390400
transform 1 0 51856 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_453
timestamp 1669390400
transform 1 0 52080 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_459
timestamp 1669390400
transform 1 0 52752 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_469
timestamp 1669390400
transform 1 0 53872 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_65_475
timestamp 1669390400
transform 1 0 54544 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_491
timestamp 1669390400
transform 1 0 56336 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_495
timestamp 1669390400
transform 1 0 56784 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_499
timestamp 1669390400
transform 1 0 57232 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_507
timestamp 1669390400
transform 1 0 58128 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_511
timestamp 1669390400
transform 1 0 58576 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_2
timestamp 1669390400
transform 1 0 1568 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_5
timestamp 1669390400
transform 1 0 1904 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_9
timestamp 1669390400
transform 1 0 2352 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_13
timestamp 1669390400
transform 1 0 2800 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_17
timestamp 1669390400
transform 1 0 3248 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_21
timestamp 1669390400
transform 1 0 3696 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_25
timestamp 1669390400
transform 1 0 4144 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_29
timestamp 1669390400
transform 1 0 4592 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_33
timestamp 1669390400
transform 1 0 5040 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_37
timestamp 1669390400
transform 1 0 5488 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_39
timestamp 1669390400
transform 1 0 5712 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_42
timestamp 1669390400
transform 1 0 6048 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_46
timestamp 1669390400
transform 1 0 6496 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_50
timestamp 1669390400
transform 1 0 6944 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_54
timestamp 1669390400
transform 1 0 7392 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_58
timestamp 1669390400
transform 1 0 7840 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_62
timestamp 1669390400
transform 1 0 8288 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_66
timestamp 1669390400
transform 1 0 8736 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_70
timestamp 1669390400
transform 1 0 9184 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_74
timestamp 1669390400
transform 1 0 9632 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_76
timestamp 1669390400
transform 1 0 9856 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_79
timestamp 1669390400
transform 1 0 10192 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_83
timestamp 1669390400
transform 1 0 10640 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_87
timestamp 1669390400
transform 1 0 11088 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_91
timestamp 1669390400
transform 1 0 11536 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_105
timestamp 1669390400
transform 1 0 13104 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_108
timestamp 1669390400
transform 1 0 13440 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_116
timestamp 1669390400
transform 1 0 14336 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_120
timestamp 1669390400
transform 1 0 14784 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_122
timestamp 1669390400
transform 1 0 15008 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_125
timestamp 1669390400
transform 1 0 15344 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_129
timestamp 1669390400
transform 1 0 15792 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_133
timestamp 1669390400
transform 1 0 16240 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_141
timestamp 1669390400
transform 1 0 17136 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_145
timestamp 1669390400
transform 1 0 17584 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_149
timestamp 1669390400
transform 1 0 18032 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_153
timestamp 1669390400
transform 1 0 18480 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_160
timestamp 1669390400
transform 1 0 19264 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_174
timestamp 1669390400
transform 1 0 20832 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_176
timestamp 1669390400
transform 1 0 21056 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_179
timestamp 1669390400
transform 1 0 21392 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_181
timestamp 1669390400
transform 1 0 21616 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_184
timestamp 1669390400
transform 1 0 21952 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_188
timestamp 1669390400
transform 1 0 22400 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_198
timestamp 1669390400
transform 1 0 23520 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_202
timestamp 1669390400
transform 1 0 23968 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_206
timestamp 1669390400
transform 1 0 24416 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_210
timestamp 1669390400
transform 1 0 24864 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_226
timestamp 1669390400
transform 1 0 26656 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_240
timestamp 1669390400
transform 1 0 28224 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_244
timestamp 1669390400
transform 1 0 28672 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_250
timestamp 1669390400
transform 1 0 29344 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_252
timestamp 1669390400
transform 1 0 29568 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_257
timestamp 1669390400
transform 1 0 30128 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_273
timestamp 1669390400
transform 1 0 31920 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_282
timestamp 1669390400
transform 1 0 32928 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_296
timestamp 1669390400
transform 1 0 34496 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_300
timestamp 1669390400
transform 1 0 34944 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_314
timestamp 1669390400
transform 1 0 36512 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_318
timestamp 1669390400
transform 1 0 36960 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_321
timestamp 1669390400
transform 1 0 37296 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_330
timestamp 1669390400
transform 1 0 38304 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_337
timestamp 1669390400
transform 1 0 39088 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_345
timestamp 1669390400
transform 1 0 39984 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_359
timestamp 1669390400
transform 1 0 41552 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_363
timestamp 1669390400
transform 1 0 42000 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_377
timestamp 1669390400
transform 1 0 43568 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_385
timestamp 1669390400
transform 1 0 44464 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_389
timestamp 1669390400
transform 1 0 44912 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_392
timestamp 1669390400
transform 1 0 45248 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_400
timestamp 1669390400
transform 1 0 46144 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_402
timestamp 1669390400
transform 1 0 46368 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_405
timestamp 1669390400
transform 1 0 46704 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_418
timestamp 1669390400
transform 1 0 48160 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_422
timestamp 1669390400
transform 1 0 48608 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_424
timestamp 1669390400
transform 1 0 48832 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_66_427
timestamp 1669390400
transform 1 0 49168 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_459
timestamp 1669390400
transform 1 0 52752 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_463
timestamp 1669390400
transform 1 0 53200 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_465
timestamp 1669390400
transform 1 0 53424 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_472
timestamp 1669390400
transform 1 0 54208 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_66_476
timestamp 1669390400
transform 1 0 54656 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_508
timestamp 1669390400
transform 1 0 58240 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_512
timestamp 1669390400
transform 1 0 58688 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_2
timestamp 1669390400
transform 1 0 1568 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_6
timestamp 1669390400
transform 1 0 2016 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_10
timestamp 1669390400
transform 1 0 2464 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_14
timestamp 1669390400
transform 1 0 2912 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_18
timestamp 1669390400
transform 1 0 3360 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_22
timestamp 1669390400
transform 1 0 3808 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_26
timestamp 1669390400
transform 1 0 4256 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_30
timestamp 1669390400
transform 1 0 4704 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_34
timestamp 1669390400
transform 1 0 5152 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_38
timestamp 1669390400
transform 1 0 5600 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_42
timestamp 1669390400
transform 1 0 6048 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_46
timestamp 1669390400
transform 1 0 6496 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_50
timestamp 1669390400
transform 1 0 6944 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_54
timestamp 1669390400
transform 1 0 7392 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_58
timestamp 1669390400
transform 1 0 7840 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_62
timestamp 1669390400
transform 1 0 8288 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_66
timestamp 1669390400
transform 1 0 8736 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_70
timestamp 1669390400
transform 1 0 9184 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_73
timestamp 1669390400
transform 1 0 9520 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_79
timestamp 1669390400
transform 1 0 10192 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_83
timestamp 1669390400
transform 1 0 10640 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_90
timestamp 1669390400
transform 1 0 11424 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_104
timestamp 1669390400
transform 1 0 12992 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_106
timestamp 1669390400
transform 1 0 13216 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_118
timestamp 1669390400
transform 1 0 14560 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_122
timestamp 1669390400
transform 1 0 15008 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_126
timestamp 1669390400
transform 1 0 15456 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_130
timestamp 1669390400
transform 1 0 15904 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_133
timestamp 1669390400
transform 1 0 16240 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_137
timestamp 1669390400
transform 1 0 16688 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_141
timestamp 1669390400
transform 1 0 17136 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_144
timestamp 1669390400
transform 1 0 17472 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_147
timestamp 1669390400
transform 1 0 17808 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_151
timestamp 1669390400
transform 1 0 18256 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_153
timestamp 1669390400
transform 1 0 18480 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_156
timestamp 1669390400
transform 1 0 18816 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_164
timestamp 1669390400
transform 1 0 19712 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_170
timestamp 1669390400
transform 1 0 20384 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_174
timestamp 1669390400
transform 1 0 20832 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_177
timestamp 1669390400
transform 1 0 21168 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_181
timestamp 1669390400
transform 1 0 21616 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_193
timestamp 1669390400
transform 1 0 22960 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_197
timestamp 1669390400
transform 1 0 23408 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_206
timestamp 1669390400
transform 1 0 24416 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_210
timestamp 1669390400
transform 1 0 24864 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_212
timestamp 1669390400
transform 1 0 25088 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_215
timestamp 1669390400
transform 1 0 25424 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_218
timestamp 1669390400
transform 1 0 25760 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_230
timestamp 1669390400
transform 1 0 27104 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_234
timestamp 1669390400
transform 1 0 27552 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_238
timestamp 1669390400
transform 1 0 28000 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_242
timestamp 1669390400
transform 1 0 28448 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_250
timestamp 1669390400
transform 1 0 29344 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_254
timestamp 1669390400
transform 1 0 29792 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_256
timestamp 1669390400
transform 1 0 30016 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_259
timestamp 1669390400
transform 1 0 30352 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_263
timestamp 1669390400
transform 1 0 30800 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_265
timestamp 1669390400
transform 1 0 31024 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_270
timestamp 1669390400
transform 1 0 31584 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_274
timestamp 1669390400
transform 1 0 32032 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_282
timestamp 1669390400
transform 1 0 32928 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_286
timestamp 1669390400
transform 1 0 33376 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_294
timestamp 1669390400
transform 1 0 34272 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_298
timestamp 1669390400
transform 1 0 34720 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_300
timestamp 1669390400
transform 1 0 34944 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_303
timestamp 1669390400
transform 1 0 35280 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_307
timestamp 1669390400
transform 1 0 35728 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_323
timestamp 1669390400
transform 1 0 37520 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_327
timestamp 1669390400
transform 1 0 37968 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_330
timestamp 1669390400
transform 1 0 38304 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_334
timestamp 1669390400
transform 1 0 38752 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_346
timestamp 1669390400
transform 1 0 40096 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_350
timestamp 1669390400
transform 1 0 40544 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_354
timestamp 1669390400
transform 1 0 40992 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_357
timestamp 1669390400
transform 1 0 41328 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_365
timestamp 1669390400
transform 1 0 42224 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_369
timestamp 1669390400
transform 1 0 42672 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_372
timestamp 1669390400
transform 1 0 43008 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_376
timestamp 1669390400
transform 1 0 43456 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_390
timestamp 1669390400
transform 1 0 45024 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_398
timestamp 1669390400
transform 1 0 45920 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_410
timestamp 1669390400
transform 1 0 47264 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_420
timestamp 1669390400
transform 1 0 48384 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_424
timestamp 1669390400
transform 1 0 48832 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_428
timestamp 1669390400
transform 1 0 49280 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_441
timestamp 1669390400
transform 1 0 50736 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_447
timestamp 1669390400
transform 1 0 51408 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_457
timestamp 1669390400
transform 1 0 52528 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_459
timestamp 1669390400
transform 1 0 52752 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_462
timestamp 1669390400
transform 1 0 53088 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_466
timestamp 1669390400
transform 1 0 53536 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_472
timestamp 1669390400
transform 1 0 54208 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_476
timestamp 1669390400
transform 1 0 54656 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_492
timestamp 1669390400
transform 1 0 56448 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_496
timestamp 1669390400
transform 1 0 56896 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_499
timestamp 1669390400
transform 1 0 57232 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_507
timestamp 1669390400
transform 1 0 58128 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_511
timestamp 1669390400
transform 1 0 58576 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_2
timestamp 1669390400
transform 1 0 1568 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_6
timestamp 1669390400
transform 1 0 2016 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_10
timestamp 1669390400
transform 1 0 2464 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_14
timestamp 1669390400
transform 1 0 2912 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_20
timestamp 1669390400
transform 1 0 3584 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_24
timestamp 1669390400
transform 1 0 4032 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_28
timestamp 1669390400
transform 1 0 4480 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_32
timestamp 1669390400
transform 1 0 4928 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_34
timestamp 1669390400
transform 1 0 5152 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_37
timestamp 1669390400
transform 1 0 5488 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_43
timestamp 1669390400
transform 1 0 6160 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_47
timestamp 1669390400
transform 1 0 6608 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_51
timestamp 1669390400
transform 1 0 7056 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_55
timestamp 1669390400
transform 1 0 7504 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_59
timestamp 1669390400
transform 1 0 7952 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_63
timestamp 1669390400
transform 1 0 8400 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_65
timestamp 1669390400
transform 1 0 8624 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_68
timestamp 1669390400
transform 1 0 8960 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_72
timestamp 1669390400
transform 1 0 9408 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_76
timestamp 1669390400
transform 1 0 9856 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_80
timestamp 1669390400
transform 1 0 10304 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_84
timestamp 1669390400
transform 1 0 10752 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_88
timestamp 1669390400
transform 1 0 11200 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_92
timestamp 1669390400
transform 1 0 11648 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_96
timestamp 1669390400
transform 1 0 12096 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_105
timestamp 1669390400
transform 1 0 13104 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_108
timestamp 1669390400
transform 1 0 13440 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_111
timestamp 1669390400
transform 1 0 13776 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_115
timestamp 1669390400
transform 1 0 14224 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_119
timestamp 1669390400
transform 1 0 14672 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_123
timestamp 1669390400
transform 1 0 15120 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_139
timestamp 1669390400
transform 1 0 16912 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_151
timestamp 1669390400
transform 1 0 18256 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_155
timestamp 1669390400
transform 1 0 18704 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_162
timestamp 1669390400
transform 1 0 19488 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_166
timestamp 1669390400
transform 1 0 19936 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_170
timestamp 1669390400
transform 1 0 20384 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_174
timestamp 1669390400
transform 1 0 20832 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_176
timestamp 1669390400
transform 1 0 21056 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_179
timestamp 1669390400
transform 1 0 21392 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_193
timestamp 1669390400
transform 1 0 22960 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_205
timestamp 1669390400
transform 1 0 24304 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_215
timestamp 1669390400
transform 1 0 25424 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_219
timestamp 1669390400
transform 1 0 25872 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_223
timestamp 1669390400
transform 1 0 26320 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_227
timestamp 1669390400
transform 1 0 26768 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_68_231
timestamp 1669390400
transform 1 0 27216 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_239
timestamp 1669390400
transform 1 0 28112 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_247
timestamp 1669390400
transform 1 0 29008 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_250
timestamp 1669390400
transform 1 0 29344 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_263
timestamp 1669390400
transform 1 0 30800 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_273
timestamp 1669390400
transform 1 0 31920 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_277
timestamp 1669390400
transform 1 0 32368 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_68_281
timestamp 1669390400
transform 1 0 32816 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_289
timestamp 1669390400
transform 1 0 33712 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_293
timestamp 1669390400
transform 1 0 34160 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_295
timestamp 1669390400
transform 1 0 34384 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_300
timestamp 1669390400
transform 1 0 34944 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_304
timestamp 1669390400
transform 1 0 35392 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_317
timestamp 1669390400
transform 1 0 36848 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_321
timestamp 1669390400
transform 1 0 37296 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_323
timestamp 1669390400
transform 1 0 37520 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_326
timestamp 1669390400
transform 1 0 37856 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_342
timestamp 1669390400
transform 1 0 39648 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_352
timestamp 1669390400
transform 1 0 40768 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_68_356
timestamp 1669390400
transform 1 0 41216 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_364
timestamp 1669390400
transform 1 0 42112 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_370
timestamp 1669390400
transform 1 0 42784 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_372
timestamp 1669390400
transform 1 0 43008 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_68_381
timestamp 1669390400
transform 1 0 44016 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_389
timestamp 1669390400
transform 1 0 44912 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_392
timestamp 1669390400
transform 1 0 45248 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_396
timestamp 1669390400
transform 1 0 45696 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_411
timestamp 1669390400
transform 1 0 47376 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_68_423
timestamp 1669390400
transform 1 0 48720 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_431
timestamp 1669390400
transform 1 0 49616 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_441
timestamp 1669390400
transform 1 0 50736 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_460
timestamp 1669390400
transform 1 0 52864 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_463
timestamp 1669390400
transform 1 0 53200 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_479
timestamp 1669390400
transform 1 0 54992 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_68_483
timestamp 1669390400
transform 1 0 55440 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_68_499
timestamp 1669390400
transform 1 0 57232 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_507
timestamp 1669390400
transform 1 0 58128 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_511
timestamp 1669390400
transform 1 0 58576 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_2
timestamp 1669390400
transform 1 0 1568 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_8
timestamp 1669390400
transform 1 0 2240 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_14
timestamp 1669390400
transform 1 0 2912 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_18
timestamp 1669390400
transform 1 0 3360 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_22
timestamp 1669390400
transform 1 0 3808 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_26
timestamp 1669390400
transform 1 0 4256 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_30
timestamp 1669390400
transform 1 0 4704 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_34
timestamp 1669390400
transform 1 0 5152 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_38
timestamp 1669390400
transform 1 0 5600 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_42
timestamp 1669390400
transform 1 0 6048 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_46
timestamp 1669390400
transform 1 0 6496 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_50
timestamp 1669390400
transform 1 0 6944 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_54
timestamp 1669390400
transform 1 0 7392 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_58
timestamp 1669390400
transform 1 0 7840 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_62
timestamp 1669390400
transform 1 0 8288 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_66
timestamp 1669390400
transform 1 0 8736 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_70
timestamp 1669390400
transform 1 0 9184 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_73
timestamp 1669390400
transform 1 0 9520 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_75
timestamp 1669390400
transform 1 0 9744 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_78
timestamp 1669390400
transform 1 0 10080 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_82
timestamp 1669390400
transform 1 0 10528 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_86
timestamp 1669390400
transform 1 0 10976 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_90
timestamp 1669390400
transform 1 0 11424 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_96
timestamp 1669390400
transform 1 0 12096 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_100
timestamp 1669390400
transform 1 0 12544 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_104
timestamp 1669390400
transform 1 0 12992 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_118
timestamp 1669390400
transform 1 0 14560 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_120
timestamp 1669390400
transform 1 0 14784 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_123
timestamp 1669390400
transform 1 0 15120 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_127
timestamp 1669390400
transform 1 0 15568 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_131
timestamp 1669390400
transform 1 0 16016 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_138
timestamp 1669390400
transform 1 0 16800 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_144
timestamp 1669390400
transform 1 0 17472 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_147
timestamp 1669390400
transform 1 0 17808 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_149
timestamp 1669390400
transform 1 0 18032 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_152
timestamp 1669390400
transform 1 0 18368 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_162
timestamp 1669390400
transform 1 0 19488 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_172
timestamp 1669390400
transform 1 0 20608 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_174
timestamp 1669390400
transform 1 0 20832 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_177
timestamp 1669390400
transform 1 0 21168 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_181
timestamp 1669390400
transform 1 0 21616 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_191
timestamp 1669390400
transform 1 0 22736 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_201
timestamp 1669390400
transform 1 0 23856 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_205
timestamp 1669390400
transform 1 0 24304 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_209
timestamp 1669390400
transform 1 0 24752 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_215
timestamp 1669390400
transform 1 0 25424 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_218
timestamp 1669390400
transform 1 0 25760 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_222
timestamp 1669390400
transform 1 0 26208 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_230
timestamp 1669390400
transform 1 0 27104 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_234
timestamp 1669390400
transform 1 0 27552 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_240
timestamp 1669390400
transform 1 0 28224 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_246
timestamp 1669390400
transform 1 0 28896 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_255
timestamp 1669390400
transform 1 0 29904 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_269
timestamp 1669390400
transform 1 0 31472 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_281
timestamp 1669390400
transform 1 0 32816 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_283
timestamp 1669390400
transform 1 0 33040 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_286
timestamp 1669390400
transform 1 0 33376 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_292
timestamp 1669390400
transform 1 0 34048 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_294
timestamp 1669390400
transform 1 0 34272 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_303
timestamp 1669390400
transform 1 0 35280 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_307
timestamp 1669390400
transform 1 0 35728 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_309
timestamp 1669390400
transform 1 0 35952 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_316
timestamp 1669390400
transform 1 0 36736 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_320
timestamp 1669390400
transform 1 0 37184 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_324
timestamp 1669390400
transform 1 0 37632 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_335
timestamp 1669390400
transform 1 0 38864 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_345
timestamp 1669390400
transform 1 0 39984 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_351
timestamp 1669390400
transform 1 0 40656 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_357
timestamp 1669390400
transform 1 0 41328 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_366
timestamp 1669390400
transform 1 0 42336 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_378
timestamp 1669390400
transform 1 0 43680 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_388
timestamp 1669390400
transform 1 0 44800 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_392
timestamp 1669390400
transform 1 0 45248 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_396
timestamp 1669390400
transform 1 0 45696 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_408
timestamp 1669390400
transform 1 0 47040 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_418
timestamp 1669390400
transform 1 0 48160 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_428
timestamp 1669390400
transform 1 0 49280 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_432
timestamp 1669390400
transform 1 0 49728 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_434
timestamp 1669390400
transform 1 0 49952 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_441
timestamp 1669390400
transform 1 0 50736 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_443
timestamp 1669390400
transform 1 0 50960 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_448
timestamp 1669390400
transform 1 0 51520 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_458
timestamp 1669390400
transform 1 0 52640 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_464
timestamp 1669390400
transform 1 0 53312 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_468
timestamp 1669390400
transform 1 0 53760 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_69_472
timestamp 1669390400
transform 1 0 54208 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_488
timestamp 1669390400
transform 1 0 56000 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_496
timestamp 1669390400
transform 1 0 56896 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_499
timestamp 1669390400
transform 1 0 57232 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_507
timestamp 1669390400
transform 1 0 58128 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_511
timestamp 1669390400
transform 1 0 58576 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_2
timestamp 1669390400
transform 1 0 1568 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_6
timestamp 1669390400
transform 1 0 2016 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_8
timestamp 1669390400
transform 1 0 2240 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_11
timestamp 1669390400
transform 1 0 2576 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_15
timestamp 1669390400
transform 1 0 3024 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_19
timestamp 1669390400
transform 1 0 3472 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_25
timestamp 1669390400
transform 1 0 4144 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_29
timestamp 1669390400
transform 1 0 4592 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_31
timestamp 1669390400
transform 1 0 4816 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_34
timestamp 1669390400
transform 1 0 5152 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_37
timestamp 1669390400
transform 1 0 5488 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_39
timestamp 1669390400
transform 1 0 5712 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_42
timestamp 1669390400
transform 1 0 6048 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_46
timestamp 1669390400
transform 1 0 6496 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_50
timestamp 1669390400
transform 1 0 6944 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_54
timestamp 1669390400
transform 1 0 7392 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_58
timestamp 1669390400
transform 1 0 7840 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_62
timestamp 1669390400
transform 1 0 8288 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_66
timestamp 1669390400
transform 1 0 8736 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_70
timestamp 1669390400
transform 1 0 9184 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_74
timestamp 1669390400
transform 1 0 9632 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_78
timestamp 1669390400
transform 1 0 10080 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_82
timestamp 1669390400
transform 1 0 10528 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_86
timestamp 1669390400
transform 1 0 10976 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_90
timestamp 1669390400
transform 1 0 11424 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_94
timestamp 1669390400
transform 1 0 11872 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_98
timestamp 1669390400
transform 1 0 12320 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_105
timestamp 1669390400
transform 1 0 13104 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_108
timestamp 1669390400
transform 1 0 13440 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_121
timestamp 1669390400
transform 1 0 14896 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_128
timestamp 1669390400
transform 1 0 15680 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_138
timestamp 1669390400
transform 1 0 16800 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_152
timestamp 1669390400
transform 1 0 18368 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_154
timestamp 1669390400
transform 1 0 18592 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_167
timestamp 1669390400
transform 1 0 20048 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_169
timestamp 1669390400
transform 1 0 20272 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_172
timestamp 1669390400
transform 1 0 20608 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_176
timestamp 1669390400
transform 1 0 21056 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_179
timestamp 1669390400
transform 1 0 21392 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_181
timestamp 1669390400
transform 1 0 21616 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_194
timestamp 1669390400
transform 1 0 23072 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_202
timestamp 1669390400
transform 1 0 23968 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_204
timestamp 1669390400
transform 1 0 24192 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_211
timestamp 1669390400
transform 1 0 24976 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_225
timestamp 1669390400
transform 1 0 26544 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_235
timestamp 1669390400
transform 1 0 27664 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_239
timestamp 1669390400
transform 1 0 28112 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_247
timestamp 1669390400
transform 1 0 29008 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_250
timestamp 1669390400
transform 1 0 29344 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_262
timestamp 1669390400
transform 1 0 30688 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_279
timestamp 1669390400
transform 1 0 32592 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_289
timestamp 1669390400
transform 1 0 33712 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_293
timestamp 1669390400
transform 1 0 34160 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_302
timestamp 1669390400
transform 1 0 35168 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_318
timestamp 1669390400
transform 1 0 36960 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_321
timestamp 1669390400
transform 1 0 37296 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_327
timestamp 1669390400
transform 1 0 37968 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_331
timestamp 1669390400
transform 1 0 38416 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_342
timestamp 1669390400
transform 1 0 39648 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_354
timestamp 1669390400
transform 1 0 40992 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_358
timestamp 1669390400
transform 1 0 41440 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_360
timestamp 1669390400
transform 1 0 41664 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_378
timestamp 1669390400
transform 1 0 43680 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_380
timestamp 1669390400
transform 1 0 43904 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_389
timestamp 1669390400
transform 1 0 44912 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_392
timestamp 1669390400
transform 1 0 45248 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_395
timestamp 1669390400
transform 1 0 45584 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_397
timestamp 1669390400
transform 1 0 45808 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_406
timestamp 1669390400
transform 1 0 46816 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_70_414
timestamp 1669390400
transform 1 0 47712 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_430
timestamp 1669390400
transform 1 0 49504 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_442
timestamp 1669390400
transform 1 0 50848 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_70_450
timestamp 1669390400
transform 1 0 51744 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_458
timestamp 1669390400
transform 1 0 52640 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_460
timestamp 1669390400
transform 1 0 52864 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_70_463
timestamp 1669390400
transform 1 0 53200 0 1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_70_495
timestamp 1669390400
transform 1 0 56784 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_511
timestamp 1669390400
transform 1 0 58576 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_71_2
timestamp 1669390400
transform 1 0 1568 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_10
timestamp 1669390400
transform 1 0 2464 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_14
timestamp 1669390400
transform 1 0 2912 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_18
timestamp 1669390400
transform 1 0 3360 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_22
timestamp 1669390400
transform 1 0 3808 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_26
timestamp 1669390400
transform 1 0 4256 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_30
timestamp 1669390400
transform 1 0 4704 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_34
timestamp 1669390400
transform 1 0 5152 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_38
timestamp 1669390400
transform 1 0 5600 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_42
timestamp 1669390400
transform 1 0 6048 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_46
timestamp 1669390400
transform 1 0 6496 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_50
timestamp 1669390400
transform 1 0 6944 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_54
timestamp 1669390400
transform 1 0 7392 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_58
timestamp 1669390400
transform 1 0 7840 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_62
timestamp 1669390400
transform 1 0 8288 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_66
timestamp 1669390400
transform 1 0 8736 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_70
timestamp 1669390400
transform 1 0 9184 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_73
timestamp 1669390400
transform 1 0 9520 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_76
timestamp 1669390400
transform 1 0 9856 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_80
timestamp 1669390400
transform 1 0 10304 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_88
timestamp 1669390400
transform 1 0 11200 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_92
timestamp 1669390400
transform 1 0 11648 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_95
timestamp 1669390400
transform 1 0 11984 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_99
timestamp 1669390400
transform 1 0 12432 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_103
timestamp 1669390400
transform 1 0 12880 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_107
timestamp 1669390400
transform 1 0 13328 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_111
timestamp 1669390400
transform 1 0 13776 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_125
timestamp 1669390400
transform 1 0 15344 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_133
timestamp 1669390400
transform 1 0 16240 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_137
timestamp 1669390400
transform 1 0 16688 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_141
timestamp 1669390400
transform 1 0 17136 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_144
timestamp 1669390400
transform 1 0 17472 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_150
timestamp 1669390400
transform 1 0 18144 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_164
timestamp 1669390400
transform 1 0 19712 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_174
timestamp 1669390400
transform 1 0 20832 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_191
timestamp 1669390400
transform 1 0 22736 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_193
timestamp 1669390400
transform 1 0 22960 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_208
timestamp 1669390400
transform 1 0 24640 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_212
timestamp 1669390400
transform 1 0 25088 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_215
timestamp 1669390400
transform 1 0 25424 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_218
timestamp 1669390400
transform 1 0 25760 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_220
timestamp 1669390400
transform 1 0 25984 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_233
timestamp 1669390400
transform 1 0 27440 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_245
timestamp 1669390400
transform 1 0 28784 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_251
timestamp 1669390400
transform 1 0 29456 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_258
timestamp 1669390400
transform 1 0 30240 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_265
timestamp 1669390400
transform 1 0 31024 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_71_269
timestamp 1669390400
transform 1 0 31472 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_282
timestamp 1669390400
transform 1 0 32928 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_286
timestamp 1669390400
transform 1 0 33376 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_297
timestamp 1669390400
transform 1 0 34608 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_307
timestamp 1669390400
transform 1 0 35728 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_316
timestamp 1669390400
transform 1 0 36736 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_320
timestamp 1669390400
transform 1 0 37184 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_324
timestamp 1669390400
transform 1 0 37632 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_326
timestamp 1669390400
transform 1 0 37856 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_332
timestamp 1669390400
transform 1 0 38528 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_342
timestamp 1669390400
transform 1 0 39648 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_352
timestamp 1669390400
transform 1 0 40768 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_354
timestamp 1669390400
transform 1 0 40992 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_357
timestamp 1669390400
transform 1 0 41328 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_360
timestamp 1669390400
transform 1 0 41664 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_370
timestamp 1669390400
transform 1 0 42784 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_380
timestamp 1669390400
transform 1 0 43904 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_390
timestamp 1669390400
transform 1 0 45024 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_396
timestamp 1669390400
transform 1 0 45696 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_71_400
timestamp 1669390400
transform 1 0 46144 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_71_416
timestamp 1669390400
transform 1 0 47936 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_424
timestamp 1669390400
transform 1 0 48832 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_428
timestamp 1669390400
transform 1 0 49280 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_492
timestamp 1669390400
transform 1 0 56448 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_496
timestamp 1669390400
transform 1 0 56896 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_71_499
timestamp 1669390400
transform 1 0 57232 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_507
timestamp 1669390400
transform 1 0 58128 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_511
timestamp 1669390400
transform 1 0 58576 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_72_2
timestamp 1669390400
transform 1 0 1568 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_18
timestamp 1669390400
transform 1 0 3360 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_22
timestamp 1669390400
transform 1 0 3808 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_26
timestamp 1669390400
transform 1 0 4256 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_30
timestamp 1669390400
transform 1 0 4704 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_34
timestamp 1669390400
transform 1 0 5152 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_37
timestamp 1669390400
transform 1 0 5488 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_41
timestamp 1669390400
transform 1 0 5936 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_45
timestamp 1669390400
transform 1 0 6384 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_49
timestamp 1669390400
transform 1 0 6832 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_53
timestamp 1669390400
transform 1 0 7280 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_57
timestamp 1669390400
transform 1 0 7728 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_61
timestamp 1669390400
transform 1 0 8176 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_65
timestamp 1669390400
transform 1 0 8624 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_69
timestamp 1669390400
transform 1 0 9072 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_72
timestamp 1669390400
transform 1 0 9408 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_76
timestamp 1669390400
transform 1 0 9856 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_78
timestamp 1669390400
transform 1 0 10080 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_93
timestamp 1669390400
transform 1 0 11760 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_99
timestamp 1669390400
transform 1 0 12432 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_101
timestamp 1669390400
transform 1 0 12656 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_104
timestamp 1669390400
transform 1 0 12992 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_107
timestamp 1669390400
transform 1 0 13328 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_110
timestamp 1669390400
transform 1 0 13664 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_114
timestamp 1669390400
transform 1 0 14112 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_124
timestamp 1669390400
transform 1 0 15232 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_126
timestamp 1669390400
transform 1 0 15456 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_129
timestamp 1669390400
transform 1 0 15792 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_133
timestamp 1669390400
transform 1 0 16240 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_137
timestamp 1669390400
transform 1 0 16688 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_139
timestamp 1669390400
transform 1 0 16912 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_142
timestamp 1669390400
transform 1 0 17248 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_146
timestamp 1669390400
transform 1 0 17696 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_150
timestamp 1669390400
transform 1 0 18144 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_156
timestamp 1669390400
transform 1 0 18816 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_160
timestamp 1669390400
transform 1 0 19264 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_162
timestamp 1669390400
transform 1 0 19488 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_165
timestamp 1669390400
transform 1 0 19824 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_169
timestamp 1669390400
transform 1 0 20272 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_173
timestamp 1669390400
transform 1 0 20720 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_177
timestamp 1669390400
transform 1 0 21168 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_180
timestamp 1669390400
transform 1 0 21504 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_184
timestamp 1669390400
transform 1 0 21952 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_188
timestamp 1669390400
transform 1 0 22400 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_201
timestamp 1669390400
transform 1 0 23856 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_205
timestamp 1669390400
transform 1 0 24304 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_209
timestamp 1669390400
transform 1 0 24752 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_212
timestamp 1669390400
transform 1 0 25088 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_72_215
timestamp 1669390400
transform 1 0 25424 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_223
timestamp 1669390400
transform 1 0 26320 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_72_231
timestamp 1669390400
transform 1 0 27216 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_239
timestamp 1669390400
transform 1 0 28112 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_243
timestamp 1669390400
transform 1 0 28560 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_247
timestamp 1669390400
transform 1 0 29008 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_251
timestamp 1669390400
transform 1 0 29456 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_253
timestamp 1669390400
transform 1 0 29680 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_256
timestamp 1669390400
transform 1 0 30016 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_72_272
timestamp 1669390400
transform 1 0 31808 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_282
timestamp 1669390400
transform 1 0 32928 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_285
timestamp 1669390400
transform 1 0 33264 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_293
timestamp 1669390400
transform 1 0 34160 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_299
timestamp 1669390400
transform 1 0 34832 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_303
timestamp 1669390400
transform 1 0 35280 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_72_306
timestamp 1669390400
transform 1 0 35616 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_314
timestamp 1669390400
transform 1 0 36512 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_72_317
timestamp 1669390400
transform 1 0 36848 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_349
timestamp 1669390400
transform 1 0 40432 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_72_352
timestamp 1669390400
transform 1 0 40768 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_368
timestamp 1669390400
transform 1 0 42560 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_372
timestamp 1669390400
transform 1 0 43008 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_376
timestamp 1669390400
transform 1 0 43456 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_381
timestamp 1669390400
transform 1 0 44016 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_387
timestamp 1669390400
transform 1 0 44688 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_72_390
timestamp 1669390400
transform 1 0 45024 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_72_406
timestamp 1669390400
transform 1 0 46816 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_414
timestamp 1669390400
transform 1 0 47712 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_418
timestamp 1669390400
transform 1 0 48160 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_72_422
timestamp 1669390400
transform 1 0 48608 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_430
timestamp 1669390400
transform 1 0 49504 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_432
timestamp 1669390400
transform 1 0 49728 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_435
timestamp 1669390400
transform 1 0 50064 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_451
timestamp 1669390400
transform 1 0 51856 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_72_457
timestamp 1669390400
transform 1 0 52528 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_489
timestamp 1669390400
transform 1 0 56112 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_72_492
timestamp 1669390400
transform 1 0 56448 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_508
timestamp 1669390400
transform 1 0 58240 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_512
timestamp 1669390400
transform 1 0 58688 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1669390400
transform -1 0 59024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1669390400
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1669390400
transform -1 0 59024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1669390400
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1669390400
transform -1 0 59024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1669390400
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1669390400
transform -1 0 59024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1669390400
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1669390400
transform -1 0 59024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1669390400
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1669390400
transform -1 0 59024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1669390400
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1669390400
transform -1 0 59024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1669390400
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1669390400
transform -1 0 59024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1669390400
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1669390400
transform -1 0 59024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1669390400
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1669390400
transform -1 0 59024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1669390400
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1669390400
transform -1 0 59024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1669390400
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1669390400
transform -1 0 59024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1669390400
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1669390400
transform -1 0 59024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1669390400
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1669390400
transform -1 0 59024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1669390400
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1669390400
transform -1 0 59024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1669390400
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1669390400
transform -1 0 59024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1669390400
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1669390400
transform -1 0 59024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1669390400
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1669390400
transform -1 0 59024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1669390400
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1669390400
transform -1 0 59024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1669390400
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1669390400
transform -1 0 59024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1669390400
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1669390400
transform -1 0 59024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1669390400
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1669390400
transform -1 0 59024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1669390400
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1669390400
transform -1 0 59024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1669390400
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1669390400
transform -1 0 59024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1669390400
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1669390400
transform -1 0 59024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1669390400
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1669390400
transform -1 0 59024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1669390400
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1669390400
transform -1 0 59024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1669390400
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1669390400
transform -1 0 59024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1669390400
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1669390400
transform -1 0 59024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1669390400
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1669390400
transform -1 0 59024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1669390400
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1669390400
transform -1 0 59024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1669390400
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1669390400
transform -1 0 59024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1669390400
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1669390400
transform -1 0 59024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1669390400
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1669390400
transform -1 0 59024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1669390400
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1669390400
transform -1 0 59024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1669390400
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1669390400
transform -1 0 59024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1669390400
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1669390400
transform -1 0 59024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1669390400
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1669390400
transform -1 0 59024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1669390400
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1669390400
transform -1 0 59024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1669390400
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1669390400
transform -1 0 59024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1669390400
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1669390400
transform -1 0 59024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1669390400
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1669390400
transform -1 0 59024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1669390400
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1669390400
transform -1 0 59024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_86
timestamp 1669390400
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_87
timestamp 1669390400
transform -1 0 59024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_88
timestamp 1669390400
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_89
timestamp 1669390400
transform -1 0 59024 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_90
timestamp 1669390400
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_91
timestamp 1669390400
transform -1 0 59024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_92
timestamp 1669390400
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_93
timestamp 1669390400
transform -1 0 59024 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_94
timestamp 1669390400
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_95
timestamp 1669390400
transform -1 0 59024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_96
timestamp 1669390400
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_97
timestamp 1669390400
transform -1 0 59024 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_98
timestamp 1669390400
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_99
timestamp 1669390400
transform -1 0 59024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_100
timestamp 1669390400
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_101
timestamp 1669390400
transform -1 0 59024 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_102
timestamp 1669390400
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_103
timestamp 1669390400
transform -1 0 59024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_104
timestamp 1669390400
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_105
timestamp 1669390400
transform -1 0 59024 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_106
timestamp 1669390400
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_107
timestamp 1669390400
transform -1 0 59024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_108
timestamp 1669390400
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_109
timestamp 1669390400
transform -1 0 59024 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_110
timestamp 1669390400
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_111
timestamp 1669390400
transform -1 0 59024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_112
timestamp 1669390400
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_113
timestamp 1669390400
transform -1 0 59024 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_114
timestamp 1669390400
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_115
timestamp 1669390400
transform -1 0 59024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_116
timestamp 1669390400
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_117
timestamp 1669390400
transform -1 0 59024 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_118
timestamp 1669390400
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_119
timestamp 1669390400
transform -1 0 59024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_120
timestamp 1669390400
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_121
timestamp 1669390400
transform -1 0 59024 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_122
timestamp 1669390400
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_123
timestamp 1669390400
transform -1 0 59024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_124
timestamp 1669390400
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_125
timestamp 1669390400
transform -1 0 59024 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_126
timestamp 1669390400
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_127
timestamp 1669390400
transform -1 0 59024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_128
timestamp 1669390400
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_129
timestamp 1669390400
transform -1 0 59024 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_130
timestamp 1669390400
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_131
timestamp 1669390400
transform -1 0 59024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_132
timestamp 1669390400
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_133
timestamp 1669390400
transform -1 0 59024 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_134
timestamp 1669390400
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_135
timestamp 1669390400
transform -1 0 59024 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_136
timestamp 1669390400
transform 1 0 1344 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_137
timestamp 1669390400
transform -1 0 59024 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_138
timestamp 1669390400
transform 1 0 1344 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_139
timestamp 1669390400
transform -1 0 59024 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_140
timestamp 1669390400
transform 1 0 1344 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_141
timestamp 1669390400
transform -1 0 59024 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_142
timestamp 1669390400
transform 1 0 1344 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_143
timestamp 1669390400
transform -1 0 59024 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_144
timestamp 1669390400
transform 1 0 1344 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_145
timestamp 1669390400
transform -1 0 59024 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_146 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_147
timestamp 1669390400
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_148
timestamp 1669390400
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_149
timestamp 1669390400
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_150
timestamp 1669390400
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_151
timestamp 1669390400
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_152
timestamp 1669390400
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_153
timestamp 1669390400
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_154
timestamp 1669390400
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_155
timestamp 1669390400
transform 1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_156
timestamp 1669390400
transform 1 0 44464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_157
timestamp 1669390400
transform 1 0 48384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_158
timestamp 1669390400
transform 1 0 52304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_159
timestamp 1669390400
transform 1 0 56224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_160
timestamp 1669390400
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_161
timestamp 1669390400
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_162
timestamp 1669390400
transform 1 0 25200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_163
timestamp 1669390400
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_164
timestamp 1669390400
transform 1 0 41104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_165
timestamp 1669390400
transform 1 0 49056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_166
timestamp 1669390400
transform 1 0 57008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_167
timestamp 1669390400
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_168
timestamp 1669390400
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_169
timestamp 1669390400
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_170
timestamp 1669390400
transform 1 0 29120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_171
timestamp 1669390400
transform 1 0 37072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_172
timestamp 1669390400
transform 1 0 45024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_173
timestamp 1669390400
transform 1 0 52976 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_174
timestamp 1669390400
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_175
timestamp 1669390400
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_176
timestamp 1669390400
transform 1 0 25200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_177
timestamp 1669390400
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_178
timestamp 1669390400
transform 1 0 41104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_179
timestamp 1669390400
transform 1 0 49056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_180
timestamp 1669390400
transform 1 0 57008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_181
timestamp 1669390400
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_182
timestamp 1669390400
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_183
timestamp 1669390400
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_184
timestamp 1669390400
transform 1 0 29120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_185
timestamp 1669390400
transform 1 0 37072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_186
timestamp 1669390400
transform 1 0 45024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_187
timestamp 1669390400
transform 1 0 52976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188
timestamp 1669390400
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1669390400
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1669390400
transform 1 0 25200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1669390400
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1669390400
transform 1 0 41104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1669390400
transform 1 0 49056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1669390400
transform 1 0 57008 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1669390400
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1669390400
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1669390400
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1669390400
transform 1 0 29120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1669390400
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1669390400
transform 1 0 45024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1669390400
transform 1 0 52976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1669390400
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1669390400
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1669390400
transform 1 0 25200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1669390400
transform 1 0 33152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1669390400
transform 1 0 41104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1669390400
transform 1 0 49056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1669390400
transform 1 0 57008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1669390400
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1669390400
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1669390400
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1669390400
transform 1 0 29120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1669390400
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1669390400
transform 1 0 45024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1669390400
transform 1 0 52976 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1669390400
transform 1 0 9296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1669390400
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1669390400
transform 1 0 25200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1669390400
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1669390400
transform 1 0 41104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1669390400
transform 1 0 49056 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1669390400
transform 1 0 57008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1669390400
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1669390400
transform 1 0 13216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1669390400
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1669390400
transform 1 0 29120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1669390400
transform 1 0 37072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1669390400
transform 1 0 45024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1669390400
transform 1 0 52976 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1669390400
transform 1 0 9296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1669390400
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1669390400
transform 1 0 25200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1669390400
transform 1 0 33152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1669390400
transform 1 0 41104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1669390400
transform 1 0 49056 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1669390400
transform 1 0 57008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1669390400
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1669390400
transform 1 0 13216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1669390400
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1669390400
transform 1 0 29120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1669390400
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1669390400
transform 1 0 45024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1669390400
transform 1 0 52976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1669390400
transform 1 0 9296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1669390400
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1669390400
transform 1 0 25200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1669390400
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1669390400
transform 1 0 41104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1669390400
transform 1 0 49056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1669390400
transform 1 0 57008 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1669390400
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1669390400
transform 1 0 13216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1669390400
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1669390400
transform 1 0 29120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1669390400
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1669390400
transform 1 0 45024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1669390400
transform 1 0 52976 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1669390400
transform 1 0 9296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1669390400
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1669390400
transform 1 0 25200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1669390400
transform 1 0 33152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1669390400
transform 1 0 41104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1669390400
transform 1 0 49056 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1669390400
transform 1 0 57008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1669390400
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1669390400
transform 1 0 13216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1669390400
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1669390400
transform 1 0 29120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1669390400
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1669390400
transform 1 0 45024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1669390400
transform 1 0 52976 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1669390400
transform 1 0 9296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1669390400
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1669390400
transform 1 0 25200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1669390400
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1669390400
transform 1 0 41104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1669390400
transform 1 0 49056 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1669390400
transform 1 0 57008 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1669390400
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1669390400
transform 1 0 13216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1669390400
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1669390400
transform 1 0 29120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1669390400
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1669390400
transform 1 0 45024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1669390400
transform 1 0 52976 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1669390400
transform 1 0 9296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1669390400
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_288
timestamp 1669390400
transform 1 0 25200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_289
timestamp 1669390400
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290
timestamp 1669390400
transform 1 0 41104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1669390400
transform 1 0 49056 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1669390400
transform 1 0 57008 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1669390400
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1669390400
transform 1 0 13216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1669390400
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1669390400
transform 1 0 29120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1669390400
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1669390400
transform 1 0 45024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1669390400
transform 1 0 52976 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1669390400
transform 1 0 9296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1669390400
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1669390400
transform 1 0 25200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1669390400
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1669390400
transform 1 0 41104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1669390400
transform 1 0 49056 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1669390400
transform 1 0 57008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1669390400
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1669390400
transform 1 0 13216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1669390400
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1669390400
transform 1 0 29120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1669390400
transform 1 0 37072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1669390400
transform 1 0 45024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1669390400
transform 1 0 52976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1669390400
transform 1 0 9296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1669390400
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1669390400
transform 1 0 25200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1669390400
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1669390400
transform 1 0 41104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1669390400
transform 1 0 49056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1669390400
transform 1 0 57008 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1669390400
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1669390400
transform 1 0 13216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1669390400
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1669390400
transform 1 0 29120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1669390400
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1669390400
transform 1 0 45024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1669390400
transform 1 0 52976 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1669390400
transform 1 0 9296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1669390400
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1669390400
transform 1 0 25200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1669390400
transform 1 0 33152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1669390400
transform 1 0 41104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1669390400
transform 1 0 49056 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1669390400
transform 1 0 57008 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1669390400
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1669390400
transform 1 0 13216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1669390400
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1669390400
transform 1 0 29120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1669390400
transform 1 0 37072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1669390400
transform 1 0 45024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1669390400
transform 1 0 52976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1669390400
transform 1 0 9296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1669390400
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1669390400
transform 1 0 25200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1669390400
transform 1 0 33152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_346
timestamp 1669390400
transform 1 0 41104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_347
timestamp 1669390400
transform 1 0 49056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_348
timestamp 1669390400
transform 1 0 57008 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_349
timestamp 1669390400
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_350
timestamp 1669390400
transform 1 0 13216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_351
timestamp 1669390400
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_352
timestamp 1669390400
transform 1 0 29120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_353
timestamp 1669390400
transform 1 0 37072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_354
timestamp 1669390400
transform 1 0 45024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_355
timestamp 1669390400
transform 1 0 52976 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_356
timestamp 1669390400
transform 1 0 9296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_357
timestamp 1669390400
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_358
timestamp 1669390400
transform 1 0 25200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_359
timestamp 1669390400
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_360
timestamp 1669390400
transform 1 0 41104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_361
timestamp 1669390400
transform 1 0 49056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_362
timestamp 1669390400
transform 1 0 57008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_363
timestamp 1669390400
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_364
timestamp 1669390400
transform 1 0 13216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_365
timestamp 1669390400
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_366
timestamp 1669390400
transform 1 0 29120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_367
timestamp 1669390400
transform 1 0 37072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_368
timestamp 1669390400
transform 1 0 45024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_369
timestamp 1669390400
transform 1 0 52976 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_370
timestamp 1669390400
transform 1 0 9296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_371
timestamp 1669390400
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_372
timestamp 1669390400
transform 1 0 25200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_373
timestamp 1669390400
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_374
timestamp 1669390400
transform 1 0 41104 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_375
timestamp 1669390400
transform 1 0 49056 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_376
timestamp 1669390400
transform 1 0 57008 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_377
timestamp 1669390400
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_378
timestamp 1669390400
transform 1 0 13216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_379
timestamp 1669390400
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_380
timestamp 1669390400
transform 1 0 29120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_381
timestamp 1669390400
transform 1 0 37072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_382
timestamp 1669390400
transform 1 0 45024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_383
timestamp 1669390400
transform 1 0 52976 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_384
timestamp 1669390400
transform 1 0 9296 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_385
timestamp 1669390400
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_386
timestamp 1669390400
transform 1 0 25200 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_387
timestamp 1669390400
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_388
timestamp 1669390400
transform 1 0 41104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_389
timestamp 1669390400
transform 1 0 49056 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_390
timestamp 1669390400
transform 1 0 57008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_391
timestamp 1669390400
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_392
timestamp 1669390400
transform 1 0 13216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_393
timestamp 1669390400
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_394
timestamp 1669390400
transform 1 0 29120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_395
timestamp 1669390400
transform 1 0 37072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_396
timestamp 1669390400
transform 1 0 45024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_397
timestamp 1669390400
transform 1 0 52976 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_398
timestamp 1669390400
transform 1 0 9296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_399
timestamp 1669390400
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_400
timestamp 1669390400
transform 1 0 25200 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_401
timestamp 1669390400
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_402
timestamp 1669390400
transform 1 0 41104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_403
timestamp 1669390400
transform 1 0 49056 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_404
timestamp 1669390400
transform 1 0 57008 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_405
timestamp 1669390400
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_406
timestamp 1669390400
transform 1 0 13216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_407
timestamp 1669390400
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_408
timestamp 1669390400
transform 1 0 29120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_409
timestamp 1669390400
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_410
timestamp 1669390400
transform 1 0 45024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_411
timestamp 1669390400
transform 1 0 52976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_412
timestamp 1669390400
transform 1 0 9296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_413
timestamp 1669390400
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_414
timestamp 1669390400
transform 1 0 25200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_415
timestamp 1669390400
transform 1 0 33152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_416
timestamp 1669390400
transform 1 0 41104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_417
timestamp 1669390400
transform 1 0 49056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_418
timestamp 1669390400
transform 1 0 57008 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_419
timestamp 1669390400
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_420
timestamp 1669390400
transform 1 0 13216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_421
timestamp 1669390400
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_422
timestamp 1669390400
transform 1 0 29120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_423
timestamp 1669390400
transform 1 0 37072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_424
timestamp 1669390400
transform 1 0 45024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_425
timestamp 1669390400
transform 1 0 52976 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_426
timestamp 1669390400
transform 1 0 9296 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_427
timestamp 1669390400
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_428
timestamp 1669390400
transform 1 0 25200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_429
timestamp 1669390400
transform 1 0 33152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_430
timestamp 1669390400
transform 1 0 41104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_431
timestamp 1669390400
transform 1 0 49056 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_432
timestamp 1669390400
transform 1 0 57008 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_433
timestamp 1669390400
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_434
timestamp 1669390400
transform 1 0 13216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_435
timestamp 1669390400
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_436
timestamp 1669390400
transform 1 0 29120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_437
timestamp 1669390400
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_438
timestamp 1669390400
transform 1 0 45024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_439
timestamp 1669390400
transform 1 0 52976 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_440
timestamp 1669390400
transform 1 0 9296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_441
timestamp 1669390400
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_442
timestamp 1669390400
transform 1 0 25200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_443
timestamp 1669390400
transform 1 0 33152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_444
timestamp 1669390400
transform 1 0 41104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_445
timestamp 1669390400
transform 1 0 49056 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_446
timestamp 1669390400
transform 1 0 57008 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_447
timestamp 1669390400
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_448
timestamp 1669390400
transform 1 0 13216 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_449
timestamp 1669390400
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_450
timestamp 1669390400
transform 1 0 29120 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_451
timestamp 1669390400
transform 1 0 37072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_452
timestamp 1669390400
transform 1 0 45024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_453
timestamp 1669390400
transform 1 0 52976 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_454
timestamp 1669390400
transform 1 0 9296 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_455
timestamp 1669390400
transform 1 0 17248 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_456
timestamp 1669390400
transform 1 0 25200 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_457
timestamp 1669390400
transform 1 0 33152 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_458
timestamp 1669390400
transform 1 0 41104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_459
timestamp 1669390400
transform 1 0 49056 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_460
timestamp 1669390400
transform 1 0 57008 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_461
timestamp 1669390400
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_462
timestamp 1669390400
transform 1 0 13216 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_463
timestamp 1669390400
transform 1 0 21168 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_464
timestamp 1669390400
transform 1 0 29120 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_465
timestamp 1669390400
transform 1 0 37072 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_466
timestamp 1669390400
transform 1 0 45024 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_467
timestamp 1669390400
transform 1 0 52976 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_468
timestamp 1669390400
transform 1 0 9296 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_469
timestamp 1669390400
transform 1 0 17248 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_470
timestamp 1669390400
transform 1 0 25200 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_471
timestamp 1669390400
transform 1 0 33152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_472
timestamp 1669390400
transform 1 0 41104 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_473
timestamp 1669390400
transform 1 0 49056 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_474
timestamp 1669390400
transform 1 0 57008 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_475
timestamp 1669390400
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_476
timestamp 1669390400
transform 1 0 13216 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_477
timestamp 1669390400
transform 1 0 21168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_478
timestamp 1669390400
transform 1 0 29120 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_479
timestamp 1669390400
transform 1 0 37072 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_480
timestamp 1669390400
transform 1 0 45024 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_481
timestamp 1669390400
transform 1 0 52976 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_482
timestamp 1669390400
transform 1 0 9296 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_483
timestamp 1669390400
transform 1 0 17248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_484
timestamp 1669390400
transform 1 0 25200 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_485
timestamp 1669390400
transform 1 0 33152 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_486
timestamp 1669390400
transform 1 0 41104 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_487
timestamp 1669390400
transform 1 0 49056 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_488
timestamp 1669390400
transform 1 0 57008 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_489
timestamp 1669390400
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_490
timestamp 1669390400
transform 1 0 13216 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_491
timestamp 1669390400
transform 1 0 21168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_492
timestamp 1669390400
transform 1 0 29120 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_493
timestamp 1669390400
transform 1 0 37072 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_494
timestamp 1669390400
transform 1 0 45024 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_495
timestamp 1669390400
transform 1 0 52976 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_496
timestamp 1669390400
transform 1 0 9296 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_497
timestamp 1669390400
transform 1 0 17248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_498
timestamp 1669390400
transform 1 0 25200 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_499
timestamp 1669390400
transform 1 0 33152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_500
timestamp 1669390400
transform 1 0 41104 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_501
timestamp 1669390400
transform 1 0 49056 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_502
timestamp 1669390400
transform 1 0 57008 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_503
timestamp 1669390400
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_504
timestamp 1669390400
transform 1 0 13216 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_505
timestamp 1669390400
transform 1 0 21168 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_506
timestamp 1669390400
transform 1 0 29120 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_507
timestamp 1669390400
transform 1 0 37072 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_508
timestamp 1669390400
transform 1 0 45024 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_509
timestamp 1669390400
transform 1 0 52976 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_510
timestamp 1669390400
transform 1 0 9296 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_511
timestamp 1669390400
transform 1 0 17248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_512
timestamp 1669390400
transform 1 0 25200 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_513
timestamp 1669390400
transform 1 0 33152 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_514
timestamp 1669390400
transform 1 0 41104 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_515
timestamp 1669390400
transform 1 0 49056 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_516
timestamp 1669390400
transform 1 0 57008 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_517
timestamp 1669390400
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_518
timestamp 1669390400
transform 1 0 13216 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_519
timestamp 1669390400
transform 1 0 21168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_520
timestamp 1669390400
transform 1 0 29120 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_521
timestamp 1669390400
transform 1 0 37072 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_522
timestamp 1669390400
transform 1 0 45024 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_523
timestamp 1669390400
transform 1 0 52976 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_524
timestamp 1669390400
transform 1 0 9296 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_525
timestamp 1669390400
transform 1 0 17248 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_526
timestamp 1669390400
transform 1 0 25200 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_527
timestamp 1669390400
transform 1 0 33152 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_528
timestamp 1669390400
transform 1 0 41104 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_529
timestamp 1669390400
transform 1 0 49056 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_530
timestamp 1669390400
transform 1 0 57008 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_531
timestamp 1669390400
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_532
timestamp 1669390400
transform 1 0 13216 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_533
timestamp 1669390400
transform 1 0 21168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_534
timestamp 1669390400
transform 1 0 29120 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_535
timestamp 1669390400
transform 1 0 37072 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_536
timestamp 1669390400
transform 1 0 45024 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_537
timestamp 1669390400
transform 1 0 52976 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_538
timestamp 1669390400
transform 1 0 9296 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_539
timestamp 1669390400
transform 1 0 17248 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_540
timestamp 1669390400
transform 1 0 25200 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_541
timestamp 1669390400
transform 1 0 33152 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_542
timestamp 1669390400
transform 1 0 41104 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_543
timestamp 1669390400
transform 1 0 49056 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_544
timestamp 1669390400
transform 1 0 57008 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_545
timestamp 1669390400
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_546
timestamp 1669390400
transform 1 0 13216 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_547
timestamp 1669390400
transform 1 0 21168 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_548
timestamp 1669390400
transform 1 0 29120 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_549
timestamp 1669390400
transform 1 0 37072 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_550
timestamp 1669390400
transform 1 0 45024 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_551
timestamp 1669390400
transform 1 0 52976 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_552
timestamp 1669390400
transform 1 0 9296 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_553
timestamp 1669390400
transform 1 0 17248 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_554
timestamp 1669390400
transform 1 0 25200 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_555
timestamp 1669390400
transform 1 0 33152 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_556
timestamp 1669390400
transform 1 0 41104 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_557
timestamp 1669390400
transform 1 0 49056 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_558
timestamp 1669390400
transform 1 0 57008 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_559
timestamp 1669390400
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_560
timestamp 1669390400
transform 1 0 13216 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_561
timestamp 1669390400
transform 1 0 21168 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_562
timestamp 1669390400
transform 1 0 29120 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_563
timestamp 1669390400
transform 1 0 37072 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_564
timestamp 1669390400
transform 1 0 45024 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_565
timestamp 1669390400
transform 1 0 52976 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_566
timestamp 1669390400
transform 1 0 9296 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_567
timestamp 1669390400
transform 1 0 17248 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_568
timestamp 1669390400
transform 1 0 25200 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_569
timestamp 1669390400
transform 1 0 33152 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_570
timestamp 1669390400
transform 1 0 41104 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_571
timestamp 1669390400
transform 1 0 49056 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_572
timestamp 1669390400
transform 1 0 57008 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_573
timestamp 1669390400
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_574
timestamp 1669390400
transform 1 0 13216 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_575
timestamp 1669390400
transform 1 0 21168 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_576
timestamp 1669390400
transform 1 0 29120 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_577
timestamp 1669390400
transform 1 0 37072 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_578
timestamp 1669390400
transform 1 0 45024 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_579
timestamp 1669390400
transform 1 0 52976 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_580
timestamp 1669390400
transform 1 0 9296 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_581
timestamp 1669390400
transform 1 0 17248 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_582
timestamp 1669390400
transform 1 0 25200 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_583
timestamp 1669390400
transform 1 0 33152 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_584
timestamp 1669390400
transform 1 0 41104 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_585
timestamp 1669390400
transform 1 0 49056 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_586
timestamp 1669390400
transform 1 0 57008 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_587
timestamp 1669390400
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_588
timestamp 1669390400
transform 1 0 13216 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_589
timestamp 1669390400
transform 1 0 21168 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_590
timestamp 1669390400
transform 1 0 29120 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_591
timestamp 1669390400
transform 1 0 37072 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_592
timestamp 1669390400
transform 1 0 45024 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_593
timestamp 1669390400
transform 1 0 52976 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_594
timestamp 1669390400
transform 1 0 9296 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_595
timestamp 1669390400
transform 1 0 17248 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_596
timestamp 1669390400
transform 1 0 25200 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_597
timestamp 1669390400
transform 1 0 33152 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_598
timestamp 1669390400
transform 1 0 41104 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_599
timestamp 1669390400
transform 1 0 49056 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_600
timestamp 1669390400
transform 1 0 57008 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_601
timestamp 1669390400
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_602
timestamp 1669390400
transform 1 0 13216 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_603
timestamp 1669390400
transform 1 0 21168 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_604
timestamp 1669390400
transform 1 0 29120 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_605
timestamp 1669390400
transform 1 0 37072 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_606
timestamp 1669390400
transform 1 0 45024 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_607
timestamp 1669390400
transform 1 0 52976 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_608
timestamp 1669390400
transform 1 0 9296 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_609
timestamp 1669390400
transform 1 0 17248 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_610
timestamp 1669390400
transform 1 0 25200 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_611
timestamp 1669390400
transform 1 0 33152 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_612
timestamp 1669390400
transform 1 0 41104 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_613
timestamp 1669390400
transform 1 0 49056 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_614
timestamp 1669390400
transform 1 0 57008 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_615
timestamp 1669390400
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_616
timestamp 1669390400
transform 1 0 13216 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_617
timestamp 1669390400
transform 1 0 21168 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_618
timestamp 1669390400
transform 1 0 29120 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_619
timestamp 1669390400
transform 1 0 37072 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_620
timestamp 1669390400
transform 1 0 45024 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_621
timestamp 1669390400
transform 1 0 52976 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_622
timestamp 1669390400
transform 1 0 9296 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_623
timestamp 1669390400
transform 1 0 17248 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_624
timestamp 1669390400
transform 1 0 25200 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_625
timestamp 1669390400
transform 1 0 33152 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_626
timestamp 1669390400
transform 1 0 41104 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_627
timestamp 1669390400
transform 1 0 49056 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_628
timestamp 1669390400
transform 1 0 57008 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_629
timestamp 1669390400
transform 1 0 5264 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_630
timestamp 1669390400
transform 1 0 13216 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_631
timestamp 1669390400
transform 1 0 21168 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_632
timestamp 1669390400
transform 1 0 29120 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_633
timestamp 1669390400
transform 1 0 37072 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_634
timestamp 1669390400
transform 1 0 45024 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_635
timestamp 1669390400
transform 1 0 52976 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_636
timestamp 1669390400
transform 1 0 9296 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_637
timestamp 1669390400
transform 1 0 17248 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_638
timestamp 1669390400
transform 1 0 25200 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_639
timestamp 1669390400
transform 1 0 33152 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_640
timestamp 1669390400
transform 1 0 41104 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_641
timestamp 1669390400
transform 1 0 49056 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_642
timestamp 1669390400
transform 1 0 57008 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_643
timestamp 1669390400
transform 1 0 5264 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_644
timestamp 1669390400
transform 1 0 13216 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_645
timestamp 1669390400
transform 1 0 21168 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_646
timestamp 1669390400
transform 1 0 29120 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_647
timestamp 1669390400
transform 1 0 37072 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_648
timestamp 1669390400
transform 1 0 45024 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_649
timestamp 1669390400
transform 1 0 52976 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_650
timestamp 1669390400
transform 1 0 9296 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_651
timestamp 1669390400
transform 1 0 17248 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_652
timestamp 1669390400
transform 1 0 25200 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_653
timestamp 1669390400
transform 1 0 33152 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_654
timestamp 1669390400
transform 1 0 41104 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_655
timestamp 1669390400
transform 1 0 49056 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_656
timestamp 1669390400
transform 1 0 57008 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_657
timestamp 1669390400
transform 1 0 5264 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_658
timestamp 1669390400
transform 1 0 9184 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_659
timestamp 1669390400
transform 1 0 13104 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_660
timestamp 1669390400
transform 1 0 17024 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_661
timestamp 1669390400
transform 1 0 20944 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_662
timestamp 1669390400
transform 1 0 24864 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_663
timestamp 1669390400
transform 1 0 28784 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_664
timestamp 1669390400
transform 1 0 32704 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_665
timestamp 1669390400
transform 1 0 36624 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_666
timestamp 1669390400
transform 1 0 40544 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_667
timestamp 1669390400
transform 1 0 44464 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_668
timestamp 1669390400
transform 1 0 48384 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_669
timestamp 1669390400
transform 1 0 52304 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_670
timestamp 1669390400
transform 1 0 56224 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1599_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 15344 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1600_
timestamp 1669390400
transform 1 0 8960 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1601_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 6384 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1602_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 17584 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1603_
timestamp 1669390400
transform 1 0 26096 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1604_
timestamp 1669390400
transform 1 0 28448 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _1605_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 14896 0 -1 26656
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1606_
timestamp 1669390400
transform 1 0 13552 0 1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1607_
timestamp 1669390400
transform 1 0 9632 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_4  _1608_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 2240 0 1 26656
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1609_
timestamp 1669390400
transform -1 0 9296 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1610_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 7616 0 1 26656
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1611_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 5152 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1612_
timestamp 1669390400
transform -1 0 9072 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_4  _1613_
timestamp 1669390400
transform 1 0 2240 0 -1 28224
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1614_
timestamp 1669390400
transform 1 0 5936 0 1 23520
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1615_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 9072 0 1 31360
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1616_
timestamp 1669390400
transform 1 0 13328 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1617_
timestamp 1669390400
transform 1 0 6160 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1618_
timestamp 1669390400
transform -1 0 3024 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_4  _1619_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 6720 0 -1 25088
box -86 -86 2438 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1620_
timestamp 1669390400
transform 1 0 7280 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1621_
timestamp 1669390400
transform -1 0 8736 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_4  _1622_
timestamp 1669390400
transform -1 0 9184 0 -1 26656
box -86 -86 2438 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1623_
timestamp 1669390400
transform 1 0 7728 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1624_
timestamp 1669390400
transform 1 0 2912 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _1625_
timestamp 1669390400
transform 1 0 2352 0 1 28224
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1626_
timestamp 1669390400
transform -1 0 4032 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  _1627_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 3248 0 1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1628_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 13216 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1629_
timestamp 1669390400
transform -1 0 15008 0 -1 25088
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1630_
timestamp 1669390400
transform 1 0 12544 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1631_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 12656 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_4  _1632_
timestamp 1669390400
transform 1 0 8400 0 1 23520
box -86 -86 2438 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1633_
timestamp 1669390400
transform -1 0 3696 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1634_
timestamp 1669390400
transform 1 0 5152 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1635_
timestamp 1669390400
transform 1 0 8848 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1636_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 11424 0 1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1637_
timestamp 1669390400
transform -1 0 2576 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_4  _1638_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 11984 0 1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1639_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 11200 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1640_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5600 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1641_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 11984 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1642_
timestamp 1669390400
transform 1 0 3248 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1643_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 15008 0 -1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1644_
timestamp 1669390400
transform 1 0 2240 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1645_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 13552 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1646_
timestamp 1669390400
transform -1 0 17024 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1647_
timestamp 1669390400
transform 1 0 3136 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1648_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 15344 0 -1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1649_
timestamp 1669390400
transform 1 0 15568 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_4  _1650_
timestamp 1669390400
transform 1 0 25536 0 -1 39200
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_4  _1651_
timestamp 1669390400
transform 1 0 13552 0 1 23520
box -86 -86 2438 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1652_
timestamp 1669390400
transform 1 0 12992 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1653_
timestamp 1669390400
transform 1 0 14784 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1654_
timestamp 1669390400
transform 1 0 17808 0 1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_4  _1655_
timestamp 1669390400
transform 1 0 20272 0 -1 50176
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1656_
timestamp 1669390400
transform 1 0 23408 0 -1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_4  _1657_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 21504 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1658_
timestamp 1669390400
transform 1 0 17360 0 1 25088
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1659_
timestamp 1669390400
transform 1 0 20720 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1660_
timestamp 1669390400
transform 1 0 14560 0 1 25088
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1661_
timestamp 1669390400
transform 1 0 11424 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1662_
timestamp 1669390400
transform 1 0 6720 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1663_
timestamp 1669390400
transform 1 0 21504 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1664_
timestamp 1669390400
transform 1 0 19040 0 1 48608
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1665_
timestamp 1669390400
transform 1 0 22512 0 1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1666_
timestamp 1669390400
transform 1 0 23632 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1667_
timestamp 1669390400
transform 1 0 25200 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1668_
timestamp 1669390400
transform 1 0 24192 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1669_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 26208 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1670_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 24976 0 1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1671_
timestamp 1669390400
transform 1 0 24304 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1672_
timestamp 1669390400
transform -1 0 21056 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1673_
timestamp 1669390400
transform 1 0 15120 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1674_
timestamp 1669390400
transform -1 0 3024 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1675_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 12432 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1676_
timestamp 1669390400
transform 1 0 5488 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1677_
timestamp 1669390400
transform -1 0 22400 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1678_
timestamp 1669390400
transform 1 0 9632 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_4  _1679_
timestamp 1669390400
transform 1 0 4032 0 -1 25088
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1680_
timestamp 1669390400
transform -1 0 5264 0 -1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1681_
timestamp 1669390400
transform 1 0 7952 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1682_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 9632 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1683_
timestamp 1669390400
transform 1 0 18368 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1684_
timestamp 1669390400
transform 1 0 21728 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1685_
timestamp 1669390400
transform -1 0 6608 0 -1 26656
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1686_
timestamp 1669390400
transform 1 0 13664 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1687_
timestamp 1669390400
transform 1 0 10528 0 -1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1688_
timestamp 1669390400
transform 1 0 2912 0 -1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1689_
timestamp 1669390400
transform -1 0 19936 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1690_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 10192 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1691_
timestamp 1669390400
transform -1 0 9072 0 -1 29792
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1692_
timestamp 1669390400
transform -1 0 18256 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1693_
timestamp 1669390400
transform 1 0 13776 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1694_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 19824 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1695_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 16016 0 1 29792
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1696_
timestamp 1669390400
transform 1 0 19152 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1697_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 28784 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1698_
timestamp 1669390400
transform -1 0 30464 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_4  _1699_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 30352 0 1 37632
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1700_
timestamp 1669390400
transform 1 0 17472 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1701_
timestamp 1669390400
transform -1 0 17024 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1702_
timestamp 1669390400
transform 1 0 16912 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1703_
timestamp 1669390400
transform -1 0 12208 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1704_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 9632 0 -1 28224
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1705_
timestamp 1669390400
transform -1 0 21616 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1706_
timestamp 1669390400
transform 1 0 21504 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _1707_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 8512 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1708_
timestamp 1669390400
transform 1 0 19936 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1709_
timestamp 1669390400
transform -1 0 11424 0 1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1710_
timestamp 1669390400
transform 1 0 14336 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1711_
timestamp 1669390400
transform -1 0 4144 0 1 29792
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1712_
timestamp 1669390400
transform 1 0 15232 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1713_
timestamp 1669390400
transform 1 0 2800 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1714_
timestamp 1669390400
transform 1 0 1792 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1715_
timestamp 1669390400
transform -1 0 18592 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1716_
timestamp 1669390400
transform -1 0 19712 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1717_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 20272 0 -1 43904
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1718_
timestamp 1669390400
transform 1 0 23408 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or3_2  _1719_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 24080 0 1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _1720_
timestamp 1669390400
transform -1 0 28000 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1721_
timestamp 1669390400
transform -1 0 28672 0 -1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1722_
timestamp 1669390400
transform -1 0 30128 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1723_
timestamp 1669390400
transform -1 0 5712 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _1724_
timestamp 1669390400
transform 1 0 1904 0 -1 29792
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1725_
timestamp 1669390400
transform -1 0 7840 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1726_
timestamp 1669390400
transform -1 0 3248 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1727_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 2912 0 1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1728_
timestamp 1669390400
transform 1 0 3248 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1729_
timestamp 1669390400
transform 1 0 3360 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1730_
timestamp 1669390400
transform 1 0 4032 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1731_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 4144 0 1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1732_
timestamp 1669390400
transform 1 0 3472 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1733_
timestamp 1669390400
transform 1 0 10864 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1734_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 8064 0 1 47040
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1735_
timestamp 1669390400
transform 1 0 4592 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1736_
timestamp 1669390400
transform 1 0 5600 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _1737_
timestamp 1669390400
transform 1 0 3248 0 1 25088
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1738_
timestamp 1669390400
transform 1 0 4592 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1739_
timestamp 1669390400
transform 1 0 4032 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1740_
timestamp 1669390400
transform 1 0 4928 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1741_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 4704 0 -1 48608
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1742_
timestamp 1669390400
transform 1 0 28224 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or3_2  _1743_
timestamp 1669390400
transform 1 0 27664 0 1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _1744_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 29456 0 -1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1745_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 16128 0 1 36064
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1746_
timestamp 1669390400
transform 1 0 13440 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1747_
timestamp 1669390400
transform -1 0 16464 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1748_
timestamp 1669390400
transform -1 0 15008 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1749_
timestamp 1669390400
transform -1 0 15904 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1750_
timestamp 1669390400
transform -1 0 9184 0 -1 28224
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1751_
timestamp 1669390400
transform -1 0 10192 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1752_
timestamp 1669390400
transform 1 0 11648 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1753_
timestamp 1669390400
transform 1 0 11648 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1754_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 7728 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1755_
timestamp 1669390400
transform -1 0 15232 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1756_
timestamp 1669390400
transform 1 0 3136 0 -1 31360
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1757_
timestamp 1669390400
transform 1 0 11536 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _1758_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 12656 0 -1 34496
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1759_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 15568 0 1 37632
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1760_
timestamp 1669390400
transform 1 0 25648 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1761_
timestamp 1669390400
transform -1 0 28224 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1762_
timestamp 1669390400
transform 1 0 26992 0 1 36064
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1763_
timestamp 1669390400
transform -1 0 31024 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1764_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 31136 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1765_
timestamp 1669390400
transform -1 0 30240 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1766_
timestamp 1669390400
transform -1 0 30576 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1767_
timestamp 1669390400
transform -1 0 32144 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1768_
timestamp 1669390400
transform -1 0 30912 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1769_
timestamp 1669390400
transform 1 0 28448 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1770_
timestamp 1669390400
transform -1 0 7616 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1771_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 3584 0 1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1772_
timestamp 1669390400
transform -1 0 7056 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1773_
timestamp 1669390400
transform -1 0 8736 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1774_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 8288 0 1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1775_
timestamp 1669390400
transform -1 0 11088 0 1 50176
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1776_
timestamp 1669390400
transform -1 0 11312 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1777_
timestamp 1669390400
transform 1 0 10528 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1778_
timestamp 1669390400
transform 1 0 17584 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1779_
timestamp 1669390400
transform -1 0 11984 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1780_
timestamp 1669390400
transform 1 0 11984 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1781_
timestamp 1669390400
transform 1 0 9968 0 1 51744
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1782_
timestamp 1669390400
transform -1 0 10976 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _1783_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 11200 0 -1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1784_
timestamp 1669390400
transform -1 0 9184 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1785_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 9632 0 -1 51744
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_4  _1786_
timestamp 1669390400
transform 1 0 26544 0 1 39200
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _1787_
timestamp 1669390400
transform 1 0 10864 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1788_
timestamp 1669390400
transform 1 0 11088 0 1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1789_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 10640 0 -1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1790_
timestamp 1669390400
transform 1 0 11536 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1791_
timestamp 1669390400
transform -1 0 6384 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1792_
timestamp 1669390400
transform -1 0 8288 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1793_
timestamp 1669390400
transform 1 0 7840 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1794_
timestamp 1669390400
transform 1 0 10752 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1795_
timestamp 1669390400
transform 1 0 9632 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1796_
timestamp 1669390400
transform 1 0 10080 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1797_
timestamp 1669390400
transform 1 0 11200 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_4  _1798_
timestamp 1669390400
transform 1 0 17920 0 -1 26656
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1799_
timestamp 1669390400
transform -1 0 6944 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1800_
timestamp 1669390400
transform -1 0 18480 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1801_
timestamp 1669390400
transform 1 0 19376 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1802_
timestamp 1669390400
transform -1 0 9184 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1803_
timestamp 1669390400
transform 1 0 19152 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1804_
timestamp 1669390400
transform 1 0 12432 0 -1 45472
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1805_
timestamp 1669390400
transform 1 0 17584 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1806_
timestamp 1669390400
transform 1 0 19600 0 -1 48608
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1807_
timestamp 1669390400
transform 1 0 18592 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1808_
timestamp 1669390400
transform 1 0 20160 0 -1 29792
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1809_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 19936 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1810_
timestamp 1669390400
transform 1 0 21504 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1811_
timestamp 1669390400
transform -1 0 20720 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1812_
timestamp 1669390400
transform -1 0 21840 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_2  _1813_
timestamp 1669390400
transform 1 0 21504 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1814_
timestamp 1669390400
transform 1 0 21056 0 -1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1815_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 28560 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1816_
timestamp 1669390400
transform -1 0 8176 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1817_
timestamp 1669390400
transform 1 0 6384 0 -1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1818_
timestamp 1669390400
transform 1 0 6048 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1819_
timestamp 1669390400
transform -1 0 5376 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1820_
timestamp 1669390400
transform 1 0 5600 0 1 37632
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1821_
timestamp 1669390400
transform -1 0 8848 0 -1 37632
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1822_
timestamp 1669390400
transform -1 0 17024 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1823_
timestamp 1669390400
transform -1 0 10192 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1824_
timestamp 1669390400
transform -1 0 11312 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1825_
timestamp 1669390400
transform 1 0 17584 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1826_
timestamp 1669390400
transform -1 0 10528 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1827_
timestamp 1669390400
transform 1 0 19040 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1828_
timestamp 1669390400
transform 1 0 19152 0 -1 31360
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__or3_2  _1829_
timestamp 1669390400
transform 1 0 27440 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1830_
timestamp 1669390400
transform 1 0 27664 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1831_
timestamp 1669390400
transform 1 0 30352 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1832_
timestamp 1669390400
transform 1 0 24192 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1833_
timestamp 1669390400
transform 1 0 29456 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _1834_
timestamp 1669390400
transform -1 0 31248 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1835_
timestamp 1669390400
transform 1 0 30688 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1836_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 21280 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1837_
timestamp 1669390400
transform 1 0 21504 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1838_
timestamp 1669390400
transform -1 0 22512 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1839_
timestamp 1669390400
transform -1 0 15680 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1840_
timestamp 1669390400
transform 1 0 15904 0 -1 36064
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1841_
timestamp 1669390400
transform 1 0 18816 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1842_
timestamp 1669390400
transform 1 0 16128 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1843_
timestamp 1669390400
transform 1 0 7616 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1844_
timestamp 1669390400
transform 1 0 2016 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1845_
timestamp 1669390400
transform -1 0 9408 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1846_
timestamp 1669390400
transform 1 0 15008 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1847_
timestamp 1669390400
transform 1 0 17248 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1848_
timestamp 1669390400
transform 1 0 25536 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1849_
timestamp 1669390400
transform 1 0 25872 0 1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_4  _1850_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 27104 0 1 29792
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1851_
timestamp 1669390400
transform -1 0 31920 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1852_
timestamp 1669390400
transform 1 0 10080 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _1853_
timestamp 1669390400
transform 1 0 16576 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1854_
timestamp 1669390400
transform -1 0 18144 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1855_
timestamp 1669390400
transform 1 0 18368 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1856_
timestamp 1669390400
transform 1 0 13552 0 1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1857_
timestamp 1669390400
transform 1 0 14112 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1858_
timestamp 1669390400
transform 1 0 18816 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1859_
timestamp 1669390400
transform 1 0 19488 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1860_
timestamp 1669390400
transform -1 0 22400 0 -1 32928
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1861_
timestamp 1669390400
transform 1 0 23968 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1862_
timestamp 1669390400
transform -1 0 27216 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _1863_
timestamp 1669390400
transform 1 0 28224 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1864_
timestamp 1669390400
transform -1 0 30800 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1865_
timestamp 1669390400
transform -1 0 7280 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _1866_
timestamp 1669390400
transform -1 0 13216 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1867_
timestamp 1669390400
transform -1 0 12992 0 -1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1868_
timestamp 1669390400
transform 1 0 15568 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1869_
timestamp 1669390400
transform 1 0 15680 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1870_
timestamp 1669390400
transform 1 0 10976 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1871_
timestamp 1669390400
transform 1 0 17696 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1872_
timestamp 1669390400
transform 1 0 19712 0 1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1873_
timestamp 1669390400
transform 1 0 19040 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1874_
timestamp 1669390400
transform -1 0 21504 0 -1 37632
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1875_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 21504 0 1 37632
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1876_
timestamp 1669390400
transform 1 0 26096 0 -1 21952
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1877_
timestamp 1669390400
transform 1 0 29568 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1878_
timestamp 1669390400
transform 1 0 30016 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1879_
timestamp 1669390400
transform 1 0 31024 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1880_
timestamp 1669390400
transform 1 0 29792 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _1881_
timestamp 1669390400
transform -1 0 30688 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1882_
timestamp 1669390400
transform -1 0 9184 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _1883_
timestamp 1669390400
transform 1 0 8736 0 1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1884_
timestamp 1669390400
transform 1 0 7504 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _1885_
timestamp 1669390400
transform 1 0 9632 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1886_
timestamp 1669390400
transform -1 0 11088 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1887_
timestamp 1669390400
transform -1 0 3920 0 1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1888_
timestamp 1669390400
transform 1 0 16240 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1889_
timestamp 1669390400
transform 1 0 19712 0 -1 45472
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1890_
timestamp 1669390400
transform 1 0 20384 0 -1 39200
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__or3_2  _1891_
timestamp 1669390400
transform 1 0 26880 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1892_
timestamp 1669390400
transform -1 0 28784 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1893_
timestamp 1669390400
transform -1 0 28336 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1894_
timestamp 1669390400
transform 1 0 28784 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1895_
timestamp 1669390400
transform 1 0 27216 0 -1 36064
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1896_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 25536 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1897_
timestamp 1669390400
transform 1 0 27664 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1898_
timestamp 1669390400
transform 1 0 27776 0 1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1899_
timestamp 1669390400
transform -1 0 27552 0 1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _1900_
timestamp 1669390400
transform 1 0 26768 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1901_
timestamp 1669390400
transform 1 0 26208 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1902_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 27328 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1903_
timestamp 1669390400
transform 1 0 26656 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1904_
timestamp 1669390400
transform -1 0 26432 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1905_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 10528 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1906_
timestamp 1669390400
transform 1 0 16688 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1907_
timestamp 1669390400
transform -1 0 16912 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1908_
timestamp 1669390400
transform 1 0 15344 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1909_
timestamp 1669390400
transform 1 0 15120 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1910_
timestamp 1669390400
transform 1 0 12208 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1911_
timestamp 1669390400
transform 1 0 14672 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1912_
timestamp 1669390400
transform -1 0 16464 0 -1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1913_
timestamp 1669390400
transform 1 0 15456 0 1 51744
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1914_
timestamp 1669390400
transform -1 0 15008 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1915_
timestamp 1669390400
transform -1 0 14896 0 1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1916_
timestamp 1669390400
transform -1 0 14896 0 -1 51744
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1917_
timestamp 1669390400
transform 1 0 22288 0 1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1918_
timestamp 1669390400
transform 1 0 17584 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1919_
timestamp 1669390400
transform 1 0 18256 0 -1 51744
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1920_
timestamp 1669390400
transform -1 0 20608 0 -1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1921_
timestamp 1669390400
transform 1 0 22400 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1922_
timestamp 1669390400
transform 1 0 17920 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1923_
timestamp 1669390400
transform 1 0 17696 0 1 51744
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1924_
timestamp 1669390400
transform 1 0 21840 0 -1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1925_
timestamp 1669390400
transform -1 0 24640 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1926_
timestamp 1669390400
transform 1 0 22848 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1927_
timestamp 1669390400
transform -1 0 15568 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1928_
timestamp 1669390400
transform -1 0 8064 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1929_
timestamp 1669390400
transform 1 0 14224 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1930_
timestamp 1669390400
transform 1 0 3920 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1931_
timestamp 1669390400
transform 1 0 9968 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1932_
timestamp 1669390400
transform -1 0 9632 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1933_
timestamp 1669390400
transform 1 0 5936 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _1934_
timestamp 1669390400
transform 1 0 9856 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1935_
timestamp 1669390400
transform -1 0 15568 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1936_
timestamp 1669390400
transform 1 0 23296 0 1 39200
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1937_
timestamp 1669390400
transform 1 0 11872 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1938_
timestamp 1669390400
transform -1 0 16016 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1939_
timestamp 1669390400
transform 1 0 2016 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _1940_
timestamp 1669390400
transform 1 0 12544 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1941_
timestamp 1669390400
transform 1 0 17584 0 -1 36064
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1942_
timestamp 1669390400
transform -1 0 14000 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1943_
timestamp 1669390400
transform -1 0 18928 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1944_
timestamp 1669390400
transform 1 0 16464 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1945_
timestamp 1669390400
transform 1 0 18144 0 1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1946_
timestamp 1669390400
transform -1 0 20272 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1947_
timestamp 1669390400
transform 1 0 23072 0 -1 40768
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1948_
timestamp 1669390400
transform -1 0 25648 0 1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1949_
timestamp 1669390400
transform 1 0 8400 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1950_
timestamp 1669390400
transform -1 0 13776 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1951_
timestamp 1669390400
transform 1 0 13440 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1952_
timestamp 1669390400
transform 1 0 13888 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1953_
timestamp 1669390400
transform 1 0 14000 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1954_
timestamp 1669390400
transform 1 0 21504 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1955_
timestamp 1669390400
transform 1 0 13552 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1956_
timestamp 1669390400
transform 1 0 18256 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1957_
timestamp 1669390400
transform 1 0 21504 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1958_
timestamp 1669390400
transform 1 0 23408 0 1 42336
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1959_
timestamp 1669390400
transform 1 0 3808 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1960_
timestamp 1669390400
transform -1 0 2800 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1961_
timestamp 1669390400
transform -1 0 3584 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _1962_
timestamp 1669390400
transform 1 0 3248 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1963_
timestamp 1669390400
transform 1 0 5264 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1964_
timestamp 1669390400
transform 1 0 4256 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1965_
timestamp 1669390400
transform 1 0 2576 0 1 36064
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1966_
timestamp 1669390400
transform -1 0 4032 0 -1 37632
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1967_
timestamp 1669390400
transform 1 0 2912 0 -1 36064
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1968_
timestamp 1669390400
transform 1 0 23968 0 1 34496
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1969_
timestamp 1669390400
transform 1 0 2352 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1970_
timestamp 1669390400
transform 1 0 3024 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1971_
timestamp 1669390400
transform 1 0 5936 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1972_
timestamp 1669390400
transform 1 0 5936 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1973_
timestamp 1669390400
transform 1 0 7168 0 -1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1974_
timestamp 1669390400
transform 1 0 8400 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1975_
timestamp 1669390400
transform 1 0 6048 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1976_
timestamp 1669390400
transform 1 0 23856 0 1 37632
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1977_
timestamp 1669390400
transform -1 0 3024 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1978_
timestamp 1669390400
transform -1 0 3696 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1979_
timestamp 1669390400
transform 1 0 3248 0 1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1980_
timestamp 1669390400
transform -1 0 10528 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1981_
timestamp 1669390400
transform -1 0 10752 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1982_
timestamp 1669390400
transform -1 0 10864 0 -1 43904
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1983_
timestamp 1669390400
transform 1 0 10528 0 1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1984_
timestamp 1669390400
transform 1 0 9072 0 1 47040
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1985_
timestamp 1669390400
transform -1 0 9184 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1986_
timestamp 1669390400
transform 1 0 23072 0 -1 36064
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1987_
timestamp 1669390400
transform 1 0 6608 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1988_
timestamp 1669390400
transform 1 0 10752 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1989_
timestamp 1669390400
transform -1 0 9968 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1990_
timestamp 1669390400
transform 1 0 10192 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1991_
timestamp 1669390400
transform -1 0 11872 0 -1 29792
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1992_
timestamp 1669390400
transform 1 0 11760 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1993_
timestamp 1669390400
transform 1 0 15008 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1994_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 15008 0 1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1995_
timestamp 1669390400
transform 1 0 16240 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1996_
timestamp 1669390400
transform 1 0 22400 0 1 29792
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1997_
timestamp 1669390400
transform 1 0 7504 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1998_
timestamp 1669390400
transform 1 0 8624 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1999_
timestamp 1669390400
transform -1 0 7504 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2000_
timestamp 1669390400
transform -1 0 7280 0 1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2001_
timestamp 1669390400
transform 1 0 6160 0 1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2002_
timestamp 1669390400
transform 1 0 6496 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2003_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5600 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2004_
timestamp 1669390400
transform 1 0 7504 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2005_
timestamp 1669390400
transform -1 0 7728 0 -1 45472
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2006_
timestamp 1669390400
transform -1 0 8176 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2007_
timestamp 1669390400
transform 1 0 22960 0 -1 50176
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2008_
timestamp 1669390400
transform 1 0 17584 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2009_
timestamp 1669390400
transform 1 0 17808 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2010_
timestamp 1669390400
transform 1 0 12208 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2011_
timestamp 1669390400
transform 1 0 13664 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2012_
timestamp 1669390400
transform 1 0 14000 0 1 28224
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2013_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 16464 0 1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2014_
timestamp 1669390400
transform -1 0 14560 0 -1 26656
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2015_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 20272 0 1 26656
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _2016_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 18480 0 1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2017_
timestamp 1669390400
transform -1 0 20496 0 -1 28224
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2018_
timestamp 1669390400
transform -1 0 37856 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2019_
timestamp 1669390400
transform -1 0 18144 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2020_
timestamp 1669390400
transform -1 0 17136 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2021_
timestamp 1669390400
transform 1 0 15456 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2022_
timestamp 1669390400
transform 1 0 15680 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2023_
timestamp 1669390400
transform 1 0 22624 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2024_
timestamp 1669390400
transform -1 0 22064 0 -1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2025_
timestamp 1669390400
transform 1 0 19936 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2026_
timestamp 1669390400
transform 1 0 21056 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2027_
timestamp 1669390400
transform 1 0 22624 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2028_
timestamp 1669390400
transform 1 0 23296 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2029_
timestamp 1669390400
transform 1 0 39536 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2030_
timestamp 1669390400
transform 1 0 40992 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2031_
timestamp 1669390400
transform 1 0 14224 0 1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2032_
timestamp 1669390400
transform 1 0 13776 0 -1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2033_
timestamp 1669390400
transform 1 0 14560 0 1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2034_
timestamp 1669390400
transform 1 0 16240 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _2035_
timestamp 1669390400
transform 1 0 16912 0 1 47040
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2036_
timestamp 1669390400
transform 1 0 17584 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _2037_
timestamp 1669390400
transform -1 0 21056 0 1 45472
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _2038_
timestamp 1669390400
transform 1 0 17696 0 -1 47040
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2039_
timestamp 1669390400
transform 1 0 23744 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2040_
timestamp 1669390400
transform -1 0 31584 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2041_
timestamp 1669390400
transform 1 0 4256 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2042_
timestamp 1669390400
transform 1 0 4928 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2043_
timestamp 1669390400
transform -1 0 8064 0 -1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2044_
timestamp 1669390400
transform 1 0 6272 0 -1 42336
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2045_
timestamp 1669390400
transform -1 0 12320 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2046_
timestamp 1669390400
transform -1 0 6048 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2047_
timestamp 1669390400
transform 1 0 5600 0 1 40768
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2048_
timestamp 1669390400
transform 1 0 22848 0 -1 29792
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2049_
timestamp 1669390400
transform 1 0 30016 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2050_
timestamp 1669390400
transform -1 0 32816 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2051_
timestamp 1669390400
transform 1 0 30240 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2052_
timestamp 1669390400
transform -1 0 30576 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2053_
timestamp 1669390400
transform -1 0 29008 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2054_
timestamp 1669390400
transform 1 0 26768 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2055_
timestamp 1669390400
transform 1 0 26880 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2056_
timestamp 1669390400
transform -1 0 27440 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2057_
timestamp 1669390400
transform 1 0 25536 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2058_
timestamp 1669390400
transform -1 0 26208 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2059_
timestamp 1669390400
transform -1 0 26544 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2060_
timestamp 1669390400
transform 1 0 24864 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2061_
timestamp 1669390400
transform -1 0 26992 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2062_
timestamp 1669390400
transform -1 0 24192 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2063_
timestamp 1669390400
transform 1 0 24864 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2064_
timestamp 1669390400
transform 1 0 24192 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2065_
timestamp 1669390400
transform -1 0 25312 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2066_
timestamp 1669390400
transform -1 0 24528 0 1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _2067_
timestamp 1669390400
transform 1 0 19600 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2068_
timestamp 1669390400
transform 1 0 20272 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _2069_
timestamp 1669390400
transform -1 0 20720 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  _2070_
timestamp 1669390400
transform 1 0 19376 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _2071_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 24192 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _2072_
timestamp 1669390400
transform 1 0 41440 0 -1 40768
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _2073_
timestamp 1669390400
transform -1 0 48944 0 1 39200
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2074_
timestamp 1669390400
transform -1 0 25088 0 -1 21952
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2075_
timestamp 1669390400
transform 1 0 21504 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2076_
timestamp 1669390400
transform 1 0 19936 0 -1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2077_
timestamp 1669390400
transform 1 0 21168 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2078_
timestamp 1669390400
transform 1 0 25872 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2079_
timestamp 1669390400
transform 1 0 45472 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2080_
timestamp 1669390400
transform 1 0 49728 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2081_
timestamp 1669390400
transform 1 0 45360 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2082_
timestamp 1669390400
transform 1 0 23408 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2083_
timestamp 1669390400
transform 1 0 23856 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _2084_
timestamp 1669390400
transform 1 0 40320 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2085_
timestamp 1669390400
transform 1 0 46032 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2086_
timestamp 1669390400
transform 1 0 47936 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2087_
timestamp 1669390400
transform 1 0 49616 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2088_
timestamp 1669390400
transform 1 0 51856 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2089_
timestamp 1669390400
transform 1 0 51968 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2090_
timestamp 1669390400
transform -1 0 54208 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2091_
timestamp 1669390400
transform 1 0 26096 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2092_
timestamp 1669390400
transform 1 0 16464 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _2093_
timestamp 1669390400
transform 1 0 21168 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  _2094_
timestamp 1669390400
transform 1 0 27216 0 1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2095_
timestamp 1669390400
transform 1 0 34048 0 -1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2096_
timestamp 1669390400
transform -1 0 21056 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2097_
timestamp 1669390400
transform 1 0 25536 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2098_
timestamp 1669390400
transform 1 0 38080 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2099_
timestamp 1669390400
transform -1 0 21056 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2100_
timestamp 1669390400
transform 1 0 19152 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2101_
timestamp 1669390400
transform -1 0 22400 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2102_
timestamp 1669390400
transform 1 0 23408 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _2103_
timestamp 1669390400
transform 1 0 38192 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2104_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 38416 0 1 31360
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2105_
timestamp 1669390400
transform 1 0 41776 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2106_
timestamp 1669390400
transform 1 0 29456 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2107_
timestamp 1669390400
transform 1 0 32480 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2108_
timestamp 1669390400
transform -1 0 27440 0 1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2109_
timestamp 1669390400
transform 1 0 26432 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _2110_
timestamp 1669390400
transform 1 0 24080 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2111_
timestamp 1669390400
transform 1 0 28560 0 -1 32928
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2112_
timestamp 1669390400
transform -1 0 36736 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2113_
timestamp 1669390400
transform 1 0 34272 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2114_
timestamp 1669390400
transform 1 0 35392 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2115_
timestamp 1669390400
transform 1 0 39872 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2116_
timestamp 1669390400
transform 1 0 25536 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2117_
timestamp 1669390400
transform 1 0 32144 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2118_
timestamp 1669390400
transform -1 0 36736 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2119_
timestamp 1669390400
transform 1 0 39648 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2120_
timestamp 1669390400
transform 1 0 41440 0 -1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2121_
timestamp 1669390400
transform 1 0 42672 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2122_
timestamp 1669390400
transform -1 0 44016 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  _2123_
timestamp 1669390400
transform 1 0 46368 0 -1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _2124_
timestamp 1669390400
transform 1 0 45808 0 1 40768
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2125_
timestamp 1669390400
transform 1 0 45248 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2126_
timestamp 1669390400
transform -1 0 47712 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2127_
timestamp 1669390400
transform 1 0 23968 0 1 32928
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2128_
timestamp 1669390400
transform 1 0 27216 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2129_
timestamp 1669390400
transform 1 0 39536 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2130_
timestamp 1669390400
transform 1 0 47936 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2131_
timestamp 1669390400
transform 1 0 49504 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2132_
timestamp 1669390400
transform 1 0 50400 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2133_
timestamp 1669390400
transform 1 0 51408 0 1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2134_
timestamp 1669390400
transform 1 0 52304 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2135_
timestamp 1669390400
transform -1 0 54208 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2136_
timestamp 1669390400
transform 1 0 29792 0 1 40768
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2137_
timestamp 1669390400
transform 1 0 36512 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2138_
timestamp 1669390400
transform -1 0 23968 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_4  _2139_
timestamp 1669390400
transform 1 0 23856 0 1 25088
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2140_
timestamp 1669390400
transform 1 0 20272 0 -1 25088
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__and2_4  _2141_
timestamp 1669390400
transform 1 0 21280 0 -1 26656
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2142_
timestamp 1669390400
transform 1 0 28000 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2143_
timestamp 1669390400
transform 1 0 23072 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2144_
timestamp 1669390400
transform -1 0 23856 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_4  _2145_
timestamp 1669390400
transform 1 0 26096 0 -1 25088
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2146_
timestamp 1669390400
transform 1 0 29456 0 1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _2147_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 30688 0 1 28224
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2148_
timestamp 1669390400
transform 1 0 37408 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _2149_
timestamp 1669390400
transform 1 0 30240 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2150_
timestamp 1669390400
transform 1 0 30240 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2151_
timestamp 1669390400
transform -1 0 33712 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2152_
timestamp 1669390400
transform -1 0 31360 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2153_
timestamp 1669390400
transform -1 0 32032 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _2154_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 35168 0 1 29792
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2155_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 30128 0 1 32928
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2156_
timestamp 1669390400
transform 1 0 43456 0 1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2157_
timestamp 1669390400
transform 1 0 42448 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2158_
timestamp 1669390400
transform 1 0 44688 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2159_
timestamp 1669390400
transform -1 0 46256 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2160_
timestamp 1669390400
transform 1 0 30688 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2161_
timestamp 1669390400
transform 1 0 29568 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2162_
timestamp 1669390400
transform -1 0 32816 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2163_
timestamp 1669390400
transform 1 0 33488 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2164_
timestamp 1669390400
transform 1 0 27888 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2165_
timestamp 1669390400
transform 1 0 29456 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _2166_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 33488 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2167_
timestamp 1669390400
transform 1 0 33936 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2168_
timestamp 1669390400
transform 1 0 34160 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _2169_
timestamp 1669390400
transform 1 0 30240 0 -1 29792
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2170_
timestamp 1669390400
transform 1 0 45360 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2171_
timestamp 1669390400
transform 1 0 45696 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2172_
timestamp 1669390400
transform 1 0 40768 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2173_
timestamp 1669390400
transform -1 0 32256 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2174_
timestamp 1669390400
transform 1 0 32032 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2175_
timestamp 1669390400
transform 1 0 40320 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2176_
timestamp 1669390400
transform 1 0 30912 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2177_
timestamp 1669390400
transform -1 0 32256 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2178_
timestamp 1669390400
transform -1 0 42784 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2179_
timestamp 1669390400
transform 1 0 42112 0 -1 34496
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2180_
timestamp 1669390400
transform 1 0 47376 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2181_
timestamp 1669390400
transform 1 0 54880 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2182_
timestamp 1669390400
transform 1 0 53312 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2183_
timestamp 1669390400
transform 1 0 55104 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2184_
timestamp 1669390400
transform -1 0 56672 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2185_
timestamp 1669390400
transform 1 0 46256 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2186_
timestamp 1669390400
transform -1 0 47824 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2187_
timestamp 1669390400
transform 1 0 45248 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2188_
timestamp 1669390400
transform 1 0 40992 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2189_
timestamp 1669390400
transform 1 0 33488 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2190_
timestamp 1669390400
transform -1 0 36400 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2191_
timestamp 1669390400
transform 1 0 34496 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2192_
timestamp 1669390400
transform 1 0 39424 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2193_
timestamp 1669390400
transform 1 0 27552 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2194_
timestamp 1669390400
transform -1 0 30352 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2195_
timestamp 1669390400
transform 1 0 39424 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2196_
timestamp 1669390400
transform 1 0 42224 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2197_
timestamp 1669390400
transform 1 0 43904 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2198_
timestamp 1669390400
transform -1 0 32592 0 -1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2199_
timestamp 1669390400
transform 1 0 33152 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2200_
timestamp 1669390400
transform 1 0 32144 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2201_
timestamp 1669390400
transform -1 0 34384 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2202_
timestamp 1669390400
transform 1 0 35056 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2203_
timestamp 1669390400
transform 1 0 24528 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  _2204_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 27104 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2205_
timestamp 1669390400
transform 1 0 31584 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _2206_
timestamp 1669390400
transform -1 0 36960 0 1 31360
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2207_
timestamp 1669390400
transform 1 0 35728 0 -1 37632
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2208_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 45808 0 -1 37632
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2209_
timestamp 1669390400
transform 1 0 52752 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2210_
timestamp 1669390400
transform 1 0 49392 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2211_
timestamp 1669390400
transform -1 0 51184 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2212_
timestamp 1669390400
transform 1 0 41552 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2213_
timestamp 1669390400
transform -1 0 44128 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2214_
timestamp 1669390400
transform 1 0 42448 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2215_
timestamp 1669390400
transform -1 0 55104 0 1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _2216_
timestamp 1669390400
transform 1 0 46704 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2217_
timestamp 1669390400
transform 1 0 42448 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2218_
timestamp 1669390400
transform 1 0 48048 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _2219_
timestamp 1669390400
transform -1 0 47936 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2220_
timestamp 1669390400
transform -1 0 48384 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2221_
timestamp 1669390400
transform 1 0 48160 0 1 34496
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2222_
timestamp 1669390400
transform 1 0 50400 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2223_
timestamp 1669390400
transform 1 0 51296 0 1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2224_
timestamp 1669390400
transform 1 0 53312 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2225_
timestamp 1669390400
transform 1 0 54320 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2226_
timestamp 1669390400
transform 1 0 56224 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2227_
timestamp 1669390400
transform 1 0 56224 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2228_
timestamp 1669390400
transform 1 0 57344 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2229_
timestamp 1669390400
transform 1 0 51856 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2230_
timestamp 1669390400
transform -1 0 54208 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2231_
timestamp 1669390400
transform 1 0 53312 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2232_
timestamp 1669390400
transform -1 0 55328 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2233_
timestamp 1669390400
transform -1 0 50736 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2234_
timestamp 1669390400
transform -1 0 50064 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2235_
timestamp 1669390400
transform -1 0 50960 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2236_
timestamp 1669390400
transform 1 0 43680 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2237_
timestamp 1669390400
transform 1 0 42560 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2238_
timestamp 1669390400
transform -1 0 44464 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2239_
timestamp 1669390400
transform 1 0 49952 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2240_
timestamp 1669390400
transform 1 0 19712 0 1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _2241_
timestamp 1669390400
transform 1 0 39648 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2242_
timestamp 1669390400
transform 1 0 39984 0 -1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2243_
timestamp 1669390400
transform 1 0 46256 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2244_
timestamp 1669390400
transform 1 0 48048 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2245_
timestamp 1669390400
transform 1 0 49392 0 -1 42336
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2246_
timestamp 1669390400
transform -1 0 51296 0 1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2247_
timestamp 1669390400
transform 1 0 49392 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2248_
timestamp 1669390400
transform 1 0 46144 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2249_
timestamp 1669390400
transform -1 0 47600 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2250_
timestamp 1669390400
transform 1 0 46480 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2251_
timestamp 1669390400
transform 1 0 39536 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2252_
timestamp 1669390400
transform -1 0 32256 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2253_
timestamp 1669390400
transform -1 0 34272 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2254_
timestamp 1669390400
transform 1 0 33936 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2255_
timestamp 1669390400
transform 1 0 21728 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2256_
timestamp 1669390400
transform -1 0 27664 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2257_
timestamp 1669390400
transform 1 0 42224 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2258_
timestamp 1669390400
transform 1 0 36736 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2259_
timestamp 1669390400
transform -1 0 38304 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2260_
timestamp 1669390400
transform 1 0 37856 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2261_
timestamp 1669390400
transform 1 0 39648 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2262_
timestamp 1669390400
transform 1 0 32368 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2263_
timestamp 1669390400
transform 1 0 34160 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2264_
timestamp 1669390400
transform 1 0 35728 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2265_
timestamp 1669390400
transform -1 0 36400 0 -1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2266_
timestamp 1669390400
transform 1 0 33712 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2267_
timestamp 1669390400
transform -1 0 34832 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2268_
timestamp 1669390400
transform 1 0 35392 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_4  _2269_
timestamp 1669390400
transform 1 0 22624 0 -1 25088
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _2270_
timestamp 1669390400
transform -1 0 23296 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_4  _2271_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 29792 0 1 39200
box -86 -86 5798 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2272_
timestamp 1669390400
transform 1 0 37408 0 1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2273_
timestamp 1669390400
transform -1 0 45024 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2274_
timestamp 1669390400
transform 1 0 43568 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2275_
timestamp 1669390400
transform 1 0 47600 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2276_
timestamp 1669390400
transform 1 0 50960 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2277_
timestamp 1669390400
transform 1 0 53088 0 -1 39200
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2278_
timestamp 1669390400
transform 1 0 56224 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2279_
timestamp 1669390400
transform -1 0 52080 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2280_
timestamp 1669390400
transform 1 0 50624 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2281_
timestamp 1669390400
transform 1 0 48048 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2282_
timestamp 1669390400
transform 1 0 49840 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2283_
timestamp 1669390400
transform 1 0 50512 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2284_
timestamp 1669390400
transform 1 0 47600 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2285_
timestamp 1669390400
transform 1 0 48720 0 1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2286_
timestamp 1669390400
transform 1 0 38192 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2287_
timestamp 1669390400
transform 1 0 38528 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2288_
timestamp 1669390400
transform -1 0 40432 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2289_
timestamp 1669390400
transform -1 0 48048 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _2290_
timestamp 1669390400
transform 1 0 25760 0 -1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2291_
timestamp 1669390400
transform -1 0 46256 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2292_
timestamp 1669390400
transform 1 0 44016 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2293_
timestamp 1669390400
transform 1 0 45360 0 1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2294_
timestamp 1669390400
transform 1 0 46368 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2295_
timestamp 1669390400
transform 1 0 47488 0 -1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2296_
timestamp 1669390400
transform 1 0 48496 0 1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2297_
timestamp 1669390400
transform 1 0 43456 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2298_
timestamp 1669390400
transform 1 0 44240 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2299_
timestamp 1669390400
transform 1 0 44464 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2300_
timestamp 1669390400
transform 1 0 36960 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2301_
timestamp 1669390400
transform -1 0 39200 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2302_
timestamp 1669390400
transform 1 0 37968 0 -1 34496
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2303_
timestamp 1669390400
transform 1 0 41888 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2304_
timestamp 1669390400
transform 1 0 37632 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2305_
timestamp 1669390400
transform -1 0 31920 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2306_
timestamp 1669390400
transform -1 0 35728 0 -1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2307_
timestamp 1669390400
transform 1 0 35504 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_4  _2308_
timestamp 1669390400
transform 1 0 31248 0 1 42336
box -86 -86 5798 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2309_
timestamp 1669390400
transform 1 0 37520 0 1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2310_
timestamp 1669390400
transform 1 0 39536 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2311_
timestamp 1669390400
transform 1 0 39536 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2312_
timestamp 1669390400
transform 1 0 41104 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2313_
timestamp 1669390400
transform 1 0 42336 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2314_
timestamp 1669390400
transform 1 0 47936 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2315_
timestamp 1669390400
transform 1 0 49392 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2316_
timestamp 1669390400
transform 1 0 50848 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2317_
timestamp 1669390400
transform 1 0 51632 0 -1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2318_
timestamp 1669390400
transform -1 0 54880 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2319_
timestamp 1669390400
transform 1 0 53424 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2320_
timestamp 1669390400
transform -1 0 54208 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2321_
timestamp 1669390400
transform 1 0 53312 0 1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2322_
timestamp 1669390400
transform -1 0 58688 0 -1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2323_
timestamp 1669390400
transform 1 0 57344 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2324_
timestamp 1669390400
transform 1 0 45472 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _2325_
timestamp 1669390400
transform -1 0 40320 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2326_
timestamp 1669390400
transform -1 0 44016 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2327_
timestamp 1669390400
transform 1 0 48160 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2328_
timestamp 1669390400
transform 1 0 49392 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2329_
timestamp 1669390400
transform 1 0 49392 0 -1 28224
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2330_
timestamp 1669390400
transform 1 0 50288 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2331_
timestamp 1669390400
transform 1 0 29792 0 -1 28224
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2332_
timestamp 1669390400
transform -1 0 33488 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2333_
timestamp 1669390400
transform 1 0 33488 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2334_
timestamp 1669390400
transform -1 0 34496 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2335_
timestamp 1669390400
transform 1 0 38752 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2336_
timestamp 1669390400
transform -1 0 39424 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2337_
timestamp 1669390400
transform 1 0 39648 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2338_
timestamp 1669390400
transform 1 0 38416 0 1 29792
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2339_
timestamp 1669390400
transform -1 0 35616 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2340_
timestamp 1669390400
transform 1 0 39312 0 1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2341_
timestamp 1669390400
transform 1 0 39648 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2342_
timestamp 1669390400
transform 1 0 53424 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2343_
timestamp 1669390400
transform 1 0 54992 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2344_
timestamp 1669390400
transform 1 0 55328 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2345_
timestamp 1669390400
transform -1 0 58240 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2346_
timestamp 1669390400
transform 1 0 31920 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2347_
timestamp 1669390400
transform 1 0 26880 0 -1 28224
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _2348_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 35280 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _2349_
timestamp 1669390400
transform -1 0 35728 0 1 26656
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2350_
timestamp 1669390400
transform -1 0 36176 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2351_
timestamp 1669390400
transform 1 0 33712 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2352_
timestamp 1669390400
transform 1 0 34384 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2353_
timestamp 1669390400
transform -1 0 36400 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2354_
timestamp 1669390400
transform 1 0 37184 0 -1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2355_
timestamp 1669390400
transform 1 0 41440 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2356_
timestamp 1669390400
transform 1 0 41440 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2357_
timestamp 1669390400
transform 1 0 43008 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2358_
timestamp 1669390400
transform -1 0 44240 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2359_
timestamp 1669390400
transform 1 0 45248 0 -1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2360_
timestamp 1669390400
transform 1 0 56896 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2361_
timestamp 1669390400
transform 1 0 54656 0 1 28224
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2362_
timestamp 1669390400
transform 1 0 57344 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2363_
timestamp 1669390400
transform 1 0 57568 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2364_
timestamp 1669390400
transform 1 0 55776 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2365_
timestamp 1669390400
transform 1 0 57008 0 1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2366_
timestamp 1669390400
transform -1 0 58016 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2367_
timestamp 1669390400
transform -1 0 58240 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2368_
timestamp 1669390400
transform 1 0 56672 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2369_
timestamp 1669390400
transform 1 0 57120 0 1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2370_
timestamp 1669390400
transform -1 0 58016 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2371_
timestamp 1669390400
transform -1 0 58240 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2372_
timestamp 1669390400
transform -1 0 58688 0 -1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2373_
timestamp 1669390400
transform 1 0 55216 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _2374_
timestamp 1669390400
transform 1 0 41440 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2375_
timestamp 1669390400
transform 1 0 25312 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2376_
timestamp 1669390400
transform 1 0 22848 0 1 28224
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _2377_
timestamp 1669390400
transform -1 0 40880 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2378_
timestamp 1669390400
transform -1 0 35392 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2379_
timestamp 1669390400
transform 1 0 34384 0 -1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2380_
timestamp 1669390400
transform -1 0 41104 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2381_
timestamp 1669390400
transform 1 0 38864 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2382_
timestamp 1669390400
transform 1 0 40320 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2383_
timestamp 1669390400
transform -1 0 42784 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2384_
timestamp 1669390400
transform 1 0 52192 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2385_
timestamp 1669390400
transform -1 0 45808 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2386_
timestamp 1669390400
transform 1 0 45808 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _2387_
timestamp 1669390400
transform 1 0 46592 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2388_
timestamp 1669390400
transform 1 0 48608 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2389_
timestamp 1669390400
transform -1 0 48944 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2390_
timestamp 1669390400
transform -1 0 50400 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2391_
timestamp 1669390400
transform -1 0 51072 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2392_
timestamp 1669390400
transform 1 0 52528 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2393_
timestamp 1669390400
transform 1 0 54208 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2394_
timestamp 1669390400
transform 1 0 53312 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2395_
timestamp 1669390400
transform 1 0 36624 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2396_
timestamp 1669390400
transform 1 0 27328 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2397_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 29456 0 1 23520
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2398_
timestamp 1669390400
transform 1 0 35504 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2399_
timestamp 1669390400
transform 1 0 34384 0 1 23520
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2400_
timestamp 1669390400
transform 1 0 35168 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2401_
timestamp 1669390400
transform 1 0 37408 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2402_
timestamp 1669390400
transform 1 0 37072 0 -1 25088
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2403_
timestamp 1669390400
transform 1 0 41440 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2404_
timestamp 1669390400
transform 1 0 43680 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2405_
timestamp 1669390400
transform 1 0 42000 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2406_
timestamp 1669390400
transform 1 0 40768 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2407_
timestamp 1669390400
transform -1 0 43232 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2408_
timestamp 1669390400
transform 1 0 42448 0 -1 28224
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2409_
timestamp 1669390400
transform 1 0 45360 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2410_
timestamp 1669390400
transform -1 0 54656 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2411_
timestamp 1669390400
transform 1 0 45360 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2412_
timestamp 1669390400
transform -1 0 53536 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2413_
timestamp 1669390400
transform -1 0 58464 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2414_
timestamp 1669390400
transform -1 0 58240 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2415_
timestamp 1669390400
transform -1 0 58240 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2416_
timestamp 1669390400
transform -1 0 56896 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2417_
timestamp 1669390400
transform -1 0 58688 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2418_
timestamp 1669390400
transform -1 0 58464 0 1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2419_
timestamp 1669390400
transform -1 0 58016 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2420_
timestamp 1669390400
transform 1 0 57008 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2421_
timestamp 1669390400
transform -1 0 58688 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2422_
timestamp 1669390400
transform -1 0 56784 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2423_
timestamp 1669390400
transform -1 0 58688 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2424_
timestamp 1669390400
transform 1 0 39984 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2425_
timestamp 1669390400
transform 1 0 38752 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2426_
timestamp 1669390400
transform 1 0 43008 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2427_
timestamp 1669390400
transform 1 0 44352 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2428_
timestamp 1669390400
transform 1 0 35728 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2429_
timestamp 1669390400
transform 1 0 42784 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2430_
timestamp 1669390400
transform 1 0 44576 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2431_
timestamp 1669390400
transform -1 0 47936 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2432_
timestamp 1669390400
transform 1 0 44352 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2433_
timestamp 1669390400
transform -1 0 46368 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2434_
timestamp 1669390400
transform 1 0 48272 0 1 23520
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2435_
timestamp 1669390400
transform 1 0 50848 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2436_
timestamp 1669390400
transform 1 0 50064 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2437_
timestamp 1669390400
transform -1 0 37968 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2438_
timestamp 1669390400
transform 1 0 35616 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2439_
timestamp 1669390400
transform 1 0 35952 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _2440_
timestamp 1669390400
transform 1 0 33488 0 -1 20384
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _2441_
timestamp 1669390400
transform -1 0 30128 0 -1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _2442_
timestamp 1669390400
transform 1 0 32368 0 1 20384
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2443_
timestamp 1669390400
transform 1 0 35392 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _2444_
timestamp 1669390400
transform 1 0 35728 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2445_
timestamp 1669390400
transform -1 0 38304 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2446_
timestamp 1669390400
transform 1 0 37632 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2447_
timestamp 1669390400
transform 1 0 46592 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2448_
timestamp 1669390400
transform 1 0 45472 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2449_
timestamp 1669390400
transform 1 0 48160 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2450_
timestamp 1669390400
transform 1 0 47040 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2451_
timestamp 1669390400
transform 1 0 43008 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2452_
timestamp 1669390400
transform 1 0 49392 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2453_
timestamp 1669390400
transform 1 0 50960 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2454_
timestamp 1669390400
transform -1 0 52528 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2455_
timestamp 1669390400
transform 1 0 52304 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2456_
timestamp 1669390400
transform 1 0 53984 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2457_
timestamp 1669390400
transform 1 0 53424 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2458_
timestamp 1669390400
transform 1 0 53648 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2459_
timestamp 1669390400
transform -1 0 58688 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2460_
timestamp 1669390400
transform -1 0 56224 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2461_
timestamp 1669390400
transform -1 0 55888 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2462_
timestamp 1669390400
transform -1 0 56896 0 1 37632
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2463_
timestamp 1669390400
transform 1 0 55888 0 -1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2464_
timestamp 1669390400
transform -1 0 56336 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2465_
timestamp 1669390400
transform -1 0 55888 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2466_
timestamp 1669390400
transform 1 0 42000 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2467_
timestamp 1669390400
transform 1 0 43680 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2468_
timestamp 1669390400
transform 1 0 40096 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2469_
timestamp 1669390400
transform 1 0 42560 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2470_
timestamp 1669390400
transform 1 0 42560 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2471_
timestamp 1669390400
transform 1 0 31584 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2472_
timestamp 1669390400
transform 1 0 32368 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2473_
timestamp 1669390400
transform 1 0 41328 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2474_
timestamp 1669390400
transform -1 0 42784 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2475_
timestamp 1669390400
transform 1 0 41776 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2476_
timestamp 1669390400
transform 1 0 42224 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2477_
timestamp 1669390400
transform 1 0 43904 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2478_
timestamp 1669390400
transform 1 0 43344 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2479_
timestamp 1669390400
transform 1 0 46704 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2480_
timestamp 1669390400
transform 1 0 48720 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2481_
timestamp 1669390400
transform 1 0 47600 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2482_
timestamp 1669390400
transform 1 0 49840 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2483_
timestamp 1669390400
transform 1 0 31472 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2484_
timestamp 1669390400
transform 1 0 32368 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2485_
timestamp 1669390400
transform 1 0 33376 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2486_
timestamp 1669390400
transform 1 0 34944 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2487_
timestamp 1669390400
transform -1 0 34944 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2488_
timestamp 1669390400
transform 1 0 35504 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2489_
timestamp 1669390400
transform 1 0 35504 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2490_
timestamp 1669390400
transform 1 0 37184 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2491_
timestamp 1669390400
transform 1 0 37520 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2492_
timestamp 1669390400
transform -1 0 39312 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2493_
timestamp 1669390400
transform 1 0 36288 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2494_
timestamp 1669390400
transform 1 0 36960 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2495_
timestamp 1669390400
transform 1 0 37072 0 -1 20384
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2496_
timestamp 1669390400
transform 1 0 45248 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2497_
timestamp 1669390400
transform 1 0 43344 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2498_
timestamp 1669390400
transform 1 0 45696 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2499_
timestamp 1669390400
transform -1 0 47712 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2500_
timestamp 1669390400
transform 1 0 46144 0 1 20384
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2501_
timestamp 1669390400
transform 1 0 49392 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2502_
timestamp 1669390400
transform 1 0 48944 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2503_
timestamp 1669390400
transform -1 0 50736 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2504_
timestamp 1669390400
transform 1 0 50176 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2505_
timestamp 1669390400
transform 1 0 50736 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2506_
timestamp 1669390400
transform 1 0 51184 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2507_
timestamp 1669390400
transform 1 0 51296 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2508_
timestamp 1669390400
transform 1 0 53312 0 1 21952
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2509_
timestamp 1669390400
transform -1 0 56896 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2510_
timestamp 1669390400
transform -1 0 55776 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2511_
timestamp 1669390400
transform 1 0 55552 0 1 23520
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2512_
timestamp 1669390400
transform 1 0 54656 0 1 18816
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2513_
timestamp 1669390400
transform -1 0 58464 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2514_
timestamp 1669390400
transform 1 0 54208 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2515_
timestamp 1669390400
transform 1 0 57344 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2516_
timestamp 1669390400
transform 1 0 39984 0 -1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2517_
timestamp 1669390400
transform 1 0 38864 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2518_
timestamp 1669390400
transform 1 0 39648 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2519_
timestamp 1669390400
transform 1 0 42224 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2520_
timestamp 1669390400
transform -1 0 43904 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2521_
timestamp 1669390400
transform 1 0 42672 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2522_
timestamp 1669390400
transform 1 0 43344 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2523_
timestamp 1669390400
transform 1 0 45584 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2524_
timestamp 1669390400
transform 1 0 46480 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2525_
timestamp 1669390400
transform 1 0 43344 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2526_
timestamp 1669390400
transform 1 0 43568 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2527_
timestamp 1669390400
transform 1 0 46816 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2528_
timestamp 1669390400
transform 1 0 49392 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2529_
timestamp 1669390400
transform 1 0 48272 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2530_
timestamp 1669390400
transform 1 0 49168 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2531_
timestamp 1669390400
transform 1 0 32480 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2532_
timestamp 1669390400
transform 1 0 35168 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2533_
timestamp 1669390400
transform -1 0 36176 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2534_
timestamp 1669390400
transform -1 0 31136 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2535_
timestamp 1669390400
transform -1 0 33712 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2536_
timestamp 1669390400
transform 1 0 33488 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2537_
timestamp 1669390400
transform -1 0 37632 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2538_
timestamp 1669390400
transform -1 0 40992 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2539_
timestamp 1669390400
transform 1 0 35616 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2540_
timestamp 1669390400
transform -1 0 38528 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2541_
timestamp 1669390400
transform 1 0 38416 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2542_
timestamp 1669390400
transform -1 0 47936 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2543_
timestamp 1669390400
transform 1 0 46256 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2544_
timestamp 1669390400
transform 1 0 46480 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2545_
timestamp 1669390400
transform -1 0 47936 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2546_
timestamp 1669390400
transform 1 0 46144 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2547_
timestamp 1669390400
transform 1 0 49056 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2548_
timestamp 1669390400
transform 1 0 49392 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2549_
timestamp 1669390400
transform -1 0 51520 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2550_
timestamp 1669390400
transform 1 0 49616 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2551_
timestamp 1669390400
transform 1 0 51520 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2552_
timestamp 1669390400
transform 1 0 51968 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2553_
timestamp 1669390400
transform -1 0 53872 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2554_
timestamp 1669390400
transform 1 0 51744 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2555_
timestamp 1669390400
transform 1 0 53312 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2556_
timestamp 1669390400
transform 1 0 52304 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2557_
timestamp 1669390400
transform -1 0 54208 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2558_
timestamp 1669390400
transform 1 0 52640 0 -1 20384
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2559_
timestamp 1669390400
transform 1 0 55888 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2560_
timestamp 1669390400
transform 1 0 53536 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2561_
timestamp 1669390400
transform -1 0 58688 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2562_
timestamp 1669390400
transform 1 0 42672 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2563_
timestamp 1669390400
transform -1 0 44464 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2564_
timestamp 1669390400
transform 1 0 45360 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2565_
timestamp 1669390400
transform 1 0 45472 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2566_
timestamp 1669390400
transform 1 0 46480 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2567_
timestamp 1669390400
transform 1 0 49392 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2568_
timestamp 1669390400
transform 1 0 48720 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2569_
timestamp 1669390400
transform 1 0 46144 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2570_
timestamp 1669390400
transform 1 0 46144 0 -1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2571_
timestamp 1669390400
transform -1 0 31472 0 1 17248
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2572_
timestamp 1669390400
transform 1 0 32368 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2573_
timestamp 1669390400
transform 1 0 33936 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2574_
timestamp 1669390400
transform 1 0 42560 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2575_
timestamp 1669390400
transform 1 0 43568 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2576_
timestamp 1669390400
transform 1 0 44128 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2577_
timestamp 1669390400
transform -1 0 45248 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2578_
timestamp 1669390400
transform 1 0 37856 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2579_
timestamp 1669390400
transform 1 0 37408 0 1 14112
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2580_
timestamp 1669390400
transform 1 0 45808 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2581_
timestamp 1669390400
transform 1 0 46144 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2582_
timestamp 1669390400
transform -1 0 47936 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2583_
timestamp 1669390400
transform 1 0 46032 0 1 12544
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2584_
timestamp 1669390400
transform 1 0 48608 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2585_
timestamp 1669390400
transform 1 0 49392 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2586_
timestamp 1669390400
transform 1 0 49840 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2587_
timestamp 1669390400
transform 1 0 50400 0 1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2588_
timestamp 1669390400
transform 1 0 52864 0 -1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_2  _2589_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 51744 0 -1 14112
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2590_
timestamp 1669390400
transform 1 0 53536 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2591_
timestamp 1669390400
transform 1 0 53760 0 1 10976
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2592_
timestamp 1669390400
transform 1 0 51408 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2593_
timestamp 1669390400
transform 1 0 33936 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2594_
timestamp 1669390400
transform -1 0 34720 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2595_
timestamp 1669390400
transform 1 0 33488 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2596_
timestamp 1669390400
transform 1 0 32032 0 -1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2597_
timestamp 1669390400
transform -1 0 35728 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2598_
timestamp 1669390400
transform 1 0 39760 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2599_
timestamp 1669390400
transform 1 0 41776 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2600_
timestamp 1669390400
transform 1 0 42560 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2601_
timestamp 1669390400
transform -1 0 43680 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2602_
timestamp 1669390400
transform -1 0 35168 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2603_
timestamp 1669390400
transform 1 0 34384 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2604_
timestamp 1669390400
transform 1 0 34720 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2605_
timestamp 1669390400
transform 1 0 43568 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2606_
timestamp 1669390400
transform 1 0 45024 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2607_
timestamp 1669390400
transform -1 0 43344 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2608_
timestamp 1669390400
transform 1 0 43568 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2609_
timestamp 1669390400
transform 1 0 45472 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2610_
timestamp 1669390400
transform 1 0 46592 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2611_
timestamp 1669390400
transform -1 0 48272 0 -1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2612_
timestamp 1669390400
transform 1 0 50288 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2613_
timestamp 1669390400
transform -1 0 51856 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2614_
timestamp 1669390400
transform 1 0 50400 0 -1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2615_
timestamp 1669390400
transform 1 0 50288 0 1 7840
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _2616_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 53312 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2617_
timestamp 1669390400
transform 1 0 52528 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2618_
timestamp 1669390400
transform 1 0 54432 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2619_
timestamp 1669390400
transform -1 0 55776 0 1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2620_
timestamp 1669390400
transform -1 0 57904 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2621_
timestamp 1669390400
transform 1 0 56224 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2622_
timestamp 1669390400
transform 1 0 56336 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2623_
timestamp 1669390400
transform 1 0 33936 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2624_
timestamp 1669390400
transform -1 0 35168 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2625_
timestamp 1669390400
transform 1 0 33376 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2626_
timestamp 1669390400
transform -1 0 36400 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2627_
timestamp 1669390400
transform 1 0 33152 0 1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2628_
timestamp 1669390400
transform 1 0 35056 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2629_
timestamp 1669390400
transform 1 0 39984 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2630_
timestamp 1669390400
transform 1 0 38752 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2631_
timestamp 1669390400
transform -1 0 39312 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2632_
timestamp 1669390400
transform 1 0 34496 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2633_
timestamp 1669390400
transform 1 0 36288 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2634_
timestamp 1669390400
transform 1 0 36288 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2635_
timestamp 1669390400
transform 1 0 36960 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2636_
timestamp 1669390400
transform 1 0 39872 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2637_
timestamp 1669390400
transform 1 0 36848 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2638_
timestamp 1669390400
transform 1 0 38640 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2639_
timestamp 1669390400
transform 1 0 40880 0 1 3136
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2640_
timestamp 1669390400
transform 1 0 41664 0 1 3136
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2641_
timestamp 1669390400
transform -1 0 45248 0 -1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2642_
timestamp 1669390400
transform 1 0 41440 0 -1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2643_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 39760 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2644_
timestamp 1669390400
transform 1 0 33936 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2645_
timestamp 1669390400
transform 1 0 34720 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2646_
timestamp 1669390400
transform 1 0 37408 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2647_
timestamp 1669390400
transform 1 0 34720 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2648_
timestamp 1669390400
transform 1 0 34832 0 -1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2649_
timestamp 1669390400
transform 1 0 37184 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2650_
timestamp 1669390400
transform 1 0 41104 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2651_
timestamp 1669390400
transform 1 0 41440 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2652_
timestamp 1669390400
transform -1 0 40992 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2653_
timestamp 1669390400
transform 1 0 37408 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2654_
timestamp 1669390400
transform -1 0 40320 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2655_
timestamp 1669390400
transform 1 0 37408 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2656_
timestamp 1669390400
transform -1 0 40096 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2657_
timestamp 1669390400
transform 1 0 39088 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2658_
timestamp 1669390400
transform 1 0 40432 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2659_
timestamp 1669390400
transform 1 0 41552 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2660_
timestamp 1669390400
transform 1 0 40432 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2661_
timestamp 1669390400
transform 1 0 36512 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2662_
timestamp 1669390400
transform 1 0 37408 0 1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2663_
timestamp 1669390400
transform 1 0 37408 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2664_
timestamp 1669390400
transform 1 0 36736 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2665_
timestamp 1669390400
transform 1 0 38752 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2666_
timestamp 1669390400
transform -1 0 39312 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2667_
timestamp 1669390400
transform 1 0 38976 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2668_
timestamp 1669390400
transform -1 0 41216 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2669_
timestamp 1669390400
transform 1 0 40880 0 1 4704
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2670_
timestamp 1669390400
transform 1 0 41440 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2671_
timestamp 1669390400
transform -1 0 43232 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2672_
timestamp 1669390400
transform -1 0 44800 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2673_
timestamp 1669390400
transform 1 0 46032 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2674_
timestamp 1669390400
transform 1 0 47040 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2675_
timestamp 1669390400
transform 1 0 45360 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2676_
timestamp 1669390400
transform 1 0 48608 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2677_
timestamp 1669390400
transform 1 0 54208 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2678_
timestamp 1669390400
transform 1 0 52976 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2679_
timestamp 1669390400
transform -1 0 54992 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2680_
timestamp 1669390400
transform 1 0 55552 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2681_
timestamp 1669390400
transform 1 0 57344 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_2  _2682_
timestamp 1669390400
transform 1 0 55552 0 1 21952
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2683_
timestamp 1669390400
transform -1 0 58688 0 1 20384
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2684_
timestamp 1669390400
transform 1 0 57344 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2685_
timestamp 1669390400
transform -1 0 58464 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2686_
timestamp 1669390400
transform -1 0 57456 0 1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2687_
timestamp 1669390400
transform -1 0 56784 0 -1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2688_
timestamp 1669390400
transform -1 0 56560 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2689_
timestamp 1669390400
transform -1 0 58688 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2690_
timestamp 1669390400
transform -1 0 58240 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2691_
timestamp 1669390400
transform 1 0 57344 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2692_
timestamp 1669390400
transform 1 0 57904 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2693_
timestamp 1669390400
transform 1 0 56784 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2694_
timestamp 1669390400
transform 1 0 43568 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2695_
timestamp 1669390400
transform 1 0 44016 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2696_
timestamp 1669390400
transform -1 0 45472 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2697_
timestamp 1669390400
transform 1 0 45360 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2698_
timestamp 1669390400
transform 1 0 46480 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2699_
timestamp 1669390400
transform 1 0 43568 0 1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2700_
timestamp 1669390400
transform 1 0 45360 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2701_
timestamp 1669390400
transform 1 0 46480 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2702_
timestamp 1669390400
transform 1 0 45360 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2703_
timestamp 1669390400
transform -1 0 43120 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2704_
timestamp 1669390400
transform -1 0 35280 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _2705_
timestamp 1669390400
transform 1 0 38752 0 -1 40768
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2706_
timestamp 1669390400
transform 1 0 40880 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2707_
timestamp 1669390400
transform -1 0 42448 0 1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2708_
timestamp 1669390400
transform 1 0 37968 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2709_
timestamp 1669390400
transform 1 0 27664 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2710_
timestamp 1669390400
transform 1 0 35840 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_4  _2711_
timestamp 1669390400
transform 1 0 31248 0 1 43904
box -86 -86 5798 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2712_
timestamp 1669390400
transform 1 0 37408 0 1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2713_
timestamp 1669390400
transform 1 0 38864 0 -1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2714_
timestamp 1669390400
transform 1 0 41328 0 1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2715_
timestamp 1669390400
transform 1 0 43120 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2716_
timestamp 1669390400
transform 1 0 45472 0 -1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2717_
timestamp 1669390400
transform 1 0 42672 0 -1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2718_
timestamp 1669390400
transform -1 0 46256 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2719_
timestamp 1669390400
transform -1 0 44912 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2720_
timestamp 1669390400
transform 1 0 42672 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2721_
timestamp 1669390400
transform -1 0 43792 0 1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2722_
timestamp 1669390400
transform 1 0 39200 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2723_
timestamp 1669390400
transform -1 0 41104 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2724_
timestamp 1669390400
transform -1 0 40992 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2725_
timestamp 1669390400
transform 1 0 42000 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2726_
timestamp 1669390400
transform 1 0 42896 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2727_
timestamp 1669390400
transform 1 0 38192 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2728_
timestamp 1669390400
transform 1 0 38640 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2729_
timestamp 1669390400
transform -1 0 40544 0 -1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2730_
timestamp 1669390400
transform 1 0 37632 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2731_
timestamp 1669390400
transform -1 0 35952 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2732_
timestamp 1669390400
transform -1 0 36176 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2733_
timestamp 1669390400
transform 1 0 34944 0 -1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _2734_
timestamp 1669390400
transform 1 0 33488 0 -1 31360
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2735_
timestamp 1669390400
transform 1 0 35168 0 -1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2736_
timestamp 1669390400
transform 1 0 37632 0 -1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2737_
timestamp 1669390400
transform 1 0 39200 0 -1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2738_
timestamp 1669390400
transform 1 0 41440 0 -1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2739_
timestamp 1669390400
transform 1 0 42784 0 -1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2740_
timestamp 1669390400
transform 1 0 45472 0 -1 51744
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2741_
timestamp 1669390400
transform 1 0 48048 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2742_
timestamp 1669390400
transform 1 0 49392 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2743_
timestamp 1669390400
transform -1 0 49840 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2744_
timestamp 1669390400
transform -1 0 48944 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2745_
timestamp 1669390400
transform 1 0 49504 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2746_
timestamp 1669390400
transform 1 0 46032 0 1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2747_
timestamp 1669390400
transform 1 0 49392 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2748_
timestamp 1669390400
transform 1 0 48048 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2749_
timestamp 1669390400
transform -1 0 49840 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2750_
timestamp 1669390400
transform 1 0 48944 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2751_
timestamp 1669390400
transform 1 0 44800 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2752_
timestamp 1669390400
transform -1 0 46480 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2753_
timestamp 1669390400
transform -1 0 47264 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2754_
timestamp 1669390400
transform 1 0 45808 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2755_
timestamp 1669390400
transform -1 0 44016 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2756_
timestamp 1669390400
transform 1 0 41664 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2757_
timestamp 1669390400
transform -1 0 42112 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2758_
timestamp 1669390400
transform 1 0 41888 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2759_
timestamp 1669390400
transform 1 0 40208 0 1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2760_
timestamp 1669390400
transform 1 0 39312 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2761_
timestamp 1669390400
transform -1 0 39760 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2762_
timestamp 1669390400
transform 1 0 38304 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2763_
timestamp 1669390400
transform -1 0 37184 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2764_
timestamp 1669390400
transform -1 0 40768 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2765_
timestamp 1669390400
transform -1 0 40096 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2766_
timestamp 1669390400
transform 1 0 35616 0 1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2767_
timestamp 1669390400
transform -1 0 36736 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2768_
timestamp 1669390400
transform 1 0 32256 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2769_
timestamp 1669390400
transform -1 0 33712 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2770_
timestamp 1669390400
transform -1 0 34832 0 -1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_4  _2771_
timestamp 1669390400
transform -1 0 35840 0 1 47040
box -86 -86 5798 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2772_
timestamp 1669390400
transform 1 0 33488 0 -1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2773_
timestamp 1669390400
transform 1 0 35392 0 1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2774_
timestamp 1669390400
transform 1 0 37408 0 1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2775_
timestamp 1669390400
transform 1 0 38304 0 -1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2776_
timestamp 1669390400
transform 1 0 39424 0 1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2777_
timestamp 1669390400
transform 1 0 42336 0 1 53312
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2778_
timestamp 1669390400
transform 1 0 45696 0 1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2779_
timestamp 1669390400
transform 1 0 49392 0 -1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2780_
timestamp 1669390400
transform 1 0 45920 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2781_
timestamp 1669390400
transform -1 0 37856 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2782_
timestamp 1669390400
transform 1 0 35392 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2783_
timestamp 1669390400
transform -1 0 36960 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2784_
timestamp 1669390400
transform -1 0 34384 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2785_
timestamp 1669390400
transform 1 0 33936 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2786_
timestamp 1669390400
transform 1 0 31472 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2787_
timestamp 1669390400
transform -1 0 29904 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2788_
timestamp 1669390400
transform 1 0 30128 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2789_
timestamp 1669390400
transform 1 0 29456 0 1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_4  _2790_
timestamp 1669390400
transform -1 0 35168 0 1 48608
box -86 -86 5798 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2791_
timestamp 1669390400
transform 1 0 29904 0 -1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2792_
timestamp 1669390400
transform 1 0 31584 0 -1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2793_
timestamp 1669390400
transform 1 0 32704 0 1 51744
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2794_
timestamp 1669390400
transform 1 0 35840 0 -1 53312
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2795_
timestamp 1669390400
transform 1 0 38976 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2796_
timestamp 1669390400
transform 1 0 39200 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2797_
timestamp 1669390400
transform 1 0 39200 0 1 53312
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2798_
timestamp 1669390400
transform 1 0 41552 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2799_
timestamp 1669390400
transform -1 0 43344 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2800_
timestamp 1669390400
transform 1 0 42560 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2801_
timestamp 1669390400
transform 1 0 42112 0 1 54880
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2802_
timestamp 1669390400
transform 1 0 45920 0 1 56448
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2803_
timestamp 1669390400
transform -1 0 51744 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2804_
timestamp 1669390400
transform 1 0 51072 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2805_
timestamp 1669390400
transform -1 0 53648 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2806_
timestamp 1669390400
transform 1 0 51184 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2807_
timestamp 1669390400
transform 1 0 53312 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2808_
timestamp 1669390400
transform 1 0 48272 0 1 50176
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2809_
timestamp 1669390400
transform 1 0 51184 0 -1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2810_
timestamp 1669390400
transform -1 0 54656 0 1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2811_
timestamp 1669390400
transform -1 0 51968 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2812_
timestamp 1669390400
transform 1 0 49392 0 -1 53312
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2813_
timestamp 1669390400
transform 1 0 51072 0 1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2814_
timestamp 1669390400
transform -1 0 52752 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2815_
timestamp 1669390400
transform -1 0 52864 0 1 56448
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2816_
timestamp 1669390400
transform 1 0 52304 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2817_
timestamp 1669390400
transform -1 0 51856 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2818_
timestamp 1669390400
transform -1 0 50848 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2819_
timestamp 1669390400
transform -1 0 48608 0 1 53312
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2820_
timestamp 1669390400
transform -1 0 47040 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2821_
timestamp 1669390400
transform -1 0 46816 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2822_
timestamp 1669390400
transform 1 0 33488 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2823_
timestamp 1669390400
transform -1 0 33936 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2824_
timestamp 1669390400
transform 1 0 32928 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2825_
timestamp 1669390400
transform -1 0 34832 0 -1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2826_
timestamp 1669390400
transform -1 0 33712 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2827_
timestamp 1669390400
transform -1 0 29680 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2828_
timestamp 1669390400
transform -1 0 29008 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2829_
timestamp 1669390400
transform -1 0 27216 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2830_
timestamp 1669390400
transform 1 0 27888 0 -1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2831_
timestamp 1669390400
transform -1 0 31584 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_4  _2832_
timestamp 1669390400
transform -1 0 32704 0 -1 48608
box -86 -86 5798 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2833_
timestamp 1669390400
transform -1 0 28448 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2834_
timestamp 1669390400
transform 1 0 26992 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2835_
timestamp 1669390400
transform 1 0 26208 0 1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2836_
timestamp 1669390400
transform 1 0 27104 0 -1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2837_
timestamp 1669390400
transform 1 0 29456 0 1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2838_
timestamp 1669390400
transform 1 0 29680 0 -1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2839_
timestamp 1669390400
transform 1 0 31696 0 -1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2840_
timestamp 1669390400
transform 1 0 33152 0 1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2841_
timestamp 1669390400
transform 1 0 34944 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2842_
timestamp 1669390400
transform 1 0 36064 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2843_
timestamp 1669390400
transform 1 0 35728 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2844_
timestamp 1669390400
transform 1 0 35168 0 1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2845_
timestamp 1669390400
transform -1 0 39872 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2846_
timestamp 1669390400
transform -1 0 42112 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2847_
timestamp 1669390400
transform -1 0 39984 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2848_
timestamp 1669390400
transform 1 0 40208 0 1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2849_
timestamp 1669390400
transform 1 0 27104 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2850_
timestamp 1669390400
transform -1 0 30128 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2851_
timestamp 1669390400
transform 1 0 29680 0 -1 53312
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2852_
timestamp 1669390400
transform 1 0 29456 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2853_
timestamp 1669390400
transform 1 0 20272 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2854_
timestamp 1669390400
transform 1 0 18928 0 1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2855_
timestamp 1669390400
transform 1 0 20272 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_4  _2856_
timestamp 1669390400
transform -1 0 32368 0 -1 47040
box -86 -86 5798 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2857_
timestamp 1669390400
transform -1 0 20272 0 -1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2858_
timestamp 1669390400
transform -1 0 27440 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2859_
timestamp 1669390400
transform -1 0 27664 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2860_
timestamp 1669390400
transform 1 0 19488 0 1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2861_
timestamp 1669390400
transform 1 0 25312 0 1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2862_
timestamp 1669390400
transform 1 0 26880 0 1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2863_
timestamp 1669390400
transform 1 0 32368 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2864_
timestamp 1669390400
transform 1 0 32032 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2865_
timestamp 1669390400
transform -1 0 30800 0 1 56448
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2866_
timestamp 1669390400
transform -1 0 35840 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2867_
timestamp 1669390400
transform -1 0 38304 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2868_
timestamp 1669390400
transform -1 0 36736 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2869_
timestamp 1669390400
transform 1 0 35616 0 1 58016
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2870_
timestamp 1669390400
transform 1 0 41440 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2871_
timestamp 1669390400
transform -1 0 45696 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2872_
timestamp 1669390400
transform 1 0 44128 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2873_
timestamp 1669390400
transform 1 0 38528 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2874_
timestamp 1669390400
transform -1 0 39648 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2875_
timestamp 1669390400
transform 1 0 36176 0 -1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2876_
timestamp 1669390400
transform 1 0 37408 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2877_
timestamp 1669390400
transform -1 0 34944 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2878_
timestamp 1669390400
transform -1 0 29008 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2879_
timestamp 1669390400
transform -1 0 27664 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2880_
timestamp 1669390400
transform 1 0 26208 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2881_
timestamp 1669390400
transform -1 0 14336 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2882_
timestamp 1669390400
transform -1 0 13440 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _2883_
timestamp 1669390400
transform -1 0 24416 0 1 48608
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2884_
timestamp 1669390400
transform 1 0 11760 0 1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2885_
timestamp 1669390400
transform 1 0 13552 0 1 58016
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2886_
timestamp 1669390400
transform -1 0 20384 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2887_
timestamp 1669390400
transform -1 0 19712 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2888_
timestamp 1669390400
transform -1 0 19264 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2889_
timestamp 1669390400
transform 1 0 18816 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2890_
timestamp 1669390400
transform 1 0 18704 0 1 58016
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2891_
timestamp 1669390400
transform 1 0 25200 0 1 58016
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2892_
timestamp 1669390400
transform 1 0 27664 0 -1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2893_
timestamp 1669390400
transform 1 0 29680 0 -1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2894_
timestamp 1669390400
transform -1 0 29008 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2895_
timestamp 1669390400
transform -1 0 31024 0 -1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2896_
timestamp 1669390400
transform 1 0 29120 0 -1 58016
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2897_
timestamp 1669390400
transform 1 0 29792 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2898_
timestamp 1669390400
transform 1 0 32368 0 -1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2899_
timestamp 1669390400
transform -1 0 35280 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2900_
timestamp 1669390400
transform 1 0 53760 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2901_
timestamp 1669390400
transform -1 0 54432 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2902_
timestamp 1669390400
transform 1 0 54096 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2903_
timestamp 1669390400
transform 1 0 55440 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_2  _2904_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 53200 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _2905_
timestamp 1669390400
transform 1 0 54768 0 -1 17248
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2906_
timestamp 1669390400
transform -1 0 56784 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2907_
timestamp 1669390400
transform -1 0 56672 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2908_
timestamp 1669390400
transform -1 0 56896 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2909_
timestamp 1669390400
transform 1 0 55552 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2910_
timestamp 1669390400
transform 1 0 47936 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2911_
timestamp 1669390400
transform 1 0 55216 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2912_
timestamp 1669390400
transform -1 0 57456 0 1 7840
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _2913_
timestamp 1669390400
transform -1 0 58688 0 1 15680
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _2914_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 55104 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2915_
timestamp 1669390400
transform 1 0 55328 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2916_
timestamp 1669390400
transform 1 0 56000 0 1 48608
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2917_
timestamp 1669390400
transform 1 0 51632 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2918_
timestamp 1669390400
transform 1 0 53312 0 1 56448
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2919_
timestamp 1669390400
transform 1 0 47040 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2920_
timestamp 1669390400
transform -1 0 42784 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2921_
timestamp 1669390400
transform 1 0 32816 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2922_
timestamp 1669390400
transform 1 0 34832 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2923_
timestamp 1669390400
transform 1 0 43008 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2924_
timestamp 1669390400
transform 1 0 37968 0 -1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2925_
timestamp 1669390400
transform 1 0 38528 0 1 58016
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2926_
timestamp 1669390400
transform 1 0 35504 0 1 56448
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2927_
timestamp 1669390400
transform 1 0 43568 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2928_
timestamp 1669390400
transform 1 0 44016 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2929_
timestamp 1669390400
transform 1 0 43120 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2930_
timestamp 1669390400
transform -1 0 38864 0 -1 58016
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2931_
timestamp 1669390400
transform 1 0 28448 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2932_
timestamp 1669390400
transform -1 0 54208 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2933_
timestamp 1669390400
transform -1 0 54544 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2934_
timestamp 1669390400
transform -1 0 53872 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2935_
timestamp 1669390400
transform -1 0 54656 0 1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2936_
timestamp 1669390400
transform 1 0 51744 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2937_
timestamp 1669390400
transform -1 0 50736 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2938_
timestamp 1669390400
transform -1 0 50736 0 -1 56448
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2939_
timestamp 1669390400
transform 1 0 47936 0 -1 54880
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2940_
timestamp 1669390400
transform -1 0 56224 0 -1 47040
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2941_
timestamp 1669390400
transform 1 0 56112 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2942_
timestamp 1669390400
transform -1 0 56000 0 -1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2943_
timestamp 1669390400
transform -1 0 53984 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2944_
timestamp 1669390400
transform -1 0 55104 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _2945_
timestamp 1669390400
transform -1 0 54880 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2946_
timestamp 1669390400
transform -1 0 56448 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2947_
timestamp 1669390400
transform 1 0 54768 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2948_
timestamp 1669390400
transform -1 0 55440 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2949_
timestamp 1669390400
transform 1 0 52304 0 -1 42336
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2950_
timestamp 1669390400
transform -1 0 54208 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2951_
timestamp 1669390400
transform -1 0 55888 0 1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2952_
timestamp 1669390400
transform 1 0 50512 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2953_
timestamp 1669390400
transform 1 0 51520 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2954_
timestamp 1669390400
transform 1 0 51632 0 -1 48608
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2955_
timestamp 1669390400
transform -1 0 54320 0 -1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2956_
timestamp 1669390400
transform 1 0 51744 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2957_
timestamp 1669390400
transform -1 0 53872 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2958_
timestamp 1669390400
transform -1 0 52864 0 1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2959_
timestamp 1669390400
transform -1 0 51408 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2960_
timestamp 1669390400
transform 1 0 49840 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2961_
timestamp 1669390400
transform -1 0 48720 0 1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2962_
timestamp 1669390400
transform -1 0 48160 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2963_
timestamp 1669390400
transform 1 0 46368 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2964_
timestamp 1669390400
transform -1 0 47712 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2965_
timestamp 1669390400
transform 1 0 46928 0 1 54880
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2966_
timestamp 1669390400
transform 1 0 36064 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2967_
timestamp 1669390400
transform -1 0 44800 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2968_
timestamp 1669390400
transform -1 0 40768 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2969_
timestamp 1669390400
transform 1 0 40208 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2970_
timestamp 1669390400
transform 1 0 39872 0 1 58016
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2971_
timestamp 1669390400
transform -1 0 43680 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2972_
timestamp 1669390400
transform 1 0 39872 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2973_
timestamp 1669390400
transform -1 0 45024 0 -1 56448
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2974_
timestamp 1669390400
transform 1 0 38976 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2975_
timestamp 1669390400
transform 1 0 18592 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2976_
timestamp 1669390400
transform 1 0 12544 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2977_
timestamp 1669390400
transform -1 0 15680 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2978_
timestamp 1669390400
transform -1 0 14336 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2979_
timestamp 1669390400
transform 1 0 10864 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2980_
timestamp 1669390400
transform -1 0 14224 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2981_
timestamp 1669390400
transform -1 0 24192 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2982_
timestamp 1669390400
transform -1 0 13104 0 1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2983_
timestamp 1669390400
transform 1 0 11648 0 -1 56448
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2984_
timestamp 1669390400
transform 1 0 13216 0 -1 58016
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2985_
timestamp 1669390400
transform -1 0 15232 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2986_
timestamp 1669390400
transform 1 0 14224 0 -1 59584
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2987_
timestamp 1669390400
transform 1 0 15568 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2988_
timestamp 1669390400
transform 1 0 18368 0 -1 59584
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2989_
timestamp 1669390400
transform 1 0 24304 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2990_
timestamp 1669390400
transform -1 0 27664 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2991_
timestamp 1669390400
transform 1 0 26096 0 -1 59584
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2992_
timestamp 1669390400
transform 1 0 28448 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2993_
timestamp 1669390400
transform 1 0 30128 0 -1 58016
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2994_
timestamp 1669390400
transform -1 0 35168 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2995_
timestamp 1669390400
transform 1 0 30912 0 1 58016
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2996_
timestamp 1669390400
transform 1 0 33824 0 -1 59584
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2997_
timestamp 1669390400
transform -1 0 32816 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2998_
timestamp 1669390400
transform 1 0 31024 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2999_
timestamp 1669390400
transform -1 0 39648 0 1 56448
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3000_
timestamp 1669390400
transform 1 0 26768 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _3001_
timestamp 1669390400
transform -1 0 28784 0 -1 59584
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3002_
timestamp 1669390400
transform 1 0 33488 0 -1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3003_
timestamp 1669390400
transform 1 0 33488 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _3004_
timestamp 1669390400
transform -1 0 43680 0 1 58016
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3005_
timestamp 1669390400
transform 1 0 12320 0 1 56448
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _3006_
timestamp 1669390400
transform 1 0 13328 0 -1 56448
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3007_
timestamp 1669390400
transform 1 0 14448 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3008_
timestamp 1669390400
transform -1 0 23408 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3009_
timestamp 1669390400
transform -1 0 17136 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _3010_
timestamp 1669390400
transform 1 0 14560 0 -1 54880
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3011_
timestamp 1669390400
transform 1 0 15568 0 1 56448
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3012_
timestamp 1669390400
transform -1 0 16800 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3013_
timestamp 1669390400
transform 1 0 19712 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3014_
timestamp 1669390400
transform 1 0 19936 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3015_
timestamp 1669390400
transform 1 0 17024 0 1 58016
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _3016_
timestamp 1669390400
transform 1 0 22624 0 1 59584
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3017_
timestamp 1669390400
transform -1 0 16800 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _3018_
timestamp 1669390400
transform 1 0 15680 0 1 53312
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _3019_
timestamp 1669390400
transform 1 0 17136 0 1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _3020_
timestamp 1669390400
transform 1 0 21840 0 1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3021_
timestamp 1669390400
transform -1 0 25088 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3022_
timestamp 1669390400
transform -1 0 25424 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _3023_
timestamp 1669390400
transform 1 0 23072 0 -1 59584
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3024_
timestamp 1669390400
transform 1 0 21728 0 1 58016
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3025_
timestamp 1669390400
transform 1 0 23296 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3026_
timestamp 1669390400
transform 1 0 21840 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _3027_
timestamp 1669390400
transform 1 0 21280 0 -1 59584
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3028_
timestamp 1669390400
transform 1 0 21952 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _3029_
timestamp 1669390400
transform 1 0 21840 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _3030_
timestamp 1669390400
transform 1 0 23184 0 1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3031_
timestamp 1669390400
transform 1 0 22848 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3032_
timestamp 1669390400
transform 1 0 22960 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3033_
timestamp 1669390400
transform 1 0 23520 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3034_
timestamp 1669390400
transform -1 0 39984 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3035_
timestamp 1669390400
transform -1 0 28896 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _3036_
timestamp 1669390400
transform -1 0 28784 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3037_
timestamp 1669390400
transform -1 0 27664 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3038_
timestamp 1669390400
transform -1 0 21840 0 1 3136
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _3039_
timestamp 1669390400
transform 1 0 28896 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _3040_
timestamp 1669390400
transform -1 0 33712 0 1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _3041_
timestamp 1669390400
transform 1 0 31136 0 -1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3042_
timestamp 1669390400
transform 1 0 31136 0 1 3136
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3043_
timestamp 1669390400
transform -1 0 34160 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _3044_
timestamp 1669390400
transform 1 0 29008 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3045_
timestamp 1669390400
transform -1 0 30800 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _3046_
timestamp 1669390400
transform 1 0 29568 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3047_
timestamp 1669390400
transform 1 0 31024 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3048_
timestamp 1669390400
transform -1 0 31136 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3049_
timestamp 1669390400
transform 1 0 32592 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3050_
timestamp 1669390400
transform 1 0 31360 0 -1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3051_
timestamp 1669390400
transform -1 0 34160 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3052_
timestamp 1669390400
transform -1 0 30016 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _3053_
timestamp 1669390400
transform -1 0 31136 0 -1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3054_
timestamp 1669390400
transform 1 0 31472 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3055_
timestamp 1669390400
transform -1 0 32592 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _3056_
timestamp 1669390400
transform 1 0 30464 0 1 9408
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3057_
timestamp 1669390400
transform -1 0 32928 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3058_
timestamp 1669390400
transform 1 0 28336 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3059_
timestamp 1669390400
transform 1 0 29456 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3060_
timestamp 1669390400
transform -1 0 29120 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3061_
timestamp 1669390400
transform 1 0 29344 0 -1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3062_
timestamp 1669390400
transform -1 0 32032 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3063_
timestamp 1669390400
transform 1 0 32368 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3064_
timestamp 1669390400
transform 1 0 31248 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3065_
timestamp 1669390400
transform 1 0 29456 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3066_
timestamp 1669390400
transform -1 0 31584 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _3067_
timestamp 1669390400
transform -1 0 29008 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3068_
timestamp 1669390400
transform -1 0 27216 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _3069_
timestamp 1669390400
transform 1 0 25648 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _3070_
timestamp 1669390400
transform 1 0 29456 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3071_
timestamp 1669390400
transform -1 0 31472 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _3072_
timestamp 1669390400
transform 1 0 25648 0 -1 14112
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3073_
timestamp 1669390400
transform -1 0 27664 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3074_
timestamp 1669390400
transform -1 0 27104 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3075_
timestamp 1669390400
transform 1 0 26992 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3076_
timestamp 1669390400
transform -1 0 27776 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3077_
timestamp 1669390400
transform -1 0 27888 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3078_
timestamp 1669390400
transform -1 0 26768 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3079_
timestamp 1669390400
transform 1 0 27440 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3080_
timestamp 1669390400
transform 1 0 26320 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3081_
timestamp 1669390400
transform -1 0 26544 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3082_
timestamp 1669390400
transform -1 0 25312 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3083_
timestamp 1669390400
transform -1 0 28112 0 1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3084_
timestamp 1669390400
transform -1 0 27328 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _3085_
timestamp 1669390400
transform 1 0 28112 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3086_
timestamp 1669390400
transform 1 0 26320 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _3087_
timestamp 1669390400
transform -1 0 26768 0 1 18816
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3088_
timestamp 1669390400
transform -1 0 24080 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3089_
timestamp 1669390400
transform 1 0 28112 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _3090_
timestamp 1669390400
transform -1 0 27888 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3091_
timestamp 1669390400
transform 1 0 27440 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3092_
timestamp 1669390400
transform -1 0 25088 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3093_
timestamp 1669390400
transform -1 0 28112 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3094_
timestamp 1669390400
transform 1 0 25536 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3095_
timestamp 1669390400
transform -1 0 25984 0 1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3096_
timestamp 1669390400
transform -1 0 22176 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _3097_
timestamp 1669390400
transform -1 0 27216 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _3098_
timestamp 1669390400
transform 1 0 25760 0 1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3099_
timestamp 1669390400
transform -1 0 23744 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3100_
timestamp 1669390400
transform 1 0 25536 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _3101_
timestamp 1669390400
transform -1 0 24080 0 1 4704
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3102_
timestamp 1669390400
transform -1 0 22512 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3103_
timestamp 1669390400
transform -1 0 27776 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3104_
timestamp 1669390400
transform -1 0 26768 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _3105_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 26992 0 1 7840
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3106_
timestamp 1669390400
transform 1 0 25536 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3107_
timestamp 1669390400
transform -1 0 24752 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3108_
timestamp 1669390400
transform 1 0 22960 0 -1 6272
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3109_
timestamp 1669390400
transform -1 0 24864 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3110_
timestamp 1669390400
transform -1 0 25200 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3111_
timestamp 1669390400
transform -1 0 20832 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3112_
timestamp 1669390400
transform -1 0 28672 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3113_
timestamp 1669390400
transform -1 0 22176 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3114_
timestamp 1669390400
transform 1 0 24192 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _3115_
timestamp 1669390400
transform 1 0 20048 0 -1 7840
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3116_
timestamp 1669390400
transform -1 0 22176 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3117_
timestamp 1669390400
transform -1 0 23968 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3118_
timestamp 1669390400
transform -1 0 25088 0 -1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3119_
timestamp 1669390400
transform -1 0 23296 0 -1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3120_
timestamp 1669390400
transform 1 0 22624 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3121_
timestamp 1669390400
transform -1 0 23632 0 -1 7840
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3122_
timestamp 1669390400
transform 1 0 22400 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3123_
timestamp 1669390400
transform -1 0 21728 0 -1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3124_
timestamp 1669390400
transform -1 0 20160 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3125_
timestamp 1669390400
transform -1 0 25424 0 1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3126_
timestamp 1669390400
transform -1 0 24640 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3127_
timestamp 1669390400
transform -1 0 23184 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3128_
timestamp 1669390400
transform 1 0 22064 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _3129_
timestamp 1669390400
transform -1 0 24080 0 1 12544
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3130_
timestamp 1669390400
transform -1 0 21952 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3131_
timestamp 1669390400
transform -1 0 24080 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3132_
timestamp 1669390400
transform -1 0 26320 0 -1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3133_
timestamp 1669390400
transform -1 0 23408 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3134_
timestamp 1669390400
transform -1 0 23072 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3135_
timestamp 1669390400
transform -1 0 23856 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3136_
timestamp 1669390400
transform 1 0 22288 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3137_
timestamp 1669390400
transform 1 0 20496 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3138_
timestamp 1669390400
transform -1 0 22176 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _3139_
timestamp 1669390400
transform -1 0 26096 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3140_
timestamp 1669390400
transform -1 0 23184 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _3141_
timestamp 1669390400
transform 1 0 22064 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _3142_
timestamp 1669390400
transform -1 0 23184 0 -1 18816
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3143_
timestamp 1669390400
transform -1 0 22400 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3144_
timestamp 1669390400
transform -1 0 23296 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3145_
timestamp 1669390400
transform -1 0 22512 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3146_
timestamp 1669390400
transform -1 0 23296 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3147_
timestamp 1669390400
transform 1 0 21728 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3148_
timestamp 1669390400
transform -1 0 10864 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3149_
timestamp 1669390400
transform -1 0 10528 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _3150_
timestamp 1669390400
transform -1 0 10640 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3151_
timestamp 1669390400
transform 1 0 3472 0 -1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3152_
timestamp 1669390400
transform 1 0 6496 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3153_
timestamp 1669390400
transform 1 0 3360 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _3154_
timestamp 1669390400
transform 1 0 3472 0 -1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3155_
timestamp 1669390400
transform 1 0 5600 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3156_
timestamp 1669390400
transform 1 0 4144 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3157_
timestamp 1669390400
transform 1 0 4144 0 1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3158_
timestamp 1669390400
transform 1 0 3808 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3159_
timestamp 1669390400
transform 1 0 5600 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _3160_
timestamp 1669390400
transform 1 0 4480 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3161_
timestamp 1669390400
transform 1 0 5600 0 1 3136
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3162_
timestamp 1669390400
transform -1 0 7056 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3163_
timestamp 1669390400
transform 1 0 4592 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _3164_
timestamp 1669390400
transform -1 0 7056 0 1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3165_
timestamp 1669390400
transform 1 0 5712 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _3166_
timestamp 1669390400
transform 1 0 7616 0 1 7840
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _3167_
timestamp 1669390400
transform 1 0 7728 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3168_
timestamp 1669390400
transform 1 0 9632 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _3169_
timestamp 1669390400
transform 1 0 6720 0 -1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3170_
timestamp 1669390400
transform -1 0 7840 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3171_
timestamp 1669390400
transform 1 0 4816 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _3172_
timestamp 1669390400
transform 1 0 7728 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _3173_
timestamp 1669390400
transform -1 0 8736 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3174_
timestamp 1669390400
transform -1 0 6384 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3175_
timestamp 1669390400
transform -1 0 13104 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3176_
timestamp 1669390400
transform 1 0 11984 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3177_
timestamp 1669390400
transform -1 0 14112 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3178_
timestamp 1669390400
transform 1 0 13552 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3179_
timestamp 1669390400
transform -1 0 13776 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3180_
timestamp 1669390400
transform -1 0 12208 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _3181_
timestamp 1669390400
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _3182_
timestamp 1669390400
transform 1 0 12208 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3183_
timestamp 1669390400
transform -1 0 11200 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3184_
timestamp 1669390400
transform -1 0 10080 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3185_
timestamp 1669390400
transform -1 0 10864 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _3186_
timestamp 1669390400
transform -1 0 10304 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3187_
timestamp 1669390400
transform -1 0 6384 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _3188_
timestamp 1669390400
transform -1 0 11984 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3189_
timestamp 1669390400
transform -1 0 16128 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3190_
timestamp 1669390400
transform -1 0 15344 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _3191_
timestamp 1669390400
transform -1 0 18256 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3192_
timestamp 1669390400
transform -1 0 17584 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3193_
timestamp 1669390400
transform -1 0 16800 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _3194_
timestamp 1669390400
transform 1 0 17696 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3195_
timestamp 1669390400
transform -1 0 19152 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3196_
timestamp 1669390400
transform -1 0 17136 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3197_
timestamp 1669390400
transform 1 0 19376 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _3198_
timestamp 1669390400
transform 1 0 18480 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _3199_
timestamp 1669390400
transform -1 0 22960 0 -1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _3200_
timestamp 1669390400
transform -1 0 19936 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _3201_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 17584 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _3202_
timestamp 1669390400
transform 1 0 9296 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  _3203_ Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 10080 0 -1 6272
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _3204_
timestamp 1669390400
transform -1 0 17136 0 -1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _3205_
timestamp 1669390400
transform 1 0 9296 0 1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _3206_
timestamp 1669390400
transform 1 0 13328 0 -1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _3207_
timestamp 1669390400
transform 1 0 10528 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _3208_
timestamp 1669390400
transform 1 0 15456 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _3209_
timestamp 1669390400
transform 1 0 15344 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _3210_
timestamp 1669390400
transform 1 0 17584 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  _3211_
timestamp 1669390400
transform 1 0 14784 0 1 7840
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  _3212_
timestamp 1669390400
transform 1 0 15008 0 1 6272
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _3213_
timestamp 1669390400
transform 1 0 15232 0 1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  _3214_
timestamp 1669390400
transform 1 0 15344 0 1 10976
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _3215_
timestamp 1669390400
transform 1 0 15344 0 1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _3216_
timestamp 1669390400
transform 1 0 15344 0 1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _3217_
timestamp 1669390400
transform 1 0 9296 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _3218_
timestamp 1669390400
transform -1 0 9184 0 -1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _3219_
timestamp 1669390400
transform 1 0 5600 0 1 12544
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _3220_
timestamp 1669390400
transform 1 0 5264 0 -1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _3221_
timestamp 1669390400
transform 1 0 5376 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _3222_
timestamp 1669390400
transform 1 0 5376 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _3223_
timestamp 1669390400
transform 1 0 9632 0 -1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _3224_
timestamp 1669390400
transform 1 0 5152 0 -1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _3225_
timestamp 1669390400
transform 1 0 5040 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _3226_
timestamp 1669390400
transform 1 0 9296 0 1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _3227_
timestamp 1669390400
transform 1 0 9296 0 1 14112
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _3228_
timestamp 1669390400
transform 1 0 8064 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _3229_
timestamp 1669390400
transform 1 0 5376 0 -1 17248
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_2  _3230_
timestamp 1669390400
transform -1 0 15120 0 -1 17248
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _3231_
timestamp 1669390400
transform 1 0 13328 0 -1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _3232_
timestamp 1669390400
transform 1 0 15344 0 1 15680
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _3233_
timestamp 1669390400
transform 1 0 15344 0 1 18816
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 11536 0 -1 12544
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1669390400
transform 1 0 7504 0 1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1669390400
transform 1 0 11424 0 -1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1669390400
transform -1 0 9184 0 -1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1669390400
transform 1 0 11424 0 -1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  fanout9
timestamp 1669390400
transform 1 0 18480 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  fanout10
timestamp 1669390400
transform 1 0 18368 0 -1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  fanout11 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 20944 0 1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout12 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 16016 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input1 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 30240 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input2
timestamp 1669390400
transform 1 0 38864 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input3
timestamp 1669390400
transform -1 0 48272 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input4
timestamp 1669390400
transform -1 0 55888 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input5 Desktop/EF/FullFlow/pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 13440 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output6
timestamp 1669390400
transform 1 0 50288 0 1 59584
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output7
timestamp 1669390400
transform -1 0 11760 0 1 59584
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output8
timestamp 1669390400
transform 1 0 30240 0 1 59584
box -86 -86 1654 870
<< labels >>
flabel metal2 s 4256 0 4368 800 0 FreeSans 448 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 30128 0 30240 800 0 FreeSans 448 90 0 0 divSel[0]
port 1 nsew signal input
flabel metal2 s 38752 0 38864 800 0 FreeSans 448 90 0 0 divSel[1]
port 2 nsew signal input
flabel metal2 s 47376 0 47488 800 0 FreeSans 448 90 0 0 divSel[2]
port 3 nsew signal input
flabel metal2 s 56000 0 56112 800 0 FreeSans 448 90 0 0 divSel[3]
port 4 nsew signal input
flabel metal2 s 21504 0 21616 800 0 FreeSans 448 90 0 0 enable
port 5 nsew signal input
flabel metal2 s 50176 63181 50288 63981 0 FreeSans 448 90 0 0 qcomplex
port 6 nsew signal tristate
flabel metal2 s 10080 63181 10192 63981 0 FreeSans 448 90 0 0 qcos
port 7 nsew signal tristate
flabel metal2 s 30128 63181 30240 63981 0 FreeSans 448 90 0 0 qsin
port 8 nsew signal tristate
flabel metal2 s 12880 0 12992 800 0 FreeSans 448 90 0 0 rst
port 9 nsew signal input
flabel metal4 s 4448 3076 4768 60428 0 FreeSans 1280 90 0 0 vdd
port 10 nsew power bidirectional
flabel metal4 s 35168 3076 35488 60428 0 FreeSans 1280 90 0 0 vdd
port 10 nsew power bidirectional
flabel metal4 s 19808 3076 20128 60428 0 FreeSans 1280 90 0 0 vss
port 11 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 60428 0 FreeSans 1280 90 0 0 vss
port 11 nsew ground bidirectional
rlabel metal1 30184 60368 30184 60368 0 vdd
rlabel metal1 30184 59584 30184 59584 0 vss
rlabel metal2 18200 5376 18200 5376 0 _0000_
rlabel metal2 15400 7392 15400 7392 0 _0001_
rlabel metal2 15736 7336 15736 7336 0 _0002_
rlabel metal2 15960 10248 15960 10248 0 _0003_
rlabel metal2 16072 11816 16072 11816 0 _0004_
rlabel metal2 16072 13608 16072 13608 0 _0005_
rlabel metal3 17024 14504 17024 14504 0 _0006_
rlabel metal2 9912 8316 9912 8316 0 _0007_
rlabel metal2 7000 11704 7000 11704 0 _0008_
rlabel metal2 6104 12096 6104 12096 0 _0009_
rlabel metal2 5992 9296 5992 9296 0 _0010_
rlabel metal2 14504 4872 14504 4872 0 _0011_
rlabel metal2 6216 4312 6216 4312 0 _0012_
rlabel metal2 6160 5880 6160 5880 0 _0013_
rlabel metal2 10248 7924 10248 7924 0 _0014_
rlabel metal2 5544 17192 5544 17192 0 _0015_
rlabel metal2 5824 21672 5824 21672 0 _0016_
rlabel metal3 11088 22120 11088 22120 0 _0017_
rlabel metal2 10024 14840 10024 14840 0 _0018_
rlabel metal2 9128 16072 9128 16072 0 _0019_
rlabel metal2 5936 20216 5936 20216 0 _0020_
rlabel metal2 14672 16856 14672 16856 0 _0021_
rlabel metal2 14280 5432 14280 5432 0 _0022_
rlabel metal2 14056 19152 14056 19152 0 _0023_
rlabel metal2 16240 16072 16240 16072 0 _0024_
rlabel metal2 16128 19208 16128 19208 0 _0025_
rlabel metal2 18648 8792 18648 8792 0 _0026_
rlabel metal2 13104 9240 13104 9240 0 _0027_
rlabel metal3 23464 11704 23464 11704 0 _0028_
rlabel metal2 24808 14000 24808 14000 0 _0029_
rlabel metal2 16184 18032 16184 18032 0 _0030_
rlabel metal2 21672 5880 21672 5880 0 _0031_
rlabel metal2 22008 5936 22008 5936 0 _0032_
rlabel metal2 43848 14504 43848 14504 0 _0033_
rlabel metal3 45640 14616 45640 14616 0 _0034_
rlabel metal3 47880 15176 47880 15176 0 _0035_
rlabel metal2 52696 14560 52696 14560 0 _0036_
rlabel metal3 49224 14616 49224 14616 0 _0037_
rlabel metal3 50680 12936 50680 12936 0 _0038_
rlabel metal2 35672 15904 35672 15904 0 _0039_
rlabel metal2 36176 15288 36176 15288 0 _0040_
rlabel metal2 35896 15568 35896 15568 0 _0041_
rlabel metal2 30856 19040 30856 19040 0 _0042_
rlabel metal2 6776 30576 6776 30576 0 _0043_
rlabel metal3 33824 17640 33824 17640 0 _0044_
rlabel metal2 36008 15400 36008 15400 0 _0045_
rlabel metal2 37352 15148 37352 15148 0 _0046_
rlabel metal2 39592 14112 39592 14112 0 _0047_
rlabel metal2 36344 15008 36344 15008 0 _0048_
rlabel metal2 46424 13272 46424 13272 0 _0049_
rlabel metal2 46088 14000 46088 14000 0 _0050_
rlabel metal2 47432 12992 47432 12992 0 _0051_
rlabel metal2 47656 12936 47656 12936 0 _0052_
rlabel metal2 47096 12264 47096 12264 0 _0053_
rlabel metal3 6608 23800 6608 23800 0 _0054_
rlabel metal3 48720 12376 48720 12376 0 _0055_
rlabel metal3 48328 13048 48328 13048 0 _0056_
rlabel metal2 51352 12768 51352 12768 0 _0057_
rlabel metal2 49672 12600 49672 12600 0 _0058_
rlabel metal2 51856 13608 51856 13608 0 _0059_
rlabel metal3 51408 14728 51408 14728 0 _0060_
rlabel metal2 52248 15008 52248 15008 0 _0061_
rlabel metal2 52752 13160 52752 13160 0 _0062_
rlabel metal2 52584 15624 52584 15624 0 _0063_
rlabel metal2 54488 14784 54488 14784 0 _0064_
rlabel metal2 4144 45192 4144 45192 0 _0065_
rlabel metal2 53704 16520 53704 16520 0 _0066_
rlabel metal2 52808 16240 52808 16240 0 _0067_
rlabel metal3 54684 16968 54684 16968 0 _0068_
rlabel metal2 56056 19936 56056 19936 0 _0069_
rlabel metal3 57120 18648 57120 18648 0 _0070_
rlabel metal3 57176 15288 57176 15288 0 _0071_
rlabel metal2 57512 15904 57512 15904 0 _0072_
rlabel metal2 43736 10920 43736 10920 0 _0073_
rlabel metal3 45192 11368 45192 11368 0 _0074_
rlabel metal2 46368 11144 46368 11144 0 _0075_
rlabel metal2 12880 46872 12880 46872 0 _0076_
rlabel metal3 46480 11256 46480 11256 0 _0077_
rlabel metal2 49560 10920 49560 10920 0 _0078_
rlabel metal2 51688 10136 51688 10136 0 _0079_
rlabel metal2 50568 7672 50568 7672 0 _0080_
rlabel metal2 46648 10304 46648 10304 0 _0081_
rlabel metal2 47432 9856 47432 9856 0 _0082_
rlabel metal3 31360 17416 31360 17416 0 _0083_
rlabel metal3 45864 9800 45864 9800 0 _0084_
rlabel metal3 44968 10024 44968 10024 0 _0085_
rlabel metal3 44240 9128 44240 9128 0 _0086_
rlabel metal2 1848 26992 1848 26992 0 _0087_
rlabel metal2 44632 8316 44632 8316 0 _0088_
rlabel metal2 44464 9128 44464 9128 0 _0089_
rlabel metal3 45752 9128 45752 9128 0 _0090_
rlabel metal2 38360 14784 38360 14784 0 _0091_
rlabel metal2 46032 8008 46032 8008 0 _0092_
rlabel metal2 47096 7952 47096 7952 0 _0093_
rlabel metal3 46928 9016 46928 9016 0 _0094_
rlabel metal3 48720 9128 48720 9128 0 _0095_
rlabel metal2 49560 9632 49560 9632 0 _0096_
rlabel metal3 50792 8008 50792 8008 0 _0097_
rlabel metal2 4200 22568 4200 22568 0 _0098_
rlabel metal2 50008 7924 50008 7924 0 _0099_
rlabel metal2 51072 8232 51072 8232 0 _0100_
rlabel metal2 53144 10920 53144 10920 0 _0101_
rlabel metal2 54040 10360 54040 10360 0 _0102_
rlabel metal2 55384 11564 55384 11564 0 _0103_
rlabel metal2 54936 11648 54936 11648 0 _0104_
rlabel metal2 56280 11984 56280 11984 0 _0105_
rlabel metal2 53480 8288 53480 8288 0 _0106_
rlabel metal2 34776 6720 34776 6720 0 _0107_
rlabel metal3 33488 13608 33488 13608 0 _0108_
rlabel metal3 13552 48216 13552 48216 0 _0109_
rlabel metal3 33096 13720 33096 13720 0 _0110_
rlabel metal3 33936 6664 33936 6664 0 _0111_
rlabel metal2 35112 7560 35112 7560 0 _0112_
rlabel metal2 42560 8232 42560 8232 0 _0113_
rlabel metal2 42280 9296 42280 9296 0 _0114_
rlabel metal2 42952 7784 42952 7784 0 _0115_
rlabel metal2 42504 6664 42504 6664 0 _0116_
rlabel metal2 34664 7000 34664 7000 0 _0117_
rlabel metal2 36176 5880 36176 5880 0 _0118_
rlabel metal2 45360 6104 45360 6104 0 _0119_
rlabel metal2 4144 26264 4144 26264 0 _0120_
rlabel metal2 45192 5768 45192 5768 0 _0121_
rlabel metal3 46704 5992 46704 5992 0 _0122_
rlabel metal2 44520 4648 44520 4648 0 _0123_
rlabel metal2 44800 4984 44800 4984 0 _0124_
rlabel metal3 46592 5880 46592 5880 0 _0125_
rlabel metal2 47880 7000 47880 7000 0 _0126_
rlabel metal2 53816 6720 53816 6720 0 _0127_
rlabel metal2 53144 7840 53144 7840 0 _0128_
rlabel metal2 54488 8036 54488 8036 0 _0129_
rlabel metal2 52808 9408 52808 9408 0 _0130_
rlabel metal2 2968 35392 2968 35392 0 _0131_
rlabel metal3 53704 8232 53704 8232 0 _0132_
rlabel metal2 55160 9296 55160 9296 0 _0133_
rlabel metal3 54040 9128 54040 9128 0 _0134_
rlabel metal2 55272 10080 55272 10080 0 _0135_
rlabel metal3 56840 12264 56840 12264 0 _0136_
rlabel metal2 57064 11760 57064 11760 0 _0137_
rlabel metal2 56504 11648 56504 11648 0 _0138_
rlabel metal2 57512 9520 57512 9520 0 _0139_
rlabel metal2 34216 12208 34216 12208 0 _0140_
rlabel metal2 33880 11648 33880 11648 0 _0141_
rlabel metal2 2352 31192 2352 31192 0 _0142_
rlabel metal2 35000 5040 35000 5040 0 _0143_
rlabel metal2 35840 4312 35840 4312 0 _0144_
rlabel metal2 34776 5432 34776 5432 0 _0145_
rlabel metal3 36232 4200 36232 4200 0 _0146_
rlabel metal2 40264 12432 40264 12432 0 _0147_
rlabel metal2 39032 11760 39032 11760 0 _0148_
rlabel metal2 38192 5096 38192 5096 0 _0149_
rlabel metal3 37072 5096 37072 5096 0 _0150_
rlabel metal3 36904 4312 36904 4312 0 _0151_
rlabel metal2 37464 5040 37464 5040 0 _0152_
rlabel metal2 4704 24024 4704 24024 0 _0153_
rlabel metal2 38808 4032 38808 4032 0 _0154_
rlabel metal2 42056 4760 42056 4760 0 _0155_
rlabel metal3 38472 4088 38472 4088 0 _0156_
rlabel metal2 41048 3808 41048 3808 0 _0157_
rlabel metal2 41608 3416 41608 3416 0 _0158_
rlabel metal2 44408 5320 44408 5320 0 _0159_
rlabel metal3 44296 5880 44296 5880 0 _0160_
rlabel metal3 42224 4984 42224 4984 0 _0161_
rlabel metal2 40488 9856 40488 9856 0 _0162_
rlabel metal3 34888 9800 34888 9800 0 _0163_
rlabel metal3 10976 49560 10976 49560 0 _0164_
rlabel metal3 36288 9688 36288 9688 0 _0165_
rlabel metal2 37856 8232 37856 8232 0 _0166_
rlabel metal2 35056 11144 35056 11144 0 _0167_
rlabel metal2 38136 8400 38136 8400 0 _0168_
rlabel metal2 39648 5096 39648 5096 0 _0169_
rlabel metal3 41832 12376 41832 12376 0 _0170_
rlabel metal3 41216 9688 41216 9688 0 _0171_
rlabel metal3 40320 8232 40320 8232 0 _0172_
rlabel metal2 41048 7728 41048 7728 0 _0173_
rlabel metal2 39648 7672 39648 7672 0 _0174_
rlabel metal3 2184 45080 2184 45080 0 _0175_
rlabel metal2 39256 5432 39256 5432 0 _0176_
rlabel metal2 41720 4984 41720 4984 0 _0177_
rlabel metal3 40432 4536 40432 4536 0 _0178_
rlabel metal2 41496 5096 41496 5096 0 _0179_
rlabel metal2 41384 9800 41384 9800 0 _0180_
rlabel metal2 41608 6384 41608 6384 0 _0181_
rlabel metal2 37520 10584 37520 10584 0 _0182_
rlabel metal2 37744 10584 37744 10584 0 _0183_
rlabel metal2 39144 8316 39144 8316 0 _0184_
rlabel metal3 38360 9016 38360 9016 0 _0185_
rlabel metal2 10808 46480 10808 46480 0 _0186_
rlabel metal2 39088 9128 39088 9128 0 _0187_
rlabel metal2 39592 8736 39592 8736 0 _0188_
rlabel metal3 40264 8008 40264 8008 0 _0189_
rlabel metal3 41216 5320 41216 5320 0 _0190_
rlabel metal2 44184 5376 44184 5376 0 _0191_
rlabel metal2 43064 5376 43064 5376 0 _0192_
rlabel metal2 43848 5544 43848 5544 0 _0193_
rlabel metal2 48776 5712 48776 5712 0 _0194_
rlabel metal2 47320 5432 47320 5432 0 _0195_
rlabel metal2 48216 5040 48216 5040 0 _0196_
rlabel metal2 11480 47096 11480 47096 0 _0197_
rlabel metal2 48104 4760 48104 4760 0 _0198_
rlabel metal2 49672 6496 49672 6496 0 _0199_
rlabel metal2 55048 7672 55048 7672 0 _0200_
rlabel metal2 53536 7672 53536 7672 0 _0201_
rlabel metal2 55664 7448 55664 7448 0 _0202_
rlabel metal2 56056 10192 56056 10192 0 _0203_
rlabel metal2 57456 16632 57456 16632 0 _0204_
rlabel metal2 56392 21448 56392 21448 0 _0205_
rlabel metal2 57400 18200 57400 18200 0 _0206_
rlabel metal2 58296 17640 58296 17640 0 _0207_
rlabel metal3 16856 48776 16856 48776 0 _0208_
rlabel metal2 58520 51240 58520 51240 0 _0209_
rlabel metal2 55048 44016 55048 44016 0 _0210_
rlabel metal2 54712 42000 54712 42000 0 _0211_
rlabel metal3 56560 50568 56560 50568 0 _0212_
rlabel metal2 58184 49280 58184 49280 0 _0213_
rlabel metal3 57120 47432 57120 47432 0 _0214_
rlabel metal2 57848 50232 57848 50232 0 _0215_
rlabel metal2 57848 50792 57848 50792 0 _0216_
rlabel metal2 52920 55888 52920 55888 0 _0217_
rlabel metal3 44968 47320 44968 47320 0 _0218_
rlabel metal2 15176 49672 15176 49672 0 _0219_
rlabel metal2 44520 45528 44520 45528 0 _0220_
rlabel metal2 45192 47488 45192 47488 0 _0221_
rlabel metal3 45024 47432 45024 47432 0 _0222_
rlabel metal2 46872 47768 46872 47768 0 _0223_
rlabel metal3 45136 46760 45136 46760 0 _0224_
rlabel metal2 46592 47320 46592 47320 0 _0225_
rlabel metal2 46088 47488 46088 47488 0 _0226_
rlabel metal2 45808 51464 45808 51464 0 _0227_
rlabel metal2 43064 48216 43064 48216 0 _0228_
rlabel metal2 41496 45360 41496 45360 0 _0229_
rlabel metal2 17752 45752 17752 45752 0 _0230_
rlabel metal3 40712 40152 40712 40152 0 _0231_
rlabel metal3 42504 45864 42504 45864 0 _0232_
rlabel metal3 41216 47320 41216 47320 0 _0233_
rlabel metal2 39592 46144 39592 46144 0 _0234_
rlabel metal2 36456 41216 36456 41216 0 _0235_
rlabel metal3 37296 45864 37296 45864 0 _0236_
rlabel metal3 37072 45976 37072 45976 0 _0237_
rlabel metal2 39312 46088 39312 46088 0 _0238_
rlabel metal3 41328 47432 41328 47432 0 _0239_
rlabel metal2 43344 48104 43344 48104 0 _0240_
rlabel metal2 14504 47768 14504 47768 0 _0241_
rlabel metal3 44128 48776 44128 48776 0 _0242_
rlabel metal2 46424 49504 46424 49504 0 _0243_
rlabel metal2 46760 49000 46760 49000 0 _0244_
rlabel metal3 45248 49000 45248 49000 0 _0245_
rlabel metal3 45360 50344 45360 50344 0 _0246_
rlabel metal2 43568 49560 43568 49560 0 _0247_
rlabel metal2 42952 51072 42952 51072 0 _0248_
rlabel metal2 39704 46704 39704 46704 0 _0249_
rlabel metal3 41440 48776 41440 48776 0 _0250_
rlabel metal2 40488 41552 40488 41552 0 _0251_
rlabel metal2 8064 26600 8064 26600 0 _0252_
rlabel metal2 42784 41720 42784 41720 0 _0253_
rlabel metal2 39704 41496 39704 41496 0 _0254_
rlabel metal3 38808 41944 38808 41944 0 _0255_
rlabel metal2 39816 42224 39816 42224 0 _0256_
rlabel metal2 39592 47544 39592 47544 0 _0257_
rlabel metal2 38136 47544 38136 47544 0 _0258_
rlabel metal3 36344 46648 36344 46648 0 _0259_
rlabel metal2 35896 44576 35896 44576 0 _0260_
rlabel metal2 36176 47432 36176 47432 0 _0261_
rlabel metal2 35672 47544 35672 47544 0 _0262_
rlabel metal3 18144 34776 18144 34776 0 _0263_
rlabel metal3 37184 48216 37184 48216 0 _0264_
rlabel metal3 39256 48104 39256 48104 0 _0265_
rlabel metal3 41160 48888 41160 48888 0 _0266_
rlabel via2 42616 50792 42616 50792 0 _0267_
rlabel metal3 46088 51352 46088 51352 0 _0268_
rlabel metal2 47992 52472 47992 52472 0 _0269_
rlabel metal3 49280 46872 49280 46872 0 _0270_
rlabel metal2 49672 47488 49672 47488 0 _0271_
rlabel metal2 49504 48440 49504 48440 0 _0272_
rlabel metal3 49168 44296 49168 44296 0 _0273_
rlabel metal3 16240 48216 16240 48216 0 _0274_
rlabel metal3 49896 49784 49896 49784 0 _0275_
rlabel metal2 48440 49392 48440 49392 0 _0276_
rlabel metal2 49784 49000 49784 49000 0 _0277_
rlabel metal2 49000 49280 49000 49280 0 _0278_
rlabel metal2 49896 50344 49896 50344 0 _0279_
rlabel metal2 49448 53872 49448 53872 0 _0280_
rlabel metal2 46312 50960 46312 50960 0 _0281_
rlabel metal2 46088 51184 46088 51184 0 _0282_
rlabel metal2 46760 51352 46760 51352 0 _0283_
rlabel metal2 46144 53704 46144 53704 0 _0284_
rlabel metal2 3248 37240 3248 37240 0 _0285_
rlabel metal2 43176 50008 43176 50008 0 _0286_
rlabel metal2 42224 49224 42224 49224 0 _0287_
rlabel metal2 41832 50904 41832 50904 0 _0288_
rlabel metal2 41832 53368 41832 53368 0 _0289_
rlabel metal2 40040 42000 40040 42000 0 _0290_
rlabel metal2 39144 50232 39144 50232 0 _0291_
rlabel metal2 39200 47432 39200 47432 0 _0292_
rlabel metal2 39144 50512 39144 50512 0 _0293_
rlabel metal3 36848 51352 36848 51352 0 _0294_
rlabel metal2 39928 50148 39928 50148 0 _0295_
rlabel metal2 16296 47768 16296 47768 0 _0296_
rlabel metal2 37688 51072 37688 51072 0 _0297_
rlabel metal3 37352 50568 37352 50568 0 _0298_
rlabel metal2 36176 49000 36176 49000 0 _0299_
rlabel metal3 33432 48216 33432 48216 0 _0300_
rlabel metal2 33936 46424 33936 46424 0 _0301_
rlabel metal2 33992 49840 33992 49840 0 _0302_
rlabel metal2 34552 48720 34552 48720 0 _0303_
rlabel metal3 35224 49672 35224 49672 0 _0304_
rlabel metal3 37296 50680 37296 50680 0 _0305_
rlabel metal2 39368 51072 39368 51072 0 _0306_
rlabel metal2 25816 38864 25816 38864 0 _0307_
rlabel metal2 39480 51520 39480 51520 0 _0308_
rlabel metal2 41720 53760 41720 53760 0 _0309_
rlabel metal3 45360 53816 45360 53816 0 _0310_
rlabel metal3 49336 53704 49336 53704 0 _0311_
rlabel metal2 51296 56168 51296 56168 0 _0312_
rlabel metal2 46424 55776 46424 55776 0 _0313_
rlabel metal2 36568 52248 36568 52248 0 _0314_
rlabel metal2 36176 50008 36176 50008 0 _0315_
rlabel metal2 36680 52192 36680 52192 0 _0316_
rlabel metal2 33432 50512 33432 50512 0 _0317_
rlabel metal2 32536 50736 32536 50736 0 _0318_
rlabel metal3 33656 50456 33656 50456 0 _0319_
rlabel metal2 32424 51184 32424 51184 0 _0320_
rlabel metal2 29960 50624 29960 50624 0 _0321_
rlabel metal2 30184 51016 30184 51016 0 _0322_
rlabel metal2 30296 52192 30296 52192 0 _0323_
rlabel metal2 30744 51464 30744 51464 0 _0324_
rlabel metal3 31500 51240 31500 51240 0 _0325_
rlabel metal3 33712 51240 33712 51240 0 _0326_
rlabel metal2 35112 52920 35112 52920 0 _0327_
rlabel metal2 38360 53368 38360 53368 0 _0328_
rlabel metal2 1960 32816 1960 32816 0 _0329_
rlabel metal2 39704 51576 39704 51576 0 _0330_
rlabel metal2 39704 54040 39704 54040 0 _0331_
rlabel metal2 41608 54208 41608 54208 0 _0332_
rlabel metal2 42616 53200 42616 53200 0 _0333_
rlabel metal2 43288 53480 43288 53480 0 _0334_
rlabel metal3 42280 54600 42280 54600 0 _0335_
rlabel metal2 46312 56224 46312 56224 0 _0336_
rlabel metal2 51576 57848 51576 57848 0 _0337_
rlabel metal2 50960 58520 50960 58520 0 _0338_
rlabel metal2 51352 57120 51352 57120 0 _0339_
rlabel metal3 19936 48888 19936 48888 0 _0340_
rlabel metal2 52640 51912 52640 51912 0 _0341_
rlabel metal3 52976 45192 52976 45192 0 _0342_
rlabel metal2 51800 50400 51800 50400 0 _0343_
rlabel metal2 51576 51016 51576 51016 0 _0344_
rlabel metal2 52472 52080 52472 52080 0 _0345_
rlabel metal3 53424 54600 53424 54600 0 _0346_
rlabel metal2 51800 52416 51800 52416 0 _0347_
rlabel metal2 51352 53368 51352 53368 0 _0348_
rlabel metal2 52248 53760 52248 53760 0 _0349_
rlabel metal2 52192 54712 52192 54712 0 _0350_
rlabel metal2 18088 49392 18088 49392 0 _0351_
rlabel metal2 52024 57008 52024 57008 0 _0352_
rlabel metal2 53032 53312 53032 53312 0 _0353_
rlabel metal2 50456 58072 50456 58072 0 _0354_
rlabel metal3 48832 58408 48832 58408 0 _0355_
rlabel metal2 48440 56560 48440 56560 0 _0356_
rlabel metal3 46816 58520 46816 58520 0 _0357_
rlabel metal2 44352 58632 44352 58632 0 _0358_
rlabel metal2 33824 54376 33824 54376 0 _0359_
rlabel metal3 33880 54264 33880 54264 0 _0360_
rlabel metal3 33936 50792 33936 50792 0 _0361_
rlabel metal3 19488 49112 19488 49112 0 _0362_
rlabel metal2 33768 51576 33768 51576 0 _0363_
rlabel metal2 32592 53592 32592 53592 0 _0364_
rlabel metal2 29176 52584 29176 52584 0 _0365_
rlabel metal2 28672 54488 28672 54488 0 _0366_
rlabel metal3 27720 54488 27720 54488 0 _0367_
rlabel metal3 29624 54488 29624 54488 0 _0368_
rlabel metal2 31304 51184 31304 51184 0 _0369_
rlabel metal3 27496 52024 27496 52024 0 _0370_
rlabel metal3 27440 50568 27440 50568 0 _0371_
rlabel metal2 26992 49672 26992 49672 0 _0372_
rlabel metal2 23352 46312 23352 46312 0 _0373_
rlabel metal2 27496 51632 27496 51632 0 _0374_
rlabel metal3 29008 52136 29008 52136 0 _0375_
rlabel metal3 29792 53704 29792 53704 0 _0376_
rlabel metal2 32536 54152 32536 54152 0 _0377_
rlabel metal3 32816 55272 32816 55272 0 _0378_
rlabel metal3 35000 55272 35000 55272 0 _0379_
rlabel metal2 35616 53704 35616 53704 0 _0380_
rlabel metal2 36456 54040 36456 54040 0 _0381_
rlabel metal2 36008 54600 36008 54600 0 _0382_
rlabel metal2 37912 55216 37912 55216 0 _0383_
rlabel metal2 24360 45920 24360 45920 0 _0384_
rlabel metal2 39368 54824 39368 54824 0 _0385_
rlabel metal2 39816 54936 39816 54936 0 _0386_
rlabel metal3 40096 55272 40096 55272 0 _0387_
rlabel metal2 41552 57512 41552 57512 0 _0388_
rlabel metal2 27608 54488 27608 54488 0 _0389_
rlabel metal2 29848 54376 29848 54376 0 _0390_
rlabel metal2 30184 53256 30184 53256 0 _0391_
rlabel metal2 26040 54544 26040 54544 0 _0392_
rlabel metal2 20552 53200 20552 53200 0 _0393_
rlabel metal2 19656 53760 19656 53760 0 _0394_
rlabel metal2 18984 21616 18984 21616 0 _0395_
rlabel metal2 19544 54544 19544 54544 0 _0396_
rlabel metal2 29344 50568 29344 50568 0 _0397_
rlabel metal3 19376 55272 19376 55272 0 _0398_
rlabel metal2 26768 50008 26768 50008 0 _0399_
rlabel metal2 27384 52304 27384 52304 0 _0400_
rlabel metal3 23128 55384 23128 55384 0 _0401_
rlabel metal2 27160 54936 27160 54936 0 _0402_
rlabel metal3 29344 56728 29344 56728 0 _0403_
rlabel metal2 32760 54488 32760 54488 0 _0404_
rlabel metal3 29680 56840 29680 56840 0 _0405_
rlabel metal3 19880 26264 19880 26264 0 _0406_
rlabel metal2 29512 58016 29512 58016 0 _0407_
rlabel metal2 29736 57008 29736 57008 0 _0408_
rlabel metal3 37072 57400 37072 57400 0 _0409_
rlabel metal2 36456 58184 36456 58184 0 _0410_
rlabel metal2 38136 59136 38136 59136 0 _0411_
rlabel metal3 43792 59304 43792 59304 0 _0412_
rlabel metal3 45192 59192 45192 59192 0 _0413_
rlabel metal2 35672 58296 35672 58296 0 _0414_
rlabel metal2 39424 59080 39424 59080 0 _0415_
rlabel metal3 38164 58296 38164 58296 0 _0416_
rlabel metal2 1848 22064 1848 22064 0 _0417_
rlabel metal3 37128 58408 37128 58408 0 _0418_
rlabel metal2 35000 58520 35000 58520 0 _0419_
rlabel metal2 34216 59696 34216 59696 0 _0420_
rlabel metal2 28616 58072 28616 58072 0 _0421_
rlabel metal2 26768 54712 26768 54712 0 _0422_
rlabel metal3 26208 58408 26208 58408 0 _0423_
rlabel metal2 14056 57512 14056 57512 0 _0424_
rlabel metal2 12488 54824 12488 54824 0 _0425_
rlabel metal4 20216 52472 20216 52472 0 _0426_
rlabel metal2 12656 58296 12656 58296 0 _0427_
rlabel metal2 11816 21392 11816 21392 0 _0428_
rlabel metal2 19208 58352 19208 58352 0 _0429_
rlabel metal3 19824 55832 19824 55832 0 _0430_
rlabel metal2 19208 56840 19208 56840 0 _0431_
rlabel metal2 18984 56056 18984 56056 0 _0432_
rlabel metal2 19096 57736 19096 57736 0 _0433_
rlabel metal3 22176 58296 22176 58296 0 _0434_
rlabel metal2 27832 58016 27832 58016 0 _0435_
rlabel metal2 28168 58856 28168 58856 0 _0436_
rlabel metal3 30464 59304 30464 59304 0 _0437_
rlabel metal2 28728 58856 28728 58856 0 _0438_
rlabel metal2 12152 36904 12152 36904 0 _0439_
rlabel metal2 29960 58744 29960 58744 0 _0440_
rlabel metal3 29400 58632 29400 58632 0 _0441_
rlabel metal2 32536 58800 32536 58800 0 _0442_
rlabel metal3 34272 59192 34272 59192 0 _0443_
rlabel metal3 35448 57064 35448 57064 0 _0444_
rlabel metal2 53816 55300 53816 55300 0 _0445_
rlabel metal2 54152 18704 54152 18704 0 _0446_
rlabel metal3 55216 15288 55216 15288 0 _0447_
rlabel metal2 55272 16408 55272 16408 0 _0448_
rlabel metal2 55048 16464 55048 16464 0 _0449_
rlabel metal2 17024 47544 17024 47544 0 _0450_
rlabel metal3 56728 16968 56728 16968 0 _0451_
rlabel metal2 55552 14616 55552 14616 0 _0452_
rlabel metal2 56448 12152 56448 12152 0 _0453_
rlabel metal2 56616 13160 56616 13160 0 _0454_
rlabel metal2 56616 8372 56616 8372 0 _0455_
rlabel metal3 51856 6440 51856 6440 0 _0456_
rlabel metal2 55944 7952 55944 7952 0 _0457_
rlabel metal2 58520 13104 58520 13104 0 _0458_
rlabel metal2 55720 16856 55720 16856 0 _0459_
rlabel metal2 54992 41272 54992 41272 0 _0460_
rlabel metal3 21056 49000 21056 49000 0 _0461_
rlabel metal2 56448 49560 56448 49560 0 _0462_
rlabel metal3 54880 55048 54880 55048 0 _0463_
rlabel metal2 52416 56168 52416 56168 0 _0464_
rlabel metal2 53816 57400 53816 57400 0 _0465_
rlabel metal2 43512 58296 43512 58296 0 _0466_
rlabel metal2 34776 58688 34776 58688 0 _0467_
rlabel metal3 34776 58408 34776 58408 0 _0468_
rlabel metal2 35616 57064 35616 57064 0 _0469_
rlabel metal3 41104 57848 41104 57848 0 _0470_
rlabel metal2 38584 58800 38584 58800 0 _0471_
rlabel metal2 23128 48832 23128 48832 0 _0472_
rlabel metal2 38136 58016 38136 58016 0 _0473_
rlabel metal3 37520 56728 37520 56728 0 _0474_
rlabel metal2 44184 59080 44184 59080 0 _0475_
rlabel metal3 43904 57848 43904 57848 0 _0476_
rlabel metal2 38472 57344 38472 57344 0 _0477_
rlabel metal2 38360 57176 38360 57176 0 _0478_
rlabel metal3 49896 48776 49896 48776 0 _0479_
rlabel metal2 53480 55048 53480 55048 0 _0480_
rlabel metal3 53984 54488 53984 54488 0 _0481_
rlabel metal2 53592 54040 53592 54040 0 _0482_
rlabel metal2 24920 45024 24920 45024 0 _0483_
rlabel metal2 53480 53816 53480 53816 0 _0484_
rlabel metal3 51296 57512 51296 57512 0 _0485_
rlabel metal2 50344 56728 50344 56728 0 _0486_
rlabel metal2 48328 54824 48328 54824 0 _0487_
rlabel metal2 47992 54936 47992 54936 0 _0488_
rlabel metal2 55384 47488 55384 47488 0 _0489_
rlabel metal2 55720 47824 55720 47824 0 _0490_
rlabel metal3 53648 48216 53648 48216 0 _0491_
rlabel metal3 54096 41272 54096 41272 0 _0492_
rlabel metal3 53928 41720 53928 41720 0 _0493_
rlabel metal3 25032 45752 25032 45752 0 _0494_
rlabel metal2 53816 42280 53816 42280 0 _0495_
rlabel metal2 55776 42728 55776 42728 0 _0496_
rlabel metal2 54992 42840 54992 42840 0 _0497_
rlabel metal2 54096 42728 54096 42728 0 _0498_
rlabel metal2 53368 42448 53368 42448 0 _0499_
rlabel metal2 51912 48216 51912 48216 0 _0500_
rlabel metal3 53256 47432 53256 47432 0 _0501_
rlabel metal2 51688 48160 51688 48160 0 _0502_
rlabel metal2 52248 47824 52248 47824 0 _0503_
rlabel metal2 52584 48720 52584 48720 0 _0504_
rlabel metal3 25480 45920 25480 45920 0 _0505_
rlabel metal2 52584 50120 52584 50120 0 _0506_
rlabel metal2 52584 49224 52584 49224 0 _0507_
rlabel metal3 52864 48888 52864 48888 0 _0508_
rlabel metal2 52024 52696 52024 52696 0 _0509_
rlabel metal2 51128 56560 51128 56560 0 _0510_
rlabel metal3 49168 56840 49168 56840 0 _0511_
rlabel metal2 46536 56392 46536 56392 0 _0512_
rlabel metal3 47320 56056 47320 56056 0 _0513_
rlabel metal2 47320 55552 47320 55552 0 _0514_
rlabel metal2 47432 54992 47432 54992 0 _0515_
rlabel metal3 25368 46648 25368 46648 0 _0516_
rlabel metal2 40376 55832 40376 55832 0 _0517_
rlabel metal3 40656 56616 40656 56616 0 _0518_
rlabel metal2 44520 58072 44520 58072 0 _0519_
rlabel metal2 40040 58688 40040 58688 0 _0520_
rlabel metal2 40544 57848 40544 57848 0 _0521_
rlabel metal2 40096 56840 40096 56840 0 _0522_
rlabel metal2 40712 57176 40712 57176 0 _0523_
rlabel metal2 39760 56056 39760 56056 0 _0524_
rlabel metal3 41832 55832 41832 55832 0 _0525_
rlabel metal2 40040 56224 40040 56224 0 _0526_
rlabel metal3 25200 44520 25200 44520 0 _0527_
rlabel metal2 19320 58520 19320 58520 0 _0528_
rlabel metal3 13720 59192 13720 59192 0 _0529_
rlabel metal2 14784 59192 14784 59192 0 _0530_
rlabel metal2 13832 56504 13832 56504 0 _0531_
rlabel metal3 11760 56056 11760 56056 0 _0532_
rlabel metal2 13720 53760 13720 53760 0 _0533_
rlabel metal3 22456 48440 22456 48440 0 _0534_
rlabel metal2 11928 54880 11928 54880 0 _0535_
rlabel metal2 14280 56840 14280 56840 0 _0536_
rlabel metal2 14616 59024 14616 59024 0 _0537_
rlabel metal2 24584 44744 24584 44744 0 _0538_
rlabel metal2 15960 59584 15960 59584 0 _0539_
rlabel metal2 15456 58968 15456 58968 0 _0540_
rlabel metal3 17360 59080 17360 59080 0 _0541_
rlabel metal2 26936 59584 26936 59584 0 _0542_
rlabel metal2 26936 58520 26936 58520 0 _0543_
rlabel metal2 26824 58800 26824 58800 0 _0544_
rlabel metal2 28392 58408 28392 58408 0 _0545_
rlabel metal3 29960 57624 29960 57624 0 _0546_
rlabel metal2 31304 58072 31304 58072 0 _0547_
rlabel metal2 32088 58296 32088 58296 0 _0548_
rlabel metal2 25032 44632 25032 44632 0 _0549_
rlabel metal2 31080 56728 31080 56728 0 _0550_
rlabel metal2 32816 57624 32816 57624 0 _0551_
rlabel metal2 31752 57176 31752 57176 0 _0552_
rlabel metal2 31416 56560 31416 56560 0 _0553_
rlabel metal2 38696 56952 38696 56952 0 _0554_
rlabel metal2 27944 59584 27944 59584 0 _0555_
rlabel metal2 23016 59528 23016 59528 0 _0556_
rlabel metal2 33936 57848 33936 57848 0 _0557_
rlabel metal2 33768 59696 33768 59696 0 _0558_
rlabel metal2 24920 59472 24920 59472 0 _0559_
rlabel metal3 22176 6664 22176 6664 0 _0560_
rlabel metal2 13496 56336 13496 56336 0 _0561_
rlabel metal3 16800 56840 16800 56840 0 _0562_
rlabel metal2 15008 53704 15008 53704 0 _0563_
rlabel metal3 16632 53984 16632 53984 0 _0564_
rlabel metal2 16632 54992 16632 54992 0 _0565_
rlabel metal3 16912 56728 16912 56728 0 _0566_
rlabel metal2 16688 56952 16688 56952 0 _0567_
rlabel metal3 16912 58408 16912 58408 0 _0568_
rlabel metal2 20440 58128 20440 58128 0 _0569_
rlabel metal3 19152 58408 19152 58408 0 _0570_
rlabel metal2 21560 40656 21560 40656 0 _0571_
rlabel metal2 22120 58576 22120 58576 0 _0572_
rlabel metal2 22008 58912 22008 58912 0 _0573_
rlabel metal3 17136 57064 17136 57064 0 _0574_
rlabel metal2 17864 56560 17864 56560 0 _0575_
rlabel metal3 20216 56728 20216 56728 0 _0576_
rlabel metal3 23408 57064 23408 57064 0 _0577_
rlabel metal2 24472 56056 24472 56056 0 _0578_
rlabel metal3 24472 56840 24472 56840 0 _0579_
rlabel metal2 21784 58968 21784 58968 0 _0580_
rlabel metal2 23184 58296 23184 58296 0 _0581_
rlabel metal2 2296 33824 2296 33824 0 _0582_
rlabel metal2 23576 57624 23576 57624 0 _0583_
rlabel metal2 22680 56728 22680 56728 0 _0584_
rlabel metal2 22344 56280 22344 56280 0 _0585_
rlabel metal3 24024 12824 24024 12824 0 _0586_
rlabel metal2 22568 56336 22568 56336 0 _0587_
rlabel metal2 38248 56336 38248 56336 0 _0588_
rlabel metal2 23352 55496 23352 55496 0 _0589_
rlabel metal3 23464 56280 23464 56280 0 _0590_
rlabel metal2 38584 55720 38584 55720 0 _0591_
rlabel metal3 2016 42840 2016 42840 0 _0592_
rlabel metal2 24584 4928 24584 4928 0 _0593_
rlabel metal2 28112 4424 28112 4424 0 _0594_
rlabel metal2 21672 3864 21672 3864 0 _0595_
rlabel metal3 24108 3528 24108 3528 0 _0596_
rlabel metal2 26656 6664 26656 6664 0 _0597_
rlabel metal2 31864 4536 31864 4536 0 _0598_
rlabel metal2 32424 4536 32424 4536 0 _0599_
rlabel metal3 33096 3640 33096 3640 0 _0600_
rlabel metal2 26376 5320 26376 5320 0 _0601_
rlabel metal2 19544 42448 19544 42448 0 _0602_
rlabel metal2 29848 7560 29848 7560 0 _0603_
rlabel metal3 30800 7336 30800 7336 0 _0604_
rlabel metal2 32256 7336 32256 7336 0 _0605_
rlabel metal3 31920 6104 31920 6104 0 _0606_
rlabel metal2 32816 6776 32816 6776 0 _0607_
rlabel metal3 33208 5880 33208 5880 0 _0608_
rlabel metal2 29792 8456 29792 8456 0 _0609_
rlabel metal2 31528 10192 31528 10192 0 _0610_
rlabel metal2 32088 6664 32088 6664 0 _0611_
rlabel metal2 22792 36960 22792 36960 0 _0612_
rlabel metal3 31808 9800 31808 9800 0 _0613_
rlabel metal2 32760 9352 32760 9352 0 _0614_
rlabel metal2 25032 10248 25032 10248 0 _0615_
rlabel metal2 29008 11928 29008 11928 0 _0616_
rlabel metal2 29232 12152 29232 12152 0 _0617_
rlabel metal3 30520 12320 30520 12320 0 _0618_
rlabel metal2 31752 9912 31752 9912 0 _0619_
rlabel metal2 32088 10472 32088 10472 0 _0620_
rlabel metal2 31472 10808 31472 10808 0 _0621_
rlabel metal3 12712 23352 12712 23352 0 _0622_
rlabel metal2 30632 11536 30632 11536 0 _0623_
rlabel metal2 25928 11200 25928 11200 0 _0624_
rlabel metal2 26208 11256 26208 11256 0 _0625_
rlabel metal2 26488 13720 26488 13720 0 _0626_
rlabel metal3 30464 12824 30464 12824 0 _0627_
rlabel metal2 26432 14280 26432 14280 0 _0628_
rlabel metal2 27552 12936 27552 12936 0 _0629_
rlabel metal2 26376 10192 26376 10192 0 _0630_
rlabel metal2 5768 24976 5768 24976 0 _0631_
rlabel metal2 27720 16296 27720 16296 0 _0632_
rlabel metal2 27496 16464 27496 16464 0 _0633_
rlabel metal3 26376 16856 26376 16856 0 _0634_
rlabel metal3 26600 13048 26600 13048 0 _0635_
rlabel metal2 27160 14616 27160 14616 0 _0636_
rlabel metal2 26488 14616 26488 14616 0 _0637_
rlabel metal2 25144 14812 25144 14812 0 _0638_
rlabel metal2 26824 14700 26824 14700 0 _0639_
rlabel metal2 26488 19264 26488 19264 0 _0640_
rlabel metal3 3584 26488 3584 26488 0 _0641_
rlabel metal3 27720 17080 27720 17080 0 _0642_
rlabel metal3 26152 18648 26152 18648 0 _0643_
rlabel metal3 24136 18536 24136 18536 0 _0644_
rlabel metal2 28392 5544 28392 5544 0 _0645_
rlabel metal2 26264 5040 26264 5040 0 _0646_
rlabel metal2 26040 4760 26040 4760 0 _0647_
rlabel metal2 24808 18480 24808 18480 0 _0648_
rlabel metal3 26992 18424 26992 18424 0 _0649_
rlabel metal2 25592 4592 25592 4592 0 _0650_
rlabel metal2 2184 43512 2184 43512 0 _0651_
rlabel metal2 24808 5880 24808 5880 0 _0652_
rlabel metal2 26264 8064 26264 8064 0 _0653_
rlabel metal3 25256 6664 25256 6664 0 _0654_
rlabel metal2 23184 4536 23184 4536 0 _0655_
rlabel metal2 24696 5208 24696 5208 0 _0656_
rlabel metal2 22008 5096 22008 5096 0 _0657_
rlabel metal2 26712 7952 26712 7952 0 _0658_
rlabel metal2 26208 7448 26208 7448 0 _0659_
rlabel metal3 20944 37464 20944 37464 0 _0660_
rlabel metal2 25704 7784 25704 7784 0 _0661_
rlabel metal3 25256 7560 25256 7560 0 _0662_
rlabel metal2 24472 6272 24472 6272 0 _0663_
rlabel metal2 23856 5880 23856 5880 0 _0664_
rlabel metal2 24248 7840 24248 7840 0 _0665_
rlabel metal2 20664 7392 20664 7392 0 _0666_
rlabel metal3 23072 8792 23072 8792 0 _0667_
rlabel metal2 21112 7924 21112 7924 0 _0668_
rlabel metal2 22232 7504 22232 7504 0 _0669_
rlabel metal2 22008 42448 22008 42448 0 _0670_
rlabel metal2 22064 7672 22064 7672 0 _0671_
rlabel metal3 23184 10584 23184 10584 0 _0672_
rlabel metal3 23688 10472 23688 10472 0 _0673_
rlabel metal2 22120 10752 22120 10752 0 _0674_
rlabel metal2 22904 8372 22904 8372 0 _0675_
rlabel metal2 22960 7784 22960 7784 0 _0676_
rlabel via2 22008 10472 22008 10472 0 _0677_
rlabel metal3 20272 10584 20272 10584 0 _0678_
rlabel metal3 24192 37240 24192 37240 0 _0679_
rlabel metal2 24584 11592 24584 11592 0 _0680_
rlabel metal2 23688 12656 23688 12656 0 _0681_
rlabel metal2 22792 10584 22792 10584 0 _0682_
rlabel metal2 22344 12208 22344 12208 0 _0683_
rlabel metal2 21784 12488 21784 12488 0 _0684_
rlabel metal2 22848 14392 22848 14392 0 _0685_
rlabel metal3 24304 14392 24304 14392 0 _0686_
rlabel metal2 22232 15456 22232 15456 0 _0687_
rlabel metal2 22792 13048 22792 13048 0 _0688_
rlabel metal3 5712 26376 5712 26376 0 _0689_
rlabel metal2 23240 12376 23240 12376 0 _0690_
rlabel metal3 21840 15960 21840 15960 0 _0691_
rlabel metal2 21840 14504 21840 14504 0 _0692_
rlabel metal2 23016 17640 23016 17640 0 _0693_
rlabel metal2 22792 15288 22792 15288 0 _0694_
rlabel metal2 21896 17360 21896 17360 0 _0695_
rlabel metal3 21672 16968 21672 16968 0 _0696_
rlabel metal3 22736 19208 22736 19208 0 _0697_
rlabel metal2 14448 25368 14448 25368 0 _0698_
rlabel metal2 22176 17640 22176 17640 0 _0699_
rlabel metal2 22568 18312 22568 18312 0 _0700_
rlabel metal2 10248 14560 10248 14560 0 _0701_
rlabel metal3 10024 10696 10024 10696 0 _0702_
rlabel metal2 4312 12432 4312 12432 0 _0703_
rlabel metal3 5768 11368 5768 11368 0 _0704_
rlabel metal2 3920 12936 3920 12936 0 _0705_
rlabel metal2 5768 12208 5768 12208 0 _0706_
rlabel metal2 19712 41048 19712 41048 0 _0707_
rlabel metal2 4312 10192 4312 10192 0 _0708_
rlabel metal2 5040 10472 5040 10472 0 _0709_
rlabel metal3 5376 9688 5376 9688 0 _0710_
rlabel metal2 5488 3528 5488 3528 0 _0711_
rlabel metal2 6720 3640 6720 3640 0 _0712_
rlabel metal3 5544 5208 5544 5208 0 _0713_
rlabel metal2 5880 6384 5880 6384 0 _0714_
rlabel metal2 18816 24024 18816 24024 0 _0715_
rlabel metal2 8120 7840 8120 7840 0 _0716_
rlabel metal3 9408 8680 9408 8680 0 _0717_
rlabel metal2 7560 21224 7560 21224 0 _0718_
rlabel metal3 5824 20328 5824 20328 0 _0719_
rlabel metal2 8232 21896 8232 21896 0 _0720_
rlabel metal3 6832 21672 6832 21672 0 _0721_
rlabel metal2 19768 41272 19768 41272 0 _0722_
rlabel metal2 12824 22624 12824 22624 0 _0723_
rlabel metal2 13384 21560 13384 21560 0 _0724_
rlabel metal3 13608 20552 13608 20552 0 _0725_
rlabel metal3 12320 19992 12320 19992 0 _0726_
rlabel metal2 12936 21280 12936 21280 0 _0727_
rlabel metal3 12040 20776 12040 20776 0 _0728_
rlabel metal2 9968 19208 9968 19208 0 _0729_
rlabel metal2 19376 43400 19376 43400 0 _0730_
rlabel metal3 10080 20888 10080 20888 0 _0731_
rlabel metal2 6216 20384 6216 20384 0 _0732_
rlabel metal2 11704 21000 11704 21000 0 _0733_
rlabel metal2 15176 21112 15176 21112 0 _0734_
rlabel metal2 17304 22792 17304 22792 0 _0735_
rlabel metal2 16464 20776 16464 20776 0 _0736_
rlabel metal2 18760 22120 18760 22120 0 _0737_
rlabel metal2 19656 43120 19656 43120 0 _0738_
rlabel metal3 17360 21672 17360 21672 0 _0739_
rlabel metal2 19488 21560 19488 21560 0 _0740_
rlabel metal2 21784 4480 21784 4480 0 _0741_
rlabel metal2 17416 35000 17416 35000 0 _0742_
rlabel metal2 18760 43456 18760 43456 0 _0743_
rlabel metal2 19488 42168 19488 42168 0 _0744_
rlabel metal4 15176 32200 15176 32200 0 _0745_
rlabel metal2 25760 39704 25760 39704 0 _0746_
rlabel metal2 30744 37744 30744 37744 0 _0747_
rlabel metal3 31080 38696 31080 38696 0 _0748_
rlabel metal2 39144 43344 39144 43344 0 _0749_
rlabel metal3 19600 48328 19600 48328 0 _0750_
rlabel metal3 16296 42616 16296 42616 0 _0751_
rlabel metal2 21896 42000 21896 42000 0 _0752_
rlabel metal2 18872 40936 18872 40936 0 _0753_
rlabel metal2 11256 25032 11256 25032 0 _0754_
rlabel metal3 21672 40600 21672 40600 0 _0755_
rlabel metal3 23352 41944 23352 41944 0 _0756_
rlabel metal3 9632 23240 9632 23240 0 _0757_
rlabel metal2 20888 44016 20888 44016 0 _0758_
rlabel metal2 10696 43120 10696 43120 0 _0759_
rlabel metal2 20440 43624 20440 43624 0 _0760_
rlabel metal3 3248 20328 3248 20328 0 _0761_
rlabel metal2 16184 40432 16184 40432 0 _0762_
rlabel metal2 2744 41384 2744 41384 0 _0763_
rlabel metal2 2912 37800 2912 37800 0 _0764_
rlabel metal3 20608 44296 20608 44296 0 _0765_
rlabel metal2 19432 43848 19432 43848 0 _0766_
rlabel metal2 24136 42616 24136 42616 0 _0767_
rlabel metal2 26712 41832 26712 41832 0 _0768_
rlabel metal2 26544 41048 26544 41048 0 _0769_
rlabel metal2 26600 47600 26600 47600 0 _0770_
rlabel metal3 28616 43736 28616 43736 0 _0771_
rlabel metal2 28840 45304 28840 45304 0 _0772_
rlabel metal2 2856 48608 2856 48608 0 _0773_
rlabel metal2 5320 21784 5320 21784 0 _0774_
rlabel metal3 18928 40600 18928 40600 0 _0775_
rlabel metal2 3024 41384 3024 41384 0 _0776_
rlabel metal2 3976 41440 3976 41440 0 _0777_
rlabel metal2 18200 32032 18200 32032 0 _0778_
rlabel metal3 19880 50344 19880 50344 0 _0779_
rlabel metal3 10864 24696 10864 24696 0 _0780_
rlabel metal2 3640 42448 3640 42448 0 _0781_
rlabel metal2 25368 57792 25368 57792 0 _0782_
rlabel metal3 2688 24024 2688 24024 0 _0783_
rlabel metal2 7560 47880 7560 47880 0 _0784_
rlabel metal2 5824 49224 5824 49224 0 _0785_
rlabel metal2 5880 48496 5880 48496 0 _0786_
rlabel metal3 4592 25256 4592 25256 0 _0787_
rlabel metal3 5152 46872 5152 46872 0 _0788_
rlabel metal2 2296 55104 2296 55104 0 _0789_
rlabel metal2 5376 45304 5376 45304 0 _0790_
rlabel metal2 25816 44520 25816 44520 0 _0791_
rlabel metal2 29624 40544 29624 40544 0 _0792_
rlabel metal2 30184 41832 30184 41832 0 _0793_
rlabel metal3 37968 49112 37968 49112 0 _0794_
rlabel metal2 14840 36736 14840 36736 0 _0795_
rlabel metal2 16072 34048 16072 34048 0 _0796_
rlabel metal3 17248 32424 17248 32424 0 _0797_
rlabel metal2 14616 38080 14616 38080 0 _0798_
rlabel metal2 24416 37464 24416 37464 0 _0799_
rlabel metal2 2072 26768 2072 26768 0 _0800_
rlabel metal2 13944 42784 13944 42784 0 _0801_
rlabel metal2 2184 40656 2184 40656 0 _0802_
rlabel metal3 13832 38136 13832 38136 0 _0803_
rlabel metal3 8120 23576 8120 23576 0 _0804_
rlabel metal2 14840 33768 14840 33768 0 _0805_
rlabel metal2 1848 36624 1848 36624 0 _0806_
rlabel metal2 2520 33376 2520 33376 0 _0807_
rlabel metal2 14392 37856 14392 37856 0 _0808_
rlabel metal2 23576 37688 23576 37688 0 _0809_
rlabel metal3 29400 36456 29400 36456 0 _0810_
rlabel metal2 28840 35952 28840 35952 0 _0811_
rlabel metal2 25256 46256 25256 46256 0 _0812_
rlabel metal2 30520 45528 30520 45528 0 _0813_
rlabel metal2 31472 55440 31472 55440 0 _0814_
rlabel metal2 32088 45192 32088 45192 0 _0815_
rlabel metal2 30072 44800 30072 44800 0 _0816_
rlabel metal2 31752 45696 31752 45696 0 _0817_
rlabel metal2 28616 45360 28616 45360 0 _0818_
rlabel metal2 26824 45472 26824 45472 0 _0819_
rlabel metal3 7952 49112 7952 49112 0 _0820_
rlabel metal2 15736 43400 15736 43400 0 _0821_
rlabel metal3 7392 50344 7392 50344 0 _0822_
rlabel metal3 9520 50008 9520 50008 0 _0823_
rlabel metal3 18648 45192 18648 45192 0 _0824_
rlabel metal2 10976 51352 10976 51352 0 _0825_
rlabel metal2 10528 48216 10528 48216 0 _0826_
rlabel metal2 1904 37464 1904 37464 0 _0827_
rlabel metal4 17864 45640 17864 45640 0 _0828_
rlabel metal3 11200 50008 11200 50008 0 _0829_
rlabel metal2 11704 51408 11704 51408 0 _0830_
rlabel metal2 11368 51464 11368 51464 0 _0831_
rlabel metal2 10696 48216 10696 48216 0 _0832_
rlabel metal3 9632 50680 9632 50680 0 _0833_
rlabel metal3 9912 51352 9912 51352 0 _0834_
rlabel metal2 22960 39704 22960 39704 0 _0835_
rlabel metal2 26768 20888 26768 20888 0 _0836_
rlabel metal3 12096 25480 12096 25480 0 _0837_
rlabel metal2 11872 24136 11872 24136 0 _0838_
rlabel metal2 11536 24696 11536 24696 0 _0839_
rlabel metal2 11928 25088 11928 25088 0 _0840_
rlabel metal2 6552 46816 6552 46816 0 _0841_
rlabel metal2 7448 39816 7448 39816 0 _0842_
rlabel metal3 11592 25312 11592 25312 0 _0843_
rlabel metal2 10584 25984 10584 25984 0 _0844_
rlabel metal2 10024 24920 10024 24920 0 _0845_
rlabel metal3 10920 25256 10920 25256 0 _0846_
rlabel metal2 18648 25872 18648 25872 0 _0847_
rlabel metal3 21504 23464 21504 23464 0 _0848_
rlabel metal2 3080 53312 3080 53312 0 _0849_
rlabel metal3 19488 38696 19488 38696 0 _0850_
rlabel metal2 20664 39928 20664 39928 0 _0851_
rlabel metal2 16744 24920 16744 24920 0 _0852_
rlabel metal3 19992 29288 19992 29288 0 _0853_
rlabel metal2 20216 45416 20216 45416 0 _0854_
rlabel metal2 20552 45584 20552 45584 0 _0855_
rlabel metal3 18648 29400 18648 29400 0 _0856_
rlabel metal2 19264 34328 19264 34328 0 _0857_
rlabel metal2 22232 22512 22232 22512 0 _0858_
rlabel metal2 21112 35112 21112 35112 0 _0859_
rlabel metal2 21784 35952 21784 35952 0 _0860_
rlabel metal2 21112 35616 21112 35616 0 _0861_
rlabel metal2 22120 20552 22120 20552 0 _0862_
rlabel metal2 22680 20328 22680 20328 0 _0863_
rlabel metal3 24556 21336 24556 21336 0 _0864_
rlabel metal2 29848 19152 29848 19152 0 _0865_
rlabel metal3 8176 36568 8176 36568 0 _0866_
rlabel metal2 10752 22456 10752 22456 0 _0867_
rlabel metal2 6608 39368 6608 39368 0 _0868_
rlabel metal2 5768 38192 5768 38192 0 _0869_
rlabel metal2 7448 37688 7448 37688 0 _0870_
rlabel metal3 10584 20496 10584 20496 0 _0871_
rlabel metal3 17304 32312 17304 32312 0 _0872_
rlabel metal2 2072 36792 2072 36792 0 _0873_
rlabel metal2 10136 32088 10136 32088 0 _0874_
rlabel metal2 18536 32200 18536 32200 0 _0875_
rlabel metal2 10136 28560 10136 28560 0 _0876_
rlabel metal2 20048 29960 20048 29960 0 _0877_
rlabel metal2 22456 29736 22456 29736 0 _0878_
rlabel metal3 30240 28504 30240 28504 0 _0879_
rlabel metal2 30240 28616 30240 28616 0 _0880_
rlabel metal2 29512 22960 29512 22960 0 _0881_
rlabel metal2 50904 49504 50904 49504 0 _0882_
rlabel metal2 29736 16352 29736 16352 0 _0883_
rlabel metal2 41272 28840 41272 28840 0 _0884_
rlabel metal2 30968 13440 30968 13440 0 _0885_
rlabel metal3 21280 41720 21280 41720 0 _0886_
rlabel metal2 22456 32592 22456 32592 0 _0887_
rlabel metal2 25928 31248 25928 31248 0 _0888_
rlabel metal2 18536 46032 18536 46032 0 _0889_
rlabel metal3 16968 35952 16968 35952 0 _0890_
rlabel metal3 18704 35672 18704 35672 0 _0891_
rlabel metal2 17416 36848 17416 36848 0 _0892_
rlabel metal2 8792 42896 8792 42896 0 _0893_
rlabel metal2 2968 45920 2968 45920 0 _0894_
rlabel metal2 18088 36176 18088 36176 0 _0895_
rlabel metal2 13048 26208 13048 26208 0 _0896_
rlabel metal3 22568 31864 22568 31864 0 _0897_
rlabel metal2 27608 30520 27608 30520 0 _0898_
rlabel metal2 27832 30576 27832 30576 0 _0899_
rlabel metal2 29512 18816 29512 18816 0 _0900_
rlabel metal3 31360 15512 31360 15512 0 _0901_
rlabel metal2 16856 39312 16856 39312 0 _0902_
rlabel metal2 18872 34272 18872 34272 0 _0903_
rlabel metal3 18144 33320 18144 33320 0 _0904_
rlabel metal2 24360 32872 24360 32872 0 _0905_
rlabel metal2 14392 31528 14392 31528 0 _0906_
rlabel metal3 17360 32648 17360 32648 0 _0907_
rlabel metal2 19096 34104 19096 34104 0 _0908_
rlabel metal3 20552 33096 20552 33096 0 _0909_
rlabel metal3 22288 32312 22288 32312 0 _0910_
rlabel metal2 28000 18984 28000 18984 0 _0911_
rlabel metal2 26600 28392 26600 28392 0 _0912_
rlabel metal2 32536 20832 32536 20832 0 _0913_
rlabel metal2 30520 15568 30520 15568 0 _0914_
rlabel metal2 2072 30128 2072 30128 0 _0915_
rlabel metal2 12264 43960 12264 43960 0 _0916_
rlabel metal3 15008 23352 15008 23352 0 _0917_
rlabel metal2 15960 43568 15960 43568 0 _0918_
rlabel metal3 16744 44072 16744 44072 0 _0919_
rlabel metal2 15400 35896 15400 35896 0 _0920_
rlabel metal3 18648 38808 18648 38808 0 _0921_
rlabel metal2 20216 41720 20216 41720 0 _0922_
rlabel metal2 19992 38304 19992 38304 0 _0923_
rlabel metal2 21672 37688 21672 37688 0 _0924_
rlabel metal4 26376 19320 26376 19320 0 _0925_
rlabel metal2 34216 19488 34216 19488 0 _0926_
rlabel metal2 30128 15064 30128 15064 0 _0927_
rlabel metal2 30800 15512 30800 15512 0 _0928_
rlabel metal2 31304 16464 31304 16464 0 _0929_
rlabel metal2 30128 17080 30128 17080 0 _0930_
rlabel metal2 29344 18312 29344 18312 0 _0931_
rlabel metal2 8960 40600 8960 40600 0 _0932_
rlabel metal2 10696 38864 10696 38864 0 _0933_
rlabel metal2 1960 46032 1960 46032 0 _0934_
rlabel metal2 10864 38920 10864 38920 0 _0935_
rlabel metal3 19656 26768 19656 26768 0 _0936_
rlabel metal2 2744 40096 2744 40096 0 _0937_
rlabel metal3 18536 40488 18536 40488 0 _0938_
rlabel metal2 21336 39256 21336 39256 0 _0939_
rlabel metal2 24472 34552 24472 34552 0 _0940_
rlabel metal2 28168 33264 28168 33264 0 _0941_
rlabel metal2 29960 32144 29960 32144 0 _0942_
rlabel metal2 26152 40208 26152 40208 0 _0943_
rlabel metal3 28952 20776 28952 20776 0 _0944_
rlabel metal2 29848 25200 29848 25200 0 _0945_
rlabel metal3 31920 53088 31920 53088 0 _0946_
rlabel metal2 28224 19880 28224 19880 0 _0947_
rlabel metal2 26936 20664 26936 20664 0 _0948_
rlabel metal2 26544 20888 26544 20888 0 _0949_
rlabel metal2 27720 44800 27720 44800 0 _0950_
rlabel metal3 26992 44296 26992 44296 0 _0951_
rlabel metal2 27384 45528 27384 45528 0 _0952_
rlabel metal2 26040 46200 26040 46200 0 _0953_
rlabel metal2 25704 46480 25704 46480 0 _0954_
rlabel metal2 13832 22736 13832 22736 0 _0955_
rlabel metal3 16072 50008 16072 50008 0 _0956_
rlabel metal2 15848 50064 15848 50064 0 _0957_
rlabel metal2 15568 51352 15568 51352 0 _0958_
rlabel metal2 14056 51296 14056 51296 0 _0959_
rlabel metal2 15960 51744 15960 51744 0 _0960_
rlabel metal2 15736 51856 15736 51856 0 _0961_
rlabel metal2 28056 50624 28056 50624 0 _0962_
rlabel metal2 14336 50008 14336 50008 0 _0963_
rlabel metal2 13944 50960 13944 50960 0 _0964_
rlabel metal2 53816 48356 53816 48356 0 _0965_
rlabel metal4 24248 53480 24248 53480 0 _0966_
rlabel metal2 18200 51352 18200 51352 0 _0967_
rlabel metal3 19376 51240 19376 51240 0 _0968_
rlabel metal2 19376 51464 19376 51464 0 _0969_
rlabel metal3 23800 51912 23800 51912 0 _0970_
rlabel metal2 18424 52472 18424 52472 0 _0971_
rlabel metal2 28280 54768 28280 54768 0 _0972_
rlabel metal2 23352 52528 23352 52528 0 _0973_
rlabel metal2 24360 52696 24360 52696 0 _0974_
rlabel metal2 23576 52248 23576 52248 0 _0975_
rlabel metal2 15288 39592 15288 39592 0 _0976_
rlabel metal2 7784 39760 7784 39760 0 _0977_
rlabel metal2 14952 39984 14952 39984 0 _0978_
rlabel metal3 3360 23352 3360 23352 0 _0979_
rlabel metal2 10808 35896 10808 35896 0 _0980_
rlabel metal3 9744 36456 9744 36456 0 _0981_
rlabel metal2 6216 36624 6216 36624 0 _0982_
rlabel metal2 14504 39592 14504 39592 0 _0983_
rlabel metal3 19320 39088 19320 39088 0 _0984_
rlabel metal2 42168 40040 42168 40040 0 _0985_
rlabel metal3 13440 27160 13440 27160 0 _0986_
rlabel metal2 15904 20888 15904 20888 0 _0987_
rlabel metal2 3192 44856 3192 44856 0 _0988_
rlabel metal2 17752 36456 17752 36456 0 _0989_
rlabel metal3 19600 39368 19600 39368 0 _0990_
rlabel metal2 15176 55412 15176 55412 0 _0991_
rlabel metal4 18872 39816 18872 39816 0 _0992_
rlabel metal3 17640 39032 17640 39032 0 _0993_
rlabel metal2 19432 39648 19432 39648 0 _0994_
rlabel metal3 21672 39704 21672 39704 0 _0995_
rlabel metal2 45304 41776 45304 41776 0 _0996_
rlabel metal2 24920 49840 24920 49840 0 _0997_
rlabel metal3 11648 41832 11648 41832 0 _0998_
rlabel metal2 14168 42056 14168 42056 0 _0999_
rlabel metal3 14168 40600 14168 40600 0 _1000_
rlabel metal2 14840 41664 14840 41664 0 _1001_
rlabel metal2 21672 42392 21672 42392 0 _1002_
rlabel metal2 22120 43512 22120 43512 0 _1003_
rlabel metal3 16352 42840 16352 42840 0 _1004_
rlabel metal2 18760 42784 18760 42784 0 _1005_
rlabel metal2 22456 42616 22456 42616 0 _1006_
rlabel metal2 46760 39648 46760 39648 0 _1007_
rlabel metal2 2632 38472 2632 38472 0 _1008_
rlabel metal3 2744 38696 2744 38696 0 _1009_
rlabel metal2 4200 36736 4200 36736 0 _1010_
rlabel metal3 4928 35000 4928 35000 0 _1011_
rlabel metal3 5264 35672 5264 35672 0 _1012_
rlabel metal2 4872 36680 4872 36680 0 _1013_
rlabel metal2 3416 35896 3416 35896 0 _1014_
rlabel metal2 3528 36344 3528 36344 0 _1015_
rlabel metal3 13440 22568 13440 22568 0 _1016_
rlabel metal2 47208 25088 47208 25088 0 _1017_
rlabel metal2 3136 38808 3136 38808 0 _1018_
rlabel metal3 4872 38808 4872 38808 0 _1019_
rlabel metal2 6888 36064 6888 36064 0 _1020_
rlabel metal2 8512 40376 8512 40376 0 _1021_
rlabel metal3 8568 38248 8568 38248 0 _1022_
rlabel metal3 7728 38360 7728 38360 0 _1023_
rlabel metal3 12488 15064 12488 15064 0 _1024_
rlabel metal2 40040 40432 40040 40432 0 _1025_
rlabel metal2 2296 47264 2296 47264 0 _1026_
rlabel metal2 3192 46928 3192 46928 0 _1027_
rlabel metal2 8792 46928 8792 46928 0 _1028_
rlabel metal2 10136 48496 10136 48496 0 _1029_
rlabel metal2 9744 47656 9744 47656 0 _1030_
rlabel metal2 9968 43736 9968 43736 0 _1031_
rlabel metal3 9912 47320 9912 47320 0 _1032_
rlabel metal2 9016 47208 9016 47208 0 _1033_
rlabel metal2 18648 45640 18648 45640 0 _1034_
rlabel metal4 26824 18984 26824 18984 0 _1035_
rlabel metal3 7448 45080 7448 45080 0 _1036_
rlabel metal3 11088 29288 11088 29288 0 _1037_
rlabel metal2 10696 28560 10696 28560 0 _1038_
rlabel metal2 11032 28728 11032 28728 0 _1039_
rlabel metal2 11368 29904 11368 29904 0 _1040_
rlabel metal2 15400 31472 15400 31472 0 _1041_
rlabel metal3 16184 30296 16184 30296 0 _1042_
rlabel metal2 16856 30688 16856 30688 0 _1043_
rlabel metal3 19992 30184 19992 30184 0 _1044_
rlabel metal3 24360 23688 24360 23688 0 _1045_
rlabel metal2 7000 50736 7000 50736 0 _1046_
rlabel metal2 9128 46256 9128 46256 0 _1047_
rlabel metal3 12880 25480 12880 25480 0 _1048_
rlabel metal2 6776 46592 6776 46592 0 _1049_
rlabel metal3 7448 50680 7448 50680 0 _1050_
rlabel metal2 6888 45248 6888 45248 0 _1051_
rlabel metal2 6944 44520 6944 44520 0 _1052_
rlabel metal2 7728 45080 7728 45080 0 _1053_
rlabel metal2 7224 45864 7224 45864 0 _1054_
rlabel metal3 21896 50568 21896 50568 0 _1055_
rlabel metal3 42896 8232 42896 8232 0 _1056_
rlabel metal2 18032 29512 18032 29512 0 _1057_
rlabel metal3 18592 28840 18592 28840 0 _1058_
rlabel metal2 12600 28504 12600 28504 0 _1059_
rlabel metal3 14784 28728 14784 28728 0 _1060_
rlabel metal2 19096 28560 19096 28560 0 _1061_
rlabel metal2 17920 28392 17920 28392 0 _1062_
rlabel metal2 14056 26488 14056 26488 0 _1063_
rlabel metal2 19320 28224 19320 28224 0 _1064_
rlabel metal3 19208 25032 19208 25032 0 _1065_
rlabel metal2 19992 27664 19992 27664 0 _1066_
rlabel metal2 40712 34048 40712 34048 0 _1067_
rlabel metal2 16296 33376 16296 33376 0 _1068_
rlabel metal2 16464 32648 16464 32648 0 _1069_
rlabel metal2 16016 33432 16016 33432 0 _1070_
rlabel metal2 23464 32648 23464 32648 0 _1071_
rlabel metal2 23016 34496 23016 34496 0 _1072_
rlabel metal2 21560 32480 21560 32480 0 _1073_
rlabel metal2 20216 31976 20216 31976 0 _1074_
rlabel metal2 22792 33320 22792 33320 0 _1075_
rlabel metal2 23576 32144 23576 32144 0 _1076_
rlabel metal3 42252 26824 42252 26824 0 _1077_
rlabel metal2 42056 13832 42056 13832 0 _1078_
rlabel metal2 40544 12376 40544 12376 0 _1079_
rlabel metal2 14952 45192 14952 45192 0 _1080_
rlabel metal2 14728 46200 14728 46200 0 _1081_
rlabel metal3 18704 45752 18704 45752 0 _1082_
rlabel metal2 16968 47152 16968 47152 0 _1083_
rlabel metal2 18536 47040 18536 47040 0 _1084_
rlabel metal2 18256 45864 18256 45864 0 _1085_
rlabel metal2 19880 46144 19880 46144 0 _1086_
rlabel metal2 24976 20104 24976 20104 0 _1087_
rlabel metal2 24864 26600 24864 26600 0 _1088_
rlabel metal4 30632 22456 30632 22456 0 _1089_
rlabel metal2 5096 44072 5096 44072 0 _1090_
rlabel metal2 5320 43680 5320 43680 0 _1091_
rlabel metal3 7112 40600 7112 40600 0 _1092_
rlabel metal2 7000 41608 7000 41608 0 _1093_
rlabel metal2 5880 40320 5880 40320 0 _1094_
rlabel metal2 5600 40600 5600 40600 0 _1095_
rlabel metal2 23576 29232 23576 29232 0 _1096_
rlabel metal3 40376 21560 40376 21560 0 _1097_
rlabel metal2 30408 21952 30408 21952 0 _1098_
rlabel metal3 31528 21784 31528 21784 0 _1099_
rlabel metal2 30520 21392 30520 21392 0 _1100_
rlabel metal3 28392 26264 28392 26264 0 _1101_
rlabel metal3 28056 26152 28056 26152 0 _1102_
rlabel metal2 27496 26488 27496 26488 0 _1103_
rlabel metal2 26152 29008 26152 29008 0 _1104_
rlabel metal3 26712 29400 26712 29400 0 _1105_
rlabel metal2 25760 30072 25760 30072 0 _1106_
rlabel metal2 25256 31584 25256 31584 0 _1107_
rlabel metal3 25536 35896 25536 35896 0 _1108_
rlabel metal3 25816 40376 25816 40376 0 _1109_
rlabel metal2 25928 44856 25928 44856 0 _1110_
rlabel metal2 25032 52584 25032 52584 0 _1111_
rlabel metal2 25088 51352 25088 51352 0 _1112_
rlabel metal2 24528 50568 24528 50568 0 _1113_
rlabel metal2 24976 51128 24976 51128 0 _1114_
rlabel metal2 20552 20944 20552 20944 0 _1115_
rlabel metal2 25928 23128 25928 23128 0 _1116_
rlabel metal2 25592 26376 25592 26376 0 _1117_
rlabel metal3 18200 23912 18200 23912 0 _1118_
rlabel metal3 46200 38696 46200 38696 0 _1119_
rlabel metal2 52696 30576 52696 30576 0 _1120_
rlabel metal2 50568 25816 50568 25816 0 _1121_
rlabel metal3 24696 23240 24696 23240 0 _1122_
rlabel metal3 22736 23240 22736 23240 0 _1123_
rlabel metal2 20664 20720 20664 20720 0 _1124_
rlabel metal2 21672 21056 21672 21056 0 _1125_
rlabel metal2 46536 26096 46536 26096 0 _1126_
rlabel metal3 47880 27160 47880 27160 0 _1127_
rlabel metal2 52304 28616 52304 28616 0 _1128_
rlabel metal2 50456 26712 50456 26712 0 _1129_
rlabel metal2 23968 20216 23968 20216 0 _1130_
rlabel metal2 39816 21504 39816 21504 0 _1131_
rlabel metal2 44072 11424 44072 11424 0 _1132_
rlabel metal2 47544 29792 47544 29792 0 _1133_
rlabel metal3 49168 30296 49168 30296 0 _1134_
rlabel metal2 52136 29736 52136 29736 0 _1135_
rlabel metal2 54152 29736 54152 29736 0 _1136_
rlabel metal3 53088 28840 53088 28840 0 _1137_
rlabel metal2 53816 30744 53816 30744 0 _1138_
rlabel metal2 33432 38080 33432 38080 0 _1139_
rlabel metal2 20664 23520 20664 23520 0 _1140_
rlabel metal2 22736 40936 22736 40936 0 _1141_
rlabel metal2 32200 24416 32200 24416 0 _1142_
rlabel metal2 39144 32816 39144 32816 0 _1143_
rlabel metal2 18872 20944 18872 20944 0 _1144_
rlabel metal2 26264 30464 26264 30464 0 _1145_
rlabel metal2 39256 32144 39256 32144 0 _1146_
rlabel metal3 21504 23688 21504 23688 0 _1147_
rlabel metal2 21896 25648 21896 25648 0 _1148_
rlabel metal2 22120 25984 22120 25984 0 _1149_
rlabel metal2 23912 26544 23912 26544 0 _1150_
rlabel metal3 29008 50456 29008 50456 0 _1151_
rlabel metal3 42448 32536 42448 32536 0 _1152_
rlabel metal2 43624 30688 43624 30688 0 _1153_
rlabel metal2 34104 30968 34104 30968 0 _1154_
rlabel metal3 37072 19208 37072 19208 0 _1155_
rlabel metal2 36568 26208 36568 26208 0 _1156_
rlabel metal2 40376 29512 40376 29512 0 _1157_
rlabel metal2 32312 40992 32312 40992 0 _1158_
rlabel metal2 38696 23912 38696 23912 0 _1159_
rlabel metal2 36792 31640 36792 31640 0 _1160_
rlabel metal3 35168 30408 35168 30408 0 _1161_
rlabel metal2 41832 30576 41832 30576 0 _1162_
rlabel metal3 40600 33096 40600 33096 0 _1163_
rlabel metal3 26544 26488 26544 26488 0 _1164_
rlabel metal2 38808 36792 38808 36792 0 _1165_
rlabel metal2 39928 32816 39928 32816 0 _1166_
rlabel metal3 41496 30856 41496 30856 0 _1167_
rlabel metal2 42728 31752 42728 31752 0 _1168_
rlabel metal2 43176 31248 43176 31248 0 _1169_
rlabel metal2 51800 31304 51800 31304 0 _1170_
rlabel metal2 28056 53424 28056 53424 0 _1171_
rlabel metal2 51240 28728 51240 28728 0 _1172_
rlabel metal2 44184 45304 44184 45304 0 _1173_
rlabel metal3 48608 31080 48608 31080 0 _1174_
rlabel metal3 46704 24696 46704 24696 0 _1175_
rlabel metal2 38808 26152 38808 26152 0 _1176_
rlabel metal3 44688 23352 44688 23352 0 _1177_
rlabel metal2 49616 31080 49616 31080 0 _1178_
rlabel metal2 51072 30856 51072 30856 0 _1179_
rlabel metal2 52472 31416 52472 31416 0 _1180_
rlabel metal3 53368 31640 53368 31640 0 _1181_
rlabel metal3 53088 31192 53088 31192 0 _1182_
rlabel metal2 53928 31920 53928 31920 0 _1183_
rlabel metal2 36456 26096 36456 26096 0 _1184_
rlabel metal2 37800 29680 37800 29680 0 _1185_
rlabel metal2 23800 25088 23800 25088 0 _1186_
rlabel metal2 26152 26152 26152 26152 0 _1187_
rlabel metal2 22008 25536 22008 25536 0 _1188_
rlabel metal3 23856 26376 23856 26376 0 _1189_
rlabel metal3 31304 27048 31304 27048 0 _1190_
rlabel metal2 23352 21448 23352 21448 0 _1191_
rlabel metal2 24696 23968 24696 23968 0 _1192_
rlabel metal2 32312 22624 32312 22624 0 _1193_
rlabel metal2 25032 28168 25032 28168 0 _1194_
rlabel metal2 37576 28840 37576 28840 0 _1195_
rlabel metal2 43848 31864 43848 31864 0 _1196_
rlabel metal2 30968 18536 30968 18536 0 _1197_
rlabel metal2 30744 33544 30744 33544 0 _1198_
rlabel metal3 33040 34888 33040 34888 0 _1199_
rlabel metal2 31080 40236 31080 40236 0 _1200_
rlabel metal2 31528 33040 31528 33040 0 _1201_
rlabel metal2 32088 32312 32088 32312 0 _1202_
rlabel metal2 44408 33040 44408 33040 0 _1203_
rlabel metal3 45304 31640 45304 31640 0 _1204_
rlabel metal3 44856 31752 44856 31752 0 _1205_
rlabel metal2 45360 31752 45360 31752 0 _1206_
rlabel metal2 55272 31640 55272 31640 0 _1207_
rlabel metal2 31976 34384 31976 34384 0 _1208_
rlabel metal2 29960 34384 29960 34384 0 _1209_
rlabel metal2 45528 33656 45528 33656 0 _1210_
rlabel metal3 34328 35672 34328 35672 0 _1211_
rlabel metal2 35112 34720 35112 34720 0 _1212_
rlabel metal2 35000 26264 35000 26264 0 _1213_
rlabel metal2 37576 26488 37576 26488 0 _1214_
rlabel metal2 34216 34384 34216 34384 0 _1215_
rlabel metal2 45864 34664 45864 34664 0 _1216_
rlabel metal3 44744 35784 44744 35784 0 _1217_
rlabel metal2 46536 34384 46536 34384 0 _1218_
rlabel metal2 47432 34440 47432 34440 0 _1219_
rlabel metal3 41944 34216 41944 34216 0 _1220_
rlabel metal2 32088 34888 32088 34888 0 _1221_
rlabel metal2 41944 34328 41944 34328 0 _1222_
rlabel metal2 40824 35616 40824 35616 0 _1223_
rlabel metal2 30968 49728 30968 49728 0 _1224_
rlabel metal2 41832 36064 41832 36064 0 _1225_
rlabel metal2 41664 35112 41664 35112 0 _1226_
rlabel metal3 46088 33992 46088 33992 0 _1227_
rlabel via2 54824 31864 54824 31864 0 _1228_
rlabel metal2 56168 33320 56168 33320 0 _1229_
rlabel metal2 54488 33040 54488 33040 0 _1230_
rlabel metal2 55888 31864 55888 31864 0 _1231_
rlabel metal2 56728 34608 56728 34608 0 _1232_
rlabel metal2 46760 34104 46760 34104 0 _1233_
rlabel metal2 53256 35448 53256 35448 0 _1234_
rlabel metal2 46536 36064 46536 36064 0 _1235_
rlabel metal3 42784 36568 42784 36568 0 _1236_
rlabel metal2 40376 17136 40376 17136 0 _1237_
rlabel metal3 35392 34888 35392 34888 0 _1238_
rlabel metal2 42728 36120 42728 36120 0 _1239_
rlabel metal2 39816 36792 39816 36792 0 _1240_
rlabel metal2 26040 48048 26040 48048 0 _1241_
rlabel metal2 39928 37296 39928 37296 0 _1242_
rlabel metal3 41664 37128 41664 37128 0 _1243_
rlabel metal3 43792 37128 43792 37128 0 _1244_
rlabel metal2 46872 37520 46872 37520 0 _1245_
rlabel metal3 35000 25368 35000 25368 0 _1246_
rlabel metal3 35336 39592 35336 39592 0 _1247_
rlabel metal2 39032 20440 39032 20440 0 _1248_
rlabel metal3 34384 39032 34384 39032 0 _1249_
rlabel metal2 35784 37464 35784 37464 0 _1250_
rlabel metal2 24864 22904 24864 22904 0 _1251_
rlabel metal2 32984 21168 32984 21168 0 _1252_
rlabel metal3 33152 31752 33152 31752 0 _1253_
rlabel metal2 35224 38668 35224 38668 0 _1254_
rlabel metal2 46312 37240 46312 37240 0 _1255_
rlabel metal2 53704 34888 53704 34888 0 _1256_
rlabel metal2 54824 36008 54824 36008 0 _1257_
rlabel metal2 50008 32256 50008 32256 0 _1258_
rlabel metal2 53816 34832 53816 34832 0 _1259_
rlabel metal3 42336 34888 42336 34888 0 _1260_
rlabel metal2 43456 34888 43456 34888 0 _1261_
rlabel metal2 51240 34608 51240 34608 0 _1262_
rlabel metal3 53032 44184 53032 44184 0 _1263_
rlabel metal2 53816 19936 53816 19936 0 _1264_
rlabel metal2 51352 29344 51352 29344 0 _1265_
rlabel metal2 49112 33880 49112 33880 0 _1266_
rlabel metal2 48776 12600 48776 12600 0 _1267_
rlabel metal2 50120 40880 50120 40880 0 _1268_
rlabel metal2 50792 35728 50792 35728 0 _1269_
rlabel metal2 51800 35280 51800 35280 0 _1270_
rlabel metal3 53088 34888 53088 34888 0 _1271_
rlabel metal2 54712 35280 54712 35280 0 _1272_
rlabel metal2 56448 35448 56448 35448 0 _1273_
rlabel metal2 57512 36176 57512 36176 0 _1274_
rlabel metal3 57344 35672 57344 35672 0 _1275_
rlabel metal2 57960 37576 57960 37576 0 _1276_
rlabel metal2 52360 35392 52360 35392 0 _1277_
rlabel metal2 53760 37912 53760 37912 0 _1278_
rlabel metal2 54096 34328 54096 34328 0 _1279_
rlabel metal2 54600 38920 54600 38920 0 _1280_
rlabel metal2 49616 34216 49616 34216 0 _1281_
rlabel metal2 49784 36120 49784 36120 0 _1282_
rlabel metal2 49896 38864 49896 38864 0 _1283_
rlabel metal2 44016 36680 44016 36680 0 _1284_
rlabel metal2 43288 36736 43288 36736 0 _1285_
rlabel metal2 51800 37968 51800 37968 0 _1286_
rlabel metal2 50176 41384 50176 41384 0 _1287_
rlabel metal2 44408 44744 44408 44744 0 _1288_
rlabel metal2 40488 11592 40488 11592 0 _1289_
rlabel metal2 50008 41608 50008 41608 0 _1290_
rlabel metal2 47320 41664 47320 41664 0 _1291_
rlabel metal3 49896 41944 49896 41944 0 _1292_
rlabel metal2 51912 38640 51912 38640 0 _1293_
rlabel metal2 50456 39088 50456 39088 0 _1294_
rlabel metal3 50960 38808 50960 38808 0 _1295_
rlabel metal2 46536 37184 46536 37184 0 _1296_
rlabel metal2 47096 37128 47096 37128 0 _1297_
rlabel metal3 47432 38808 47432 38808 0 _1298_
rlabel metal2 40152 38724 40152 38724 0 _1299_
rlabel metal2 33880 25424 33880 25424 0 _1300_
rlabel metal2 34048 36568 34048 36568 0 _1301_
rlabel metal3 36288 38024 36288 38024 0 _1302_
rlabel metal2 39592 25144 39592 25144 0 _1303_
rlabel metal2 25704 50204 25704 50204 0 _1304_
rlabel metal3 27832 52920 27832 52920 0 _1305_
rlabel metal2 37520 34888 37520 34888 0 _1306_
rlabel metal2 38360 38668 38360 38668 0 _1307_
rlabel metal2 40320 38696 40320 38696 0 _1308_
rlabel metal2 44408 39592 44408 39592 0 _1309_
rlabel metal2 34216 42336 34216 42336 0 _1310_
rlabel metal2 35560 39480 35560 39480 0 _1311_
rlabel metal2 36008 39088 36008 39088 0 _1312_
rlabel metal2 43736 40656 43736 40656 0 _1313_
rlabel metal2 34552 44352 34552 44352 0 _1314_
rlabel metal2 35672 41608 35672 41608 0 _1315_
rlabel metal2 37912 41832 37912 41832 0 _1316_
rlabel metal2 27944 51464 27944 51464 0 _1317_
rlabel metal2 28392 52640 28392 52640 0 _1318_
rlabel metal2 37688 40768 37688 40768 0 _1319_
rlabel metal2 44632 40656 44632 40656 0 _1320_
rlabel metal2 43848 39984 43848 39984 0 _1321_
rlabel metal2 48216 40096 48216 40096 0 _1322_
rlabel metal2 16072 19824 16072 19824 0 _1323_
rlabel metal2 50008 39088 50008 39088 0 _1324_
rlabel metal2 53592 39200 53592 39200 0 _1325_
rlabel metal3 57008 38696 57008 38696 0 _1326_
rlabel metal2 56784 48104 56784 48104 0 _1327_
rlabel metal2 51576 38808 51576 38808 0 _1328_
rlabel metal2 52024 44968 52024 44968 0 _1329_
rlabel metal3 49672 40488 49672 40488 0 _1330_
rlabel metal2 50344 39984 50344 39984 0 _1331_
rlabel metal2 51352 45080 51352 45080 0 _1332_
rlabel metal2 48776 42392 48776 42392 0 _1333_
rlabel metal2 3080 28224 3080 28224 0 _1334_
rlabel metal2 49784 46312 49784 46312 0 _1335_
rlabel metal2 38696 37464 38696 37464 0 _1336_
rlabel metal2 39032 37520 39032 37520 0 _1337_
rlabel metal2 47152 46536 47152 46536 0 _1338_
rlabel metal3 47432 45080 47432 45080 0 _1339_
rlabel metal2 46200 44352 46200 44352 0 _1340_
rlabel metal2 45416 42952 45416 42952 0 _1341_
rlabel metal3 45080 44408 45080 44408 0 _1342_
rlabel metal2 46648 44632 46648 44632 0 _1343_
rlabel metal2 47992 46424 47992 46424 0 _1344_
rlabel metal2 7000 23296 7000 23296 0 _1345_
rlabel metal2 48776 46312 48776 46312 0 _1346_
rlabel metal3 49336 45080 49336 45080 0 _1347_
rlabel metal2 43960 41664 43960 41664 0 _1348_
rlabel metal2 44576 41384 44576 41384 0 _1349_
rlabel metal2 48440 44184 48440 44184 0 _1350_
rlabel metal2 43960 43568 43960 43568 0 _1351_
rlabel metal2 39256 34328 39256 34328 0 _1352_
rlabel metal2 43736 42896 43736 42896 0 _1353_
rlabel metal2 42784 44296 42784 44296 0 _1354_
rlabel metal2 39816 44688 39816 44688 0 _1355_
rlabel metal2 18760 24864 18760 24864 0 _1356_
rlabel metal2 34888 44576 34888 44576 0 _1357_
rlabel metal3 35448 45080 35448 45080 0 _1358_
rlabel metal3 37464 45192 37464 45192 0 _1359_
rlabel metal2 37912 44016 37912 44016 0 _1360_
rlabel metal3 39368 44408 39368 44408 0 _1361_
rlabel metal2 41384 44632 41384 44632 0 _1362_
rlabel metal3 40656 44296 40656 44296 0 _1363_
rlabel metal3 42112 44296 42112 44296 0 _1364_
rlabel metal2 48328 44296 48328 44296 0 _1365_
rlabel via2 49112 44968 49112 44968 0 _1366_
rlabel metal3 24136 41272 24136 41272 0 _1367_
rlabel metal3 50848 44968 50848 44968 0 _1368_
rlabel metal2 52136 44688 52136 44688 0 _1369_
rlabel metal3 53368 45864 53368 45864 0 _1370_
rlabel metal2 54152 38696 54152 38696 0 _1371_
rlabel metal2 53592 38080 53592 38080 0 _1372_
rlabel metal3 54600 45640 54600 45640 0 _1373_
rlabel metal2 54488 46872 54488 46872 0 _1374_
rlabel metal2 55384 48440 55384 48440 0 _1375_
rlabel metal2 58128 45864 58128 45864 0 _1376_
rlabel metal3 47208 26824 47208 26824 0 _1377_
rlabel metal2 24360 44968 24360 44968 0 _1378_
rlabel metal2 43960 11144 43960 11144 0 _1379_
rlabel metal3 46032 26488 46032 26488 0 _1380_
rlabel metal2 50680 27552 50680 27552 0 _1381_
rlabel metal3 50120 27160 50120 27160 0 _1382_
rlabel metal3 52136 27720 52136 27720 0 _1383_
rlabel metal2 55048 27888 55048 27888 0 _1384_
rlabel metal2 32200 25536 32200 25536 0 _1385_
rlabel metal3 33600 25592 33600 25592 0 _1386_
rlabel metal2 34216 25872 34216 25872 0 _1387_
rlabel via2 42056 30072 42056 30072 0 _1388_
rlabel metal2 14224 25592 14224 25592 0 _1389_
rlabel metal3 39648 30856 39648 30856 0 _1390_
rlabel metal2 39816 31248 39816 31248 0 _1391_
rlabel metal2 39872 29400 39872 29400 0 _1392_
rlabel metal3 41104 29400 41104 29400 0 _1393_
rlabel metal2 39144 27496 39144 27496 0 _1394_
rlabel metal2 40712 29120 40712 29120 0 _1395_
rlabel metal2 55160 29176 55160 29176 0 _1396_
rlabel metal3 54992 29288 54992 29288 0 _1397_
rlabel metal2 58072 29288 58072 29288 0 _1398_
rlabel metal3 56784 29512 56784 29512 0 _1399_
rlabel metal2 15904 40936 15904 40936 0 _1400_
rlabel metal2 57848 30772 57848 30772 0 _1401_
rlabel metal3 33040 18312 33040 18312 0 _1402_
rlabel metal2 24584 26992 24584 26992 0 _1403_
rlabel metal2 34776 24472 34776 24472 0 _1404_
rlabel metal2 35560 26096 35560 26096 0 _1405_
rlabel metal2 35896 25032 35896 25032 0 _1406_
rlabel metal2 34944 25368 34944 25368 0 _1407_
rlabel metal3 35392 23240 35392 23240 0 _1408_
rlabel metal2 43512 29456 43512 29456 0 _1409_
rlabel metal2 41608 28840 41608 28840 0 _1410_
rlabel metal2 7672 3920 7672 3920 0 _1411_
rlabel metal3 42840 28504 42840 28504 0 _1412_
rlabel metal2 44072 28448 44072 28448 0 _1413_
rlabel metal2 43512 28896 43512 28896 0 _1414_
rlabel metal2 56728 29120 56728 29120 0 _1415_
rlabel metal2 56840 30800 56840 30800 0 _1416_
rlabel metal2 58072 28616 58072 28616 0 _1417_
rlabel metal2 57456 28504 57456 28504 0 _1418_
rlabel metal2 58296 29680 58296 29680 0 _1419_
rlabel metal2 57624 30240 57624 30240 0 _1420_
rlabel metal3 57400 32536 57400 32536 0 _1421_
rlabel metal2 2744 24248 2744 24248 0 _1422_
rlabel metal2 58128 33320 58128 33320 0 _1423_
rlabel metal2 57512 33040 57512 33040 0 _1424_
rlabel metal2 57736 36736 57736 36736 0 _1425_
rlabel metal2 57848 37744 57848 37744 0 _1426_
rlabel metal2 58408 40712 58408 40712 0 _1427_
rlabel metal2 57568 37464 57568 37464 0 _1428_
rlabel metal2 57848 46312 57848 46312 0 _1429_
rlabel metal2 55272 48160 55272 48160 0 _1430_
rlabel metal2 55944 51016 55944 51016 0 _1431_
rlabel metal2 44240 10584 44240 10584 0 _1432_
rlabel metal2 5992 26208 5992 26208 0 _1433_
rlabel metal2 39256 26040 39256 26040 0 _1434_
rlabel metal3 40488 13944 40488 13944 0 _1435_
rlabel metal3 41160 26152 41160 26152 0 _1436_
rlabel metal2 35112 28280 35112 28280 0 _1437_
rlabel metal2 40712 25760 40712 25760 0 _1438_
rlabel metal3 40096 27048 40096 27048 0 _1439_
rlabel metal2 41048 26600 41048 26600 0 _1440_
rlabel metal3 41944 25592 41944 25592 0 _1441_
rlabel metal2 52136 26768 52136 26768 0 _1442_
rlabel metal2 53480 26544 53480 26544 0 _1443_
rlabel metal2 7112 31360 7112 31360 0 _1444_
rlabel metal2 46368 24472 46368 24472 0 _1445_
rlabel metal2 46872 24752 46872 24752 0 _1446_
rlabel metal3 48272 24920 48272 24920 0 _1447_
rlabel metal2 50232 24192 50232 24192 0 _1448_
rlabel metal2 48440 25144 48440 25144 0 _1449_
rlabel metal2 50120 25144 50120 25144 0 _1450_
rlabel metal3 52360 25480 52360 25480 0 _1451_
rlabel metal2 54376 25816 54376 25816 0 _1452_
rlabel metal2 54488 26712 54488 26712 0 _1453_
rlabel metal2 56504 26656 56504 26656 0 _1454_
rlabel metal3 2296 36456 2296 36456 0 _1455_
rlabel metal2 38024 23800 38024 23800 0 _1456_
rlabel metal2 28504 23968 28504 23968 0 _1457_
rlabel metal2 38808 21952 38808 21952 0 _1458_
rlabel metal2 36232 23632 36232 23632 0 _1459_
rlabel metal3 37520 23800 37520 23800 0 _1460_
rlabel metal3 37688 23688 37688 23688 0 _1461_
rlabel metal2 42056 23520 42056 23520 0 _1462_
rlabel metal3 40320 24136 40320 24136 0 _1463_
rlabel metal3 43064 23128 43064 23128 0 _1464_
rlabel metal3 43400 25480 43400 25480 0 _1465_
rlabel metal3 3024 30184 3024 30184 0 _1466_
rlabel metal2 43176 24752 43176 24752 0 _1467_
rlabel metal3 42000 23800 42000 23800 0 _1468_
rlabel metal3 44408 23912 44408 23912 0 _1469_
rlabel metal2 45528 24696 45528 24696 0 _1470_
rlabel metal2 52696 23464 52696 23464 0 _1471_
rlabel metal2 53368 23912 53368 23912 0 _1472_
rlabel metal2 52808 25032 52808 25032 0 _1473_
rlabel metal2 57960 25480 57960 25480 0 _1474_
rlabel metal2 57176 26264 57176 26264 0 _1475_
rlabel metal2 56952 25872 56952 25872 0 _1476_
rlabel metal2 6888 21952 6888 21952 0 _1477_
rlabel metal3 56896 24920 56896 24920 0 _1478_
rlabel metal2 56616 27776 56616 27776 0 _1479_
rlabel metal2 57344 39592 57344 39592 0 _1480_
rlabel metal3 57400 41160 57400 41160 0 _1481_
rlabel metal2 57568 40600 57568 40600 0 _1482_
rlabel metal2 56448 45192 56448 45192 0 _1483_
rlabel metal3 57064 43736 57064 43736 0 _1484_
rlabel metal2 56168 46312 56168 46312 0 _1485_
rlabel metal2 56392 42000 56392 42000 0 _1486_
rlabel metal2 42056 21056 42056 21056 0 _1487_
rlabel metal2 6496 25480 6496 25480 0 _1488_
rlabel metal2 38976 12264 38976 12264 0 _1489_
rlabel metal3 44352 21448 44352 21448 0 _1490_
rlabel metal2 45976 21840 45976 21840 0 _1491_
rlabel metal2 43960 23240 43960 23240 0 _1492_
rlabel metal2 44856 23800 44856 23800 0 _1493_
rlabel metal2 45752 22288 45752 22288 0 _1494_
rlabel metal3 46928 22120 46928 22120 0 _1495_
rlabel metal3 45192 22344 45192 22344 0 _1496_
rlabel metal2 51128 22792 51128 22792 0 _1497_
rlabel metal2 51016 22736 51016 22736 0 _1498_
rlabel metal3 1960 38136 1960 38136 0 _1499_
rlabel metal2 54040 22792 54040 22792 0 _1500_
rlabel metal2 51240 21504 51240 21504 0 _1501_
rlabel metal2 36344 27328 36344 27328 0 _1502_
rlabel metal2 36232 28224 36232 28224 0 _1503_
rlabel via1 39144 21000 39144 21000 0 _1504_
rlabel metal2 35784 19544 35784 19544 0 _1505_
rlabel metal3 33544 20776 33544 20776 0 _1506_
rlabel metal2 35784 20888 35784 20888 0 _1507_
rlabel metal2 38136 20832 38136 20832 0 _1508_
rlabel metal3 37128 20776 37128 20776 0 _1509_
rlabel metal3 12432 26488 12432 26488 0 _1510_
rlabel metal2 46536 20496 46536 20496 0 _1511_
rlabel metal2 46760 22792 46760 22792 0 _1512_
rlabel metal3 47152 21784 47152 21784 0 _1513_
rlabel metal2 47208 21336 47208 21336 0 _1514_
rlabel metal2 47880 21504 47880 21504 0 _1515_
rlabel metal3 48608 21560 48608 21560 0 _1516_
rlabel metal2 52136 21392 52136 21392 0 _1517_
rlabel metal3 51464 21672 51464 21672 0 _1518_
rlabel metal2 51744 21784 51744 21784 0 _1519_
rlabel metal2 53592 22400 53592 22400 0 _1520_
rlabel metal2 2632 31192 2632 31192 0 _1521_
rlabel metal3 53984 23016 53984 23016 0 _1522_
rlabel metal2 54712 22624 54712 22624 0 _1523_
rlabel metal2 54152 22848 54152 22848 0 _1524_
rlabel metal2 55160 24304 55160 24304 0 _1525_
rlabel metal2 57288 23128 57288 23128 0 _1526_
rlabel metal2 55832 28000 55832 28000 0 _1527_
rlabel metal2 55552 24472 55552 24472 0 _1528_
rlabel metal2 56280 39984 56280 39984 0 _1529_
rlabel metal2 55944 44772 55944 44772 0 _1530_
rlabel metal2 55384 49672 55384 49672 0 _1531_
rlabel metal2 2464 35000 2464 35000 0 _1532_
rlabel metal3 54824 55944 54824 55944 0 _1533_
rlabel metal2 43904 7336 43904 7336 0 _1534_
rlabel metal3 44240 7672 44240 7672 0 _1535_
rlabel metal3 41608 14952 41608 14952 0 _1536_
rlabel metal2 42840 16576 42840 16576 0 _1537_
rlabel metal3 43400 17640 43400 17640 0 _1538_
rlabel metal3 33544 19768 33544 19768 0 _1539_
rlabel metal2 42616 19600 42616 19600 0 _1540_
rlabel metal2 42280 19600 42280 19600 0 _1541_
rlabel metal2 42504 20216 42504 20216 0 _1542_
rlabel metal2 7448 25032 7448 25032 0 _1543_
rlabel metal2 42952 19600 42952 19600 0 _1544_
rlabel metal2 43512 18872 43512 18872 0 _1545_
rlabel metal2 44296 18424 44296 18424 0 _1546_
rlabel metal3 45864 18424 45864 18424 0 _1547_
rlabel metal2 47824 18424 47824 18424 0 _1548_
rlabel metal2 52136 18144 52136 18144 0 _1549_
rlabel metal3 49392 17752 49392 17752 0 _1550_
rlabel metal2 50176 17864 50176 17864 0 _1551_
rlabel metal3 33264 21672 33264 21672 0 _1552_
rlabel metal2 32872 21616 32872 21616 0 _1553_
rlabel metal3 1848 26488 1848 26488 0 _1554_
rlabel metal2 38808 19376 38808 19376 0 _1555_
rlabel metal2 36400 15624 36400 15624 0 _1556_
rlabel metal3 35280 17640 35280 17640 0 _1557_
rlabel metal3 36960 17416 36960 17416 0 _1558_
rlabel metal3 37184 17864 37184 17864 0 _1559_
rlabel metal2 39144 18088 39144 18088 0 _1560_
rlabel metal2 38024 18144 38024 18144 0 _1561_
rlabel metal2 45640 18480 45640 18480 0 _1562_
rlabel metal3 37184 20104 37184 20104 0 _1563_
rlabel metal2 37464 20720 37464 20720 0 _1564_
rlabel metal2 16632 44520 16632 44520 0 _1565_
rlabel metal3 42784 19432 42784 19432 0 _1566_
rlabel metal2 46536 18704 46536 18704 0 _1567_
rlabel metal3 45584 17752 45584 17752 0 _1568_
rlabel metal2 46872 19264 46872 19264 0 _1569_
rlabel metal3 48328 19096 48328 19096 0 _1570_
rlabel metal3 48888 19208 48888 19208 0 _1571_
rlabel metal2 50736 18984 50736 18984 0 _1572_
rlabel metal2 49672 19208 49672 19208 0 _1573_
rlabel metal2 51464 18312 51464 18312 0 _1574_
rlabel metal2 51352 18424 51352 18424 0 _1575_
rlabel metal2 9800 28112 9800 28112 0 _1576_
rlabel metal2 52136 17640 52136 17640 0 _1577_
rlabel metal2 51688 18704 51688 18704 0 _1578_
rlabel metal2 53480 18424 53480 18424 0 _1579_
rlabel metal2 55384 21896 55384 21896 0 _1580_
rlabel metal3 55832 19208 55832 19208 0 _1581_
rlabel metal2 55048 20888 55048 20888 0 _1582_
rlabel metal3 57232 20104 57232 20104 0 _1583_
rlabel metal3 56952 18536 56952 18536 0 _1584_
rlabel metal2 57456 21560 57456 21560 0 _1585_
rlabel metal3 57064 20664 57064 20664 0 _1586_
rlabel metal2 3808 26488 3808 26488 0 _1587_
rlabel metal3 57120 21448 57120 21448 0 _1588_
rlabel metal2 43736 16352 43736 16352 0 _1589_
rlabel metal2 39704 12824 39704 12824 0 _1590_
rlabel metal2 40768 15400 40768 15400 0 _1591_
rlabel metal2 42952 15792 42952 15792 0 _1592_
rlabel metal2 43624 13216 43624 13216 0 _1593_
rlabel metal2 44296 14448 44296 14448 0 _1594_
rlabel metal2 48664 15680 48664 15680 0 _1595_
rlabel metal2 46368 16184 46368 16184 0 _1596_
rlabel metal2 46872 14812 46872 14812 0 _1597_
rlabel metal2 2800 49000 2800 49000 0 _1598_
rlabel metal2 4312 2422 4312 2422 0 clk
rlabel metal2 7336 14952 7336 14952 0 clknet_0_clk
rlabel metal2 5656 5096 5656 5096 0 clknet_2_0__leaf_clk
rlabel metal2 15064 7448 15064 7448 0 clknet_2_1__leaf_clk
rlabel metal2 5096 17752 5096 17752 0 clknet_2_2__leaf_clk
rlabel metal3 15624 10584 15624 10584 0 clknet_2_3__leaf_clk
rlabel metal2 9016 12040 9016 12040 0 csTable.address\[0\]
rlabel metal2 8960 9240 8960 9240 0 csTable.address\[1\]
rlabel metal3 9464 4312 9464 4312 0 csTable.address\[2\]
rlabel metal2 6664 5600 6664 5600 0 csTable.address\[3\]
rlabel metal2 8344 7336 8344 7336 0 csTable.address\[4\]
rlabel metal3 7672 20776 7672 20776 0 csTable.address\[5\]
rlabel metal2 8960 22120 8960 22120 0 csTable.address\[6\]
rlabel metal2 13048 21644 13048 21644 0 csTable.address\[7\]
rlabel metal3 28840 3416 28840 3416 0 divSel[0]
rlabel metal2 38808 2086 38808 2086 0 divSel[1]
rlabel metal2 48104 3136 48104 3136 0 divSel[2]
rlabel metal2 55888 3416 55888 3416 0 divSel[3]
rlabel metal3 21784 4312 21784 4312 0 freeRunCntr\[0\]
rlabel metal2 26040 8288 26040 8288 0 freeRunCntr\[10\]
rlabel metal3 23632 8232 23632 8232 0 freeRunCntr\[11\]
rlabel metal2 23576 10304 23576 10304 0 freeRunCntr\[12\]
rlabel metal2 23576 12488 23576 12488 0 freeRunCntr\[13\]
rlabel metal2 23520 13944 23520 13944 0 freeRunCntr\[14\]
rlabel metal2 19096 14924 19096 14924 0 freeRunCntr\[15\]
rlabel metal2 12992 8344 12992 8344 0 freeRunCntr\[16\]
rlabel metal3 4816 12152 4816 12152 0 freeRunCntr\[17\]
rlabel metal2 20216 5600 20216 5600 0 freeRunCntr\[1\]
rlabel metal2 13272 17360 13272 17360 0 freeRunCntr\[26\]
rlabel metal2 10528 21672 10528 21672 0 freeRunCntr\[27\]
rlabel metal3 9184 20776 9184 20776 0 freeRunCntr\[28\]
rlabel metal3 51800 40936 51800 40936 0 freeRunCntr\[2\]
rlabel metal2 50456 48104 50456 48104 0 freeRunCntr\[3\]
rlabel metal2 51464 49224 51464 49224 0 freeRunCntr\[4\]
rlabel metal2 24304 12712 24304 12712 0 freeRunCntr\[5\]
rlabel metal2 24248 13888 24248 13888 0 freeRunCntr\[6\]
rlabel metal2 23968 14616 23968 14616 0 freeRunCntr\[7\]
rlabel metal2 24136 4704 24136 4704 0 freeRunCntr\[8\]
rlabel metal2 20888 5376 20888 5376 0 freeRunCntr\[9\]
rlabel metal2 26376 3864 26376 3864 0 net1
rlabel metal2 12208 17080 12208 17080 0 net10
rlabel metal2 7784 15736 7784 15736 0 net11
rlabel metal2 20216 6384 20216 6384 0 net12
rlabel metal2 26432 6664 26432 6664 0 net2
rlabel metal2 26824 7280 26824 7280 0 net3
rlabel metal3 45584 3304 45584 3304 0 net4
rlabel metal2 15624 3640 15624 3640 0 net5
rlabel metal2 50456 59864 50456 59864 0 net6
rlabel metal2 11032 59696 11032 59696 0 net7
rlabel metal2 30408 59864 30408 59864 0 net8
rlabel metal2 8344 6384 8344 6384 0 net9
rlabel metal2 50232 61642 50232 61642 0 qcomplex
rlabel metal2 10136 62678 10136 62678 0 qcos
rlabel metal3 30632 60088 30632 60088 0 qsin
rlabel metal2 12936 2086 12936 2086 0 rst
rlabel metal3 11256 16912 11256 16912 0 sigRom.address\[0\]
rlabel metal2 17080 19264 17080 19264 0 sigRom.address\[1\]
rlabel metal2 19096 17080 19096 17080 0 sigRom.address\[2\]
rlabel metal2 19096 19544 19096 19544 0 sigRom.address\[3\]
<< properties >>
string FIXED_BBOX 0 0 60397 63981
<< end >>
