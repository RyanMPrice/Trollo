VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO WavePWM
  CLASS BLOCK ;
  FOREIGN WavePWM ;
  ORIGIN 0.000 0.000 ;
  SIZE 301.985 BY 319.905 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 21.280 0.000 21.840 4.000 ;
    END
  END clk
  PIN divSel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 150.640 0.000 151.200 4.000 ;
    END
  END divSel[0]
  PIN divSel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 193.760 0.000 194.320 4.000 ;
    END
  END divSel[1]
  PIN divSel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 236.880 0.000 237.440 4.000 ;
    END
  END divSel[2]
  PIN divSel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 280.000 0.000 280.560 4.000 ;
    END
  END divSel[3]
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 107.520 0.000 108.080 4.000 ;
    END
  END enable
  PIN qcomplex
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 250.880 315.905 251.440 319.905 ;
    END
  END qcomplex
  PIN qcos
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 315.905 50.960 319.905 ;
    END
  END qcos
  PIN qsin
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 150.640 315.905 151.200 319.905 ;
    END
  END qsin
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 64.400 0.000 64.960 4.000 ;
    END
  END rst
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 302.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 302.140 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 302.140 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 302.140 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 14.710 295.120 302.140 ;
      LAYER Metal2 ;
        RECT 4.620 315.605 50.100 315.905 ;
        RECT 51.260 315.605 150.340 315.905 ;
        RECT 151.500 315.605 250.580 315.905 ;
        RECT 251.740 315.605 293.860 315.905 ;
        RECT 4.620 4.300 293.860 315.605 ;
        RECT 4.620 4.000 20.980 4.300 ;
        RECT 22.140 4.000 64.100 4.300 ;
        RECT 65.260 4.000 107.220 4.300 ;
        RECT 108.380 4.000 150.340 4.300 ;
        RECT 151.500 4.000 193.460 4.300 ;
        RECT 194.620 4.000 236.580 4.300 ;
        RECT 237.740 4.000 279.700 4.300 ;
        RECT 280.860 4.000 293.860 4.300 ;
      LAYER Metal3 ;
        RECT 4.570 15.540 293.910 304.500 ;
      LAYER Metal4 ;
        RECT 10.780 302.440 288.820 304.550 ;
        RECT 10.780 37.610 21.940 302.440 ;
        RECT 24.140 37.610 98.740 302.440 ;
        RECT 100.940 37.610 175.540 302.440 ;
        RECT 177.740 37.610 252.340 302.440 ;
        RECT 254.540 37.610 288.820 302.440 ;
  END
END WavePWM
END LIBRARY

