magic
tech gf180mcuC
magscale 1 5
timestamp 1670260637
<< obsm1 >>
rect 672 1538 4392 3166
<< metal2 >>
rect 1232 4600 1288 5000
rect 3696 4600 3752 5000
rect 840 0 896 400
rect 2464 0 2520 400
rect 4088 0 4144 400
<< obsm2 >>
rect 854 4570 1202 4600
rect 1318 4570 3666 4600
rect 3782 4570 4378 4600
rect 854 430 4378 4570
rect 926 400 2434 430
rect 2550 400 4058 430
rect 4174 400 4378 430
<< metal3 >>
rect 0 3696 400 3752
rect 0 1232 400 1288
<< obsm3 >>
rect 430 3666 4383 3738
rect 400 1318 4383 3666
rect 430 1246 4383 1318
<< metal4 >>
rect 1047 1538 1207 3166
rect 1502 1538 1662 3166
rect 1957 1538 2117 3166
rect 2412 1538 2572 3166
rect 2867 1538 3027 3166
rect 3322 1538 3482 3166
rect 3777 1538 3937 3166
rect 4232 1538 4392 3166
<< labels >>
rlabel metal2 s 2464 0 2520 400 6 INmb
port 1 nsew signal input
rlabel metal2 s 840 0 896 400 6 INpb
port 2 nsew signal input
rlabel metal3 s 0 3696 400 3752 6 cmnmos
port 3 nsew signal output
rlabel metal3 s 0 1232 400 1288 6 cmpmos
port 4 nsew signal output
rlabel metal2 s 4088 0 4144 400 6 oe
port 5 nsew signal input
rlabel metal2 s 3696 4600 3752 5000 6 onmos
port 6 nsew signal output
rlabel metal2 s 1232 4600 1288 5000 6 opmos
port 7 nsew signal output
rlabel metal4 s 1047 1538 1207 3166 6 vdd
port 8 nsew power bidirectional
rlabel metal4 s 1957 1538 2117 3166 6 vdd
port 8 nsew power bidirectional
rlabel metal4 s 2867 1538 3027 3166 6 vdd
port 8 nsew power bidirectional
rlabel metal4 s 3777 1538 3937 3166 6 vdd
port 8 nsew power bidirectional
rlabel metal4 s 1502 1538 1662 3166 6 vss
port 9 nsew ground bidirectional
rlabel metal4 s 2412 1538 2572 3166 6 vss
port 9 nsew ground bidirectional
rlabel metal4 s 3322 1538 3482 3166 6 vss
port 9 nsew ground bidirectional
rlabel metal4 s 4232 1538 4392 3166 6 vss
port 9 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 5000 5000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 75984
string GDS_FILE /mnt/c/Users/rmprice/Documents/Github/Trollo/openlane/user_Digota/runs/22_12_05_10_15/results/signoff/DIGOTA.magic.gds
string GDS_START 39552
<< end >>

