* NGSPICE file created from WavePWM.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_4 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_4 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_4 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_4 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

.subckt WavePWM clk divSel[0] divSel[1] divSel[2] divSel[3] enable qcomplex qcos qsin
+ rst vdd vss
XTAP_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3155_ _0706_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3086_ _0634_ _0637_ _0642_ _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2106_ _0941_ _0942_ _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2037_ _1085_ _0757_ _0854_ _0855_ _0889_ _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_35_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2939_ _0479_ _0484_ _0487_ _0946_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_10_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2954__A1 freeRunCntr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1757__A2 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2706__A1 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1693__A1 _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3198__A1 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1748__A2 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2945__A1 freeRunCntr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2103__I _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2173__A2 _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1987__A2 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3189__A1 _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2936__A1 _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1739__A2 _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2724_ _1120_ _0231_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2655_ _0149_ _0150_ _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1606_ _1389_ _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_2586_ _0080_ _0097_ _0099_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__3113__A1 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3207_ _0029_ net10 clknet_2_2__leaf_clk freeRunCntr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_67_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3138_ _0692_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1801__B _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3069_ _0624_ _0593_ _0625_ _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_27_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1978__A2 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1902__A2 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3104__A1 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1666__A1 freeRunCntr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1666__B2 freeRunCntr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1969__A2 _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2091__A1 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2440_ _0913_ _1248_ _1252_ _0926_ _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_2371_ _1340_ _1427_ _1428_ _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2854__B1 _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2082__A1 _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2707_ _0229_ _0232_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2385__A2 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2790__C1 _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2638_ _0154_ _0156_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2688__A3 _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2569_ _0073_ _0075_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1648__A1 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2073__A1 _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1820__A1 _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2376__A2 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2128__A2 _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1639__A1 _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2064__A1 freeRunCntr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1940_ _0787_ _0806_ _0988_ _0783_ _0602_ _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1811__A1 _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1871_ _0873_ _0874_ _0920_ _0762_ _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2423_ _1290_ _1481_ _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2354_ _1185_ _1195_ _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2285_ _1172_ _1268_ _1333_ _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_37_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2055__A1 freeRunCntr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1802__A1 _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2046__A1 _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2597__A2 _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2349__A2 _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3216__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2070_ sigRom.address\[3\] _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__2285__A1 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2972_ _0518_ _0522_ _0523_ _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1923_ _0955_ _0971_ _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_1854_ _0873_ _0874_ _0890_ _0857_ _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1785_ _0750_ _0823_ _0825_ _0831_ _0834_ _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XANTENNA__3117__I freeRunCntr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2406_ _1462_ _1463_ _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2337_ _1390_ _1391_ _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2268_ _1314_ _1315_ _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2177__B _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2199_ _1139_ _1246_ _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2028__A1 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1787__B1 _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2019__A1 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3171_ _0719_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2122_ _1153_ _1168_ _1169_ _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_47_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2053_ _0882_ _1067_ _1045_ freeRunCntr\[6\] _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2258__A1 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2258__B2 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2955_ _0480_ _0346_ _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2886_ _0397_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1906_ _1323_ _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__2430__A1 _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2981__A2 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1837_ _0775_ _0754_ _0857_ _0208_ _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2733__A2 _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1768_ _0813_ _0817_ _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1699_ _0747_ _0748_ _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_66_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1804__B _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2421__A1 _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput7 net7 qcos vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_48_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2488__A1 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2488__B2 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2660__A1 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2740_ _0227_ _0246_ _0268_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_12_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2671_ _0177_ _0192_ _0161_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1622_ _1345_ _1433_ _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_4
X_3223_ _0014_ net9 clknet_2_0__leaf_clk csTable.address\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2479__A1 _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3154_ _1433_ _0705_ _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_39_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3085_ _0479_ _0601_ _0632_ _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2105_ _1152_ _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2036_ _0778_ _0787_ _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_50_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2651__A1 _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2938_ _0312_ _0486_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2869_ _0407_ _0410_ _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_58_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1693__A2 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2642__A1 _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1709__B _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2945__A2 freeRunCntr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2881__A1 _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1684__A2 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3189__A2 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2936__A2 _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2723_ _0233_ _0239_ _0249_ _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2654_ _0172_ _0173_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2585_ _0095_ _0096_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1605_ _1345_ csTable.address\[5\] _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_3206_ _0028_ net10 clknet_2_3__leaf_clk freeRunCntr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__2872__A1 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3137_ _0687_ _0691_ _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3068_ net2 _0597_ _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2019_ _0857_ _0890_ _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3035__I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1666__A2 _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2091__A2 _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2918__A2 _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3040__A1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2370_ _1425_ _1426_ _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2854__B2 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2854__A1 _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2606__A1 _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2082__A2 _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3031__A1 freeRunCntr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2706_ _1265_ _0231_ _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2790__B1 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2790__C2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2637_ _0146_ _0151_ _0152_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_2568_ _1267_ _0078_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_59_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2499_ _1567_ _1568_ _1569_ _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3098__A1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1648__A2 _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2073__A2 _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3022__A1 freeRunCntr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3089__A1 _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1639__A2 _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2064__A2 _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1811__A2 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1870_ _0827_ _0774_ _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1683__I _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2422_ _1483_ _1484_ _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1878__A2 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2353_ _1406_ _1407_ _1408_ _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2284_ _1290_ _1292_ _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_64_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2055__A2 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1802__A2 _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3004__A1 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1999_ _0054_ _0761_ _1576_ _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2285__A2 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2971_ _0470_ _0476_ _0560_ _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2037__A2 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1922_ _0450_ _0967_ _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1853_ _0763_ _0827_ _0902_ _0754_ _0651_ _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_1784_ _0750_ _0833_ _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2405_ _1465_ _1441_ _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_29_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2336_ _1143_ _1146_ _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2267_ _0373_ _1310_ _1156_ _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2198_ _0747_ _0748_ _1197_ _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1787__B2 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1787__A1 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1711__A1 _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1778__A1 _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1950__A1 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3170_ csTable.address\[5\] _0718_ _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1702__A1 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2121_ _1162_ _1167_ _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2052_ freeRunCntr\[4\] _1056_ _1067_ _0882_ _1100_ _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_47_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2258__A2 _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2954_ freeRunCntr\[4\] _0491_ _0500_ _0502_ _0503_ _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_1905_ _0954_ net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2885_ _0424_ _0427_ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_30_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1836_ _0592_ _0765_ _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1767_ _0814_ _0815_ _0816_ _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2194__A1 _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1941__A1 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1698_ _0679_ _0746_ _1378_ _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_66_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2319_ _1280_ _1325_ _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_72_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2249__A2 _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3206__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2185__A1 _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput8 net8 qsin vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__1932__A1 _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2670_ _0181_ _0179_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1621_ _1554_ _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__2176__A1 _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1923__A1 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3222_ _0013_ net9 clknet_2_0__leaf_clk csTable.address\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_67_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3153_ freeRunCntr\[17\] _0703_ _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input3_I divSel[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2104_ _1143_ _1146_ _1097_ _1151_ _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_3084_ _0601_ _0639_ _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2035_ _0849_ _0991_ _1083_ _0738_ _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__3229__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1640__B _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2100__A1 sigRom.address\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2937_ _0354_ _0485_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2868_ _0408_ _0409_ _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2799_ _0289_ _0309_ _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1819_ _0763_ _1598_ _0783_ _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1914__A1 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2158__A1 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2330__B2 _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2881__A2 _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1887__S _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1686__I _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2722_ _0234_ _0238_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2397__A1 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2653_ _0166_ _0168_ _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2584_ _0095_ _0096_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1604_ _1367_ _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_67_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3205_ _0027_ net10 clknet_2_0__leaf_clk freeRunCntr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3136_ _0688_ _0683_ _0690_ _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3067_ net3 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_27_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2018_ _1065_ _1066_ _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_42_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2388__A1 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1899__B1 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2379__B2 _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2379__A1 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3040__A2 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2000__B1 _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2854__A2 _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2705_ _1025_ _1151_ _1305_ _0996_ _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__2790__A1 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2790__B2 _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2636_ _1079_ _0113_ _0147_ _1379_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2567_ _1267_ _0078_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2542__A1 _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2498_ _1562_ _1566_ _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__3098__A2 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1648__A3 _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3119_ _0672_ _0673_ _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2058__B1 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1639__A3 _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2834__B _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2049__B1 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2421_ _1340_ _1427_ _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_43_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2352_ _1402_ _1404_ _1405_ _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_69_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2283_ _1330_ _1331_ _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1998_ _1565_ _0849_ _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2619_ _0129_ _0134_ _0135_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__2515__A1 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1717__C _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2829__B _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2970_ _0519_ _0520_ _0467_ _0521_ _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1921_ freeRunCntr\[15\] _0969_ _0965_ freeRunCntr\[14\] _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__2442__B1 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1852_ _0175_ _0582_ _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1783_ _0783_ _0821_ _0164_ _0832_ _0779_ _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__3226__RN net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout9 net12 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_2404_ _1432_ _1436_ _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3170__A1 csTable.address\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2335_ _1097_ _1150_ _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2266_ _0472_ _1197_ _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2197_ _1236_ _1244_ _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2520__I1 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1787__A2 _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3217__RN net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3161__A1 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1711__A2 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1778__A2 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2727__A1 _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3208__RN net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1950__A2 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1702__A2 _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2120_ _1162_ _1167_ _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2051_ _1089_ _1098_ _1099_ _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_47_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2953_ freeRunCntr\[3\] _0501_ _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_22_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1904_ _0516_ _0953_ _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2884_ _0425_ _0426_ _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_30_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1835_ freeRunCntr\[3\] _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1766_ freeRunCntr\[12\] _0812_ _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2194__A2 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1697_ _1378_ _0679_ _0746_ _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2318_ _1280_ _1325_ _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2249_ _1235_ _1255_ _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1820__C _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2957__A1 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2709__A1 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1932__A2 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3134__A1 freeRunCntr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1696__A1 _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1696__B2 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1620_ _1543_ _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__2176__A2 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3221_ _0012_ net9 clknet_2_0__leaf_clk csTable.address\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__1687__A1 _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3152_ _0704_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2103_ _1150_ _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_3083_ net2 net1 _0624_ _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2034_ _0571_ _0937_ _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_54_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2939__A1 _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2936_ _1533_ _0217_ _0350_ _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2939__B2 _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2867_ _0385_ _0383_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1611__A1 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1818_ _0763_ _0849_ _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2798_ _0289_ _0309_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1749_ _0795_ _0798_ _1400_ _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1678__A1 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1602__A1 _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2158__A2 _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3107__A1 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1669__A1 freeRunCntr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1841__A1 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2721_ _0221_ _0247_ _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_8_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2652_ _1432_ _0171_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_8_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2583_ _0049_ _0050_ _0052_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_1603_ _1356_ _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_3204_ _0026_ net9 clknet_2_1__leaf_clk freeRunCntr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__2321__A2 _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3135_ freeRunCntr\[13\] _0681_ _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3066_ _0623_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2017_ _1058_ _1061_ _1064_ _0395_ _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__2085__A1 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2919_ _0355_ _0357_ _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1826__B _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1899__A1 freeRunCntr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1899__B2 freeRunCntr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1823__A1 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2379__A2 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3040__A3 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3219__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2000__B2 _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2303__A2 _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1814__A1 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2704_ _0815_ _1314_ _1357_ _1358_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2790__A2 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2635_ _0146_ _0151_ _0152_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2566_ _0073_ _0075_ _0077_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2542__A2 _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2497_ _1538_ _1545_ _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1648__A4 _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3118_ _0624_ _0653_ _0615_ _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3049_ _0596_ _0599_ _0606_ _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2058__B2 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2058__A1 freeRunCntr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1805__A1 _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2297__A1 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_2_2__f_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2049__B2 freeRunCntr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2049__A1 freeRunCntr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2221__A1 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2420_ _1290_ _1481_ _1482_ _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2351_ _1387_ _1386_ _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2282_ _1295_ _1324_ _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1997_ _0849_ _0785_ _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2212__A1 _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2763__A2 _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2618_ _0100_ _0101_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2549_ _0038_ _0057_ _0058_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1962__B1 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1920_ _0395_ _0968_ _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2442__B2 _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2442__A1 _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1851_ _0885_ _0900_ _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1782_ _0175_ _0186_ _0698_ _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2403_ _1462_ _1463_ _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2334_ _1300_ _1385_ _1386_ _1387_ _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2265_ _1311_ _1312_ _1254_ _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_65_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2196_ _1239_ _1243_ _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1795__I0 _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3161__A2 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2424__A1 _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2727__A2 _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2050_ freeRunCntr\[3\] _1097_ _1056_ freeRunCntr\[4\] _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_19_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2952_ freeRunCntr\[3\] _0501_ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1903_ _0549_ _0819_ _0952_ _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_15_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2883_ _0472_ _1317_ _1318_ _0373_ _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_1834_ _0863_ _0864_ _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_1765_ _0792_ _0793_ _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1696_ _0450_ _0722_ _0744_ _0745_ _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1941__A3 _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2317_ _1329_ _1369_ _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2248_ _1235_ _1255_ _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2179_ _1220_ _1222_ _1226_ _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_25_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2709__A2 _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1917__B1 _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2893__A1 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2645__A1 _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3125__A2 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3220_ _0010_ net9 clknet_2_0__leaf_clk csTable.address\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3151_ freeRunCntr\[17\] _0703_ _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1687__A2 _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2102_ _1148_ _1149_ _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3082_ _0638_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2033_ _0651_ _1080_ _1081_ _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__2636__A1 _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2636__B2 _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2939__A2 _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2935_ _0349_ _0482_ _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3061__A1 freeRunCntr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2866_ _0379_ _0382_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1817_ _1422_ _1444_ _1488_ _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2797_ _0328_ _0331_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_7_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2572__B1 _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1748_ _0796_ _0797_ _0285_ _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1679_ _1466_ _1433_ _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_4
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2627__A1 _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3104__B freeRunCntr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3052__A1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1602__A2 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1669__A2 _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1741__C _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1841__A2 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2720_ _0229_ _0232_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2651_ _1079_ _1590_ _0170_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1602_ _1323_ _1345_ _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2582_ _0082_ _0093_ _0094_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_4_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1932__B _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3203_ _0022_ net9 clknet_2_0__leaf_clk freeRunCntr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_67_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3134_ freeRunCntr\[13\] _0681_ _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3065_ _0618_ _0621_ _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2016_ _0395_ _1058_ _1061_ _1064_ _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XANTENNA__2085__A2 _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2918_ _0445_ _0463_ _0464_ _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_31_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2849_ _0366_ _0367_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1899__A2 _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2076__A2 sigRom.address\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3025__A1 freeRunCntr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3040__A4 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2000__A2 _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1814__A2 _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2703_ _1354_ _1364_ _1362_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2634_ _0116_ _0118_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2565_ _1535_ _1541_ _1596_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2378__I0 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2496_ _1562_ _1566_ _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_67_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3117_ freeRunCntr\[12\] _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3048_ freeRunCntr\[1\] _0598_ _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2058__A2 _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1805__A2 _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1837__B _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2049__A2 _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1980__A1 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2350_ _1402_ _1404_ _1405_ _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2281_ _1298_ _1322_ _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1996_ _1323_ _1044_ _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_20_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1971__A1 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2617_ _0100_ _0130_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2548_ _0055_ _0056_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1723__A1 _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2479_ _1173_ _1446_ _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3209__CLK clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1962__A1 _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1962__B2 _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2442__A2 _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1850_ _0898_ _0899_ _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_4
X_1781_ _0826_ _0829_ _0830_ _0602_ _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__1953__A1 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1953__B2 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2402_ _1456_ _1405_ _1407_ _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__1705__A1 _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2333_ _0770_ _1248_ _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2264_ _1247_ _1249_ _1310_ _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_65_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2195_ _1240_ _1242_ _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2130__A1 _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1979_ _1026_ _1027_ _0439_ _0230_ _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_4_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1795__I1 _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3107__B _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2011__B _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2681__B _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2424__A2 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1935__A1 _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2360__A1 _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2951_ _1430_ _0489_ _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1902_ _0818_ _0949_ _0950_ _0951_ _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_2882_ _0965_ _1304_ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1833_ freeRunCntr\[4\] _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1764_ freeRunCntr\[11\] _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1926__A1 freeRunCntr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1695_ _1389_ _0087_ _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_2316_ _1332_ _1368_ _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_57_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2247_ _1283_ _1294_ _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2178_ _1223_ _1225_ _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1896__I freeRunCntr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1917__A1 freeRunCntr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1917__B2 freeRunCntr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2342__A1 _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2893__A2 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3070__A2 _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1755__B _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3150_ freeRunCntr\[16\] _0701_ _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2333__A1 _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2884__A2 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3081_ _0634_ _0637_ _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2101_ sigRom.address\[1\] _1147_ _1115_ _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2032_ _0778_ _1047_ _0991_ _0917_ _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_35_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2934_ _0480_ _0481_ _0353_ _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2865_ _0403_ _0405_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1816_ _0778_ _0802_ _0651_ _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2796_ _0291_ _0308_ _0330_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2572__B2 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2572__A1 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1747_ _0065_ _1598_ _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1678_ _1422_ _1576_ _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2324__A1 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2875__A2 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3120__B freeRunCntr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3052__A2 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2563__A1 _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2079__B1 _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2650_ _1536_ _1590_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1601_ _1334_ _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_59_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2581_ _0090_ _0092_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3202_ _0011_ net9 clknet_2_0__leaf_clk freeRunCntr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__2857__A2 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input1_I divSel[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3133_ _0685_ _0686_ _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3064_ _0619_ _0613_ _0620_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2015_ _1389_ _1062_ _0987_ _1063_ _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_35_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3034__A2 _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2917_ _0312_ _0337_ _0350_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2848_ _0383_ _0387_ _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2779_ _0280_ _0311_ _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2076__A3 _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2536__A1 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3016__A2 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2702_ _0218_ _0222_ _0226_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_13_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2633_ _0149_ _0150_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2104__B _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2564_ _1132_ _0074_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2378__I1 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1943__B _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2495_ _1563_ _1564_ _1504_ _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3116_ _0671_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3047_ freeRunCntr\[2\] _0604_ _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3007__A2 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1837__C _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2014__B _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2518__A1 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2949__B freeRunCntr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3191__A1 _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2206__B1 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2221__A3 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1980__A2 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2280_ _1283_ _1294_ _1328_ _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2996__A1 _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1938__B _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3229__RN net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1995_ _1040_ _1042_ _1043_ _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_2616_ _0106_ _0127_ _0128_ _0132_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__1971__A2 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2769__B _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3173__A1 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2547_ _0055_ _0056_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2920__A1 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2478_ _1538_ _1545_ _1546_ _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1723__A2 _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1962__A2 _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3164__A1 csTable.address\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2978__A1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1650__A1 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1780_ _0821_ _0743_ _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2401_ _1456_ _1458_ _1459_ _1460_ _1461_ _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__1705__A2 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2332_ _1246_ _0749_ _1385_ _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2263_ _1310_ _1247_ _1249_ _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_37_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2194_ _1067_ _1164_ _1241_ _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1940__C _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2130__A2 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1641__A1 _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1641__B2 _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1978_ _0821_ _0894_ _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1944__A2 _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3146__A1 freeRunCntr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2011__C _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2424__A3 _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1632__A1 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2188__A2 _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2360__A2 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1871__A1 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2950_ _0495_ _0498_ _0499_ _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2881_ _0969_ _1151_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1901_ freeRunCntr\[8\] _0848_ _0771_ _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1832_ freeRunCntr\[5\] _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_30_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2179__A2 _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1763_ freeRunCntr\[11\] _0794_ _0812_ freeRunCntr\[12\] _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1926__A2 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1694_ _0571_ _0730_ _0738_ _0742_ _0743_ _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_57_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2315_ _1347_ _1366_ _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_38_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2246_ _1286_ _1293_ _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_72_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2177_ _1056_ _1164_ _1224_ _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1614__A1 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1917__A2 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1853__A1 _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1853__B2 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1605__A1 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2581__A2 _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2333__A2 _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3080_ _0635_ _0628_ _0636_ _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2100_ sigRom.address\[1\] _1147_ _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2031_ _0778_ _0762_ _0631_ _0821_ _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2097__A1 _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1844__A1 _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2933_ _0346_ _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2864_ _0360_ _0378_ _0404_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2795_ _0293_ _0306_ _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1815_ _0863_ _0864_ _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1746_ _1554_ _0120_ _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__2021__A1 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2021__B2 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2572__A2 _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1677_ _0571_ _0592_ _0602_ _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2324__A2 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2229_ _1262_ _1270_ _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1700__I _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2017__B _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2563__A2 _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2079__B2 _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2079__A1 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1826__A1 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2003__A1 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1600_ csTable.address\[6\] _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2580_ _0090_ _0092_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3201_ _0000_ net9 clknet_2_1__leaf_clk freeRunCntr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_67_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2711__C1 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3132_ _0624_ _0653_ _0630_ _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3063_ freeRunCntr\[3\] _0610_ _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1817__A1 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2014_ _1554_ _0120_ _0153_ _0087_ _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2916_ _0460_ _0462_ _0215_ _0213_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__2242__A1 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2847_ _0385_ _0386_ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2778_ _0284_ _0310_ _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1729_ _0329_ _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_2_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1753__B1 _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1808__A1 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2233__A1 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1992__B1 _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2536__A2 _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2472__A1 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3016__A3 _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2701_ _0223_ _0225_ _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2632_ _0143_ _0145_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2104__C _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2563_ _1379_ _1432_ _0073_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_4_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2494_ _1458_ _1507_ _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3115_ freeRunCntr\[11\] _0668_ _0669_ _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_67_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3046_ net3 _0601_ _0603_ _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2215__A1 _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1853__C _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3191__A2 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2256__I _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2206__B2 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1965__B1 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3232__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2693__A1 _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3202__D _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2445__A1 _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1994_ _0428_ _1510_ _0874_ _0917_ _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_9_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2615_ _0129_ _0100_ _0130_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2546_ _1567_ _1568_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2477_ _1540_ _1544_ _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2785__B _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3029_ freeRunCntr\[14\] _0584_ _0585_ _0586_ _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_34_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2025__B _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2978__A2 _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1758__C _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1650__A2 _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2400_ _1161_ _1437_ _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_40_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2331_ _0879_ _0880_ _1197_ _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_2262_ _0373_ _1197_ _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2193_ _0406_ _1141_ _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2418__A1 _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1641__A2 _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1977_ _0131_ _0780_ _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1684__B _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2529_ _1595_ _0035_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1880__A2 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1632__A2 csTable.address\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2896__A1 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2648__A1 _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1871__A2 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2880_ _0392_ _0401_ _0422_ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1900_ _0560_ _0749_ _0770_ freeRunCntr\[10\] _0549_ _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_15_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1831_ _0879_ _0880_ _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_30_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1762_ _0810_ _0811_ _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_1693_ _1565_ _0698_ _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2314_ _1350_ _1365_ _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2245_ _1287_ _1290_ _1292_ _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__2639__A1 _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2176_ _0472_ _1197_ _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_38_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1614__A2 csTable.address\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1853__A2 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1605__A2 csTable.address\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2869__A1 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2030_ _1078_ _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2097__A2 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1844__A2 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3046__A1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2932_ _0445_ _0463_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_62_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2863_ _0364_ _0377_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2794_ _0314_ _0316_ _0327_ _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_1814_ _0858_ _0862_ _0417_ _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__2021__A2 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1745_ _1455_ _1499_ _0761_ _1532_ _0329_ _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__1780__A1 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1676_ _0329_ _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2332__I0 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2228_ _1183_ _1274_ _1275_ _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2159_ _1204_ _1205_ _1206_ _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3037__A1 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1771__A1 _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1872__B _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2079__A2 _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1826__A2 _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2251__A2 _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2003__A2 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1782__B _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3200_ _0741_ _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2711__B1 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2711__C2 _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3131_ freeRunCntr\[14\] _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3205__D _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3062_ freeRunCntr\[3\] _0610_ _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2013_ _0252_ _0738_ _0873_ _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_23_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2118__B _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2915_ _1431_ _0210_ _0211_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__2242__A2 _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2846_ _0332_ _0335_ _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2777_ _0286_ _0289_ _0309_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__2788__B _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1728_ _1532_ _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__1753__A1 _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1659_ _0406_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__1753__B2 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1867__B _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2233__A2 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1992__A1 _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1992__B2 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1621__I _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2700_ _0224_ _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1983__A1 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2631_ _1379_ _0148_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2562_ _1056_ _1379_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1735__A1 _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2493_ _1159_ _1505_ _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2535__I0 _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3114_ _0662_ _0665_ _0661_ _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_28_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3045_ net2 _0597_ _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2999__B1 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1687__B _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2215__A2 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2829_ _0969_ _1305_ _1340_ _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1726__A1 _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2151__A1 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2206__A2 _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1965__A1 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1965__B2 _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2142__A1 _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1993_ _0745_ _1041_ _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1956__A1 _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1954__C _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2614_ _0038_ _0057_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1708__A1 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2545_ _0051_ _0052_ _0053_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2476_ _1540_ _1544_ _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_68_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2133__A1 _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3028_ freeRunCntr\[13\] _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_70_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2092__I sigRom.address\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1947__A1 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2124__A1 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2832__C1 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2330_ _1128_ _1381_ _1382_ _1383_ _1129_ _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__1790__B _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2378__S _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2261_ _1299_ _1308_ _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2115__A1 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2192_ _1045_ _1150_ _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2126__B _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1976_ _0395_ _1024_ _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__1929__A1 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2528_ _1595_ _0035_ _1121_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2459_ _1454_ _1476_ _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_56_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3222__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2593__A1 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2896__A2 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1830_ _0871_ _0878_ _1367_ _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1761_ _0799_ _0809_ _1367_ _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1692_ _0582_ _1598_ _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2336__A1 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2313_ _1354_ _1364_ _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2244_ _1121_ _1263_ _1291_ _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_38_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2175_ _1067_ _1150_ _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1847__B1 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2571__S _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2575__A1 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1959_ _0582_ _1587_ _0761_ _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1714__I _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1624__I _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3046__A2 _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_50_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2931_ freeRunCntr\[6\] _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0_clk clk clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_30_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2862_ _0389_ _0402_ _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2793_ _0317_ _0319_ _0326_ _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__2557__A1 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1813_ _0417_ _0858_ _0862_ _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_30_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1744_ _0792_ _0793_ _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_7_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1780__A2 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1675_ _0175_ _0582_ _0186_ _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1962__C _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3210__RN net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2227_ _1232_ _1273_ _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2332__I1 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2158_ _1196_ _1203_ _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2089_ _1128_ _1135_ _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_41_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2796__A1 _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1771__A2 _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1872__C _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2720__A1 _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3201__RN net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2571__I1 _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2787__A1 _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2003__A3 _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2711__B2 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2711__A1 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3130_ _0684_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2386__S _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3061_ freeRunCntr\[4\] _0617_ _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2012_ _0906_ _1059_ _1060_ _0428_ _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_35_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2914_ _0206_ _0451_ _0452_ _0459_ _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
X_2845_ _0328_ _0331_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2776_ _0291_ _0308_ _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1727_ _0764_ _0773_ _0775_ _0776_ _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__1753__A2 _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1658_ _0395_ _1345_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2769__A1 _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1992__A2 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3194__A1 _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2154__C1 _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2630_ _1078_ _1489_ _0147_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2561_ _1265_ _0071_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1735__A2 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2492_ _1555_ _1560_ _1561_ _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2535__I1 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3113_ _0653_ _0667_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3044_ net4 _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_63_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2828_ _0365_ _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3176__A1 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2759_ _1120_ _0231_ _0256_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2923__A1 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1726__A2 _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2151__A2 _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3167__A1 csTable.address\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2142__A2 _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1653__A1 _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1992_ _0186_ _0806_ _0801_ _0689_ _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_9_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1807__I _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2613_ _0079_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1708__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2544_ _0049_ _0050_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2475_ _1541_ _1542_ _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_68_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1892__A1 _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3027_ _0580_ _0572_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_24_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1698__B _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2124__A2 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1883__B2 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1883__A1 _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2832__B1 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2832__C2 _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1938__A2 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1627__I _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2260_ _1302_ _1307_ _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_49_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2115__A2 _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2191_ _1212_ _1237_ _1238_ _1211_ _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1874__A1 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1975_ _0450_ _1019_ _1023_ _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1965__C _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2527_ _1597_ _0034_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2458_ _1500_ _1523_ _1524_ _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_29_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2389_ _1447_ _1448_ _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2290__A1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2593__A2 _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1856__A1 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1608__A1 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2033__A1 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1760_ _1356_ _0799_ _0809_ _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1691_ _1477_ _1576_ _0043_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_2312_ _1362_ _1363_ _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2243_ _0965_ _1007_ _1171_ _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1847__A1 _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2174_ _1213_ _1221_ _1199_ _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1847__B2 _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2024__A1 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1958_ _0395_ _1006_ _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__1783__B1 _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1889_ _1499_ _0824_ _0757_ _0854_ _0779_ _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_0_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1838__A1 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1886__B _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2015__A1 _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1905__I _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1829__A1 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2930_ freeRunCntr\[10\] _0473_ _0477_ _0560_ _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_62_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2254__A1 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1796__B _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2006__A1 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2861_ _0392_ _0401_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2792_ _0320_ _0325_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1812_ _0859_ _0860_ _0861_ _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1743_ _1367_ _0782_ _0791_ _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_7_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1674_ _1422_ _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3212__CLK clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2226_ _1232_ _1273_ _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2493__A1 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2157_ _1152_ _1168_ _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2088_ _1128_ _1135_ _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_53_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2787__A2 _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2003__A4 _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1635__I _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2711__A2 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3060_ _0601_ _0616_ _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2011_ _0796_ _0622_ _0867_ _0329_ _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2913_ _0448_ _0449_ _0454_ _0458_ _1584_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_2844_ _0379_ _0382_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1973__C _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2775_ _0293_ _0306_ _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1726_ _0763_ _1532_ _0329_ _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1657_ _1323_ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XANTENNA__1753__A3 _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2466__A1 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3189_ _1140_ _0733_ _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2209_ _1234_ _1256_ _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2218__A1 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2769__A2 _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2044__C _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1883__C _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2154__B1 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_2_0__f_clk clknet_0_clk clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__1680__A2 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1793__C _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2560_ _0063_ _0064_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2932__A2 _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2491_ _1558_ _1559_ _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2696__A1 _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3112_ _0624_ _0609_ _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2160__A3 _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3043_ _0600_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2827_ _0321_ _0322_ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2758_ _0287_ _0288_ _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1709_ _0175_ _0153_ _0698_ _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2689_ _1327_ _1374_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2439__A1 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3100__A2 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1653__A2 _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1991_ _1036_ _1037_ _1039_ _0098_ _0428_ _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_9_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2612_ _0080_ _0097_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2543_ _1597_ _0034_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2474_ _1132_ _1489_ _1487_ _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1979__B _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1892__A2 _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3026_ _0573_ _0576_ _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_63_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1733__I _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1883__A2 _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3085__A1 _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2832__A1 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2832__B2 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2348__B1 _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2899__A1 _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2190_ _1213_ _1214_ _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1874__A2 _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3076__A1 _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1974_ _1020_ _1021_ _1022_ _0439_ _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1981__C _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2526_ _0033_ _1594_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2457_ _1520_ _1522_ _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_68_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2388_ _1267_ _1380_ _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_68_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3009_ _0972_ _1304_ _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2290__A2 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1728__I _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1856__A2 _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3058__A1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1608__A2 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1638__I _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1690_ _1565_ _0582_ _0186_ _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_51_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1792__A1 _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2311_ _1355_ _1361_ _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2242_ _1288_ _1289_ _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2173_ _0945_ _1142_ _1184_ _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_65_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3049__A1 _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2647__I1 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2024__A2 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1957_ _0670_ _1002_ _1003_ _1005_ _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1783__A1 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1888_ _0783_ _0937_ _0230_ _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2509_ _1579_ _1580_ _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1774__A1 _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1829__A2 _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2860_ _0398_ _0400_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1811_ _0208_ _0828_ _0857_ _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2791_ _0323_ _0324_ _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1742_ _0782_ _0791_ _1367_ _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_11_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1673_ _0131_ _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2190__A1 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2225_ _1257_ _1272_ _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_26_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2156_ _1196_ _1203_ _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2087_ _1129_ _1134_ _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_53_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2245__A2 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2989_ _0423_ _0434_ _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1756__A1 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2705__B1 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2181__A1 _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2484__A2 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1747__A1 _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2010_ _0252_ _1038_ _0098_ _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_63_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2912_ _0127_ _0455_ _0456_ _0457_ _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_31_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1986__A1 _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2843_ _0314_ _0380_ _0381_ _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2774_ _0298_ _0305_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1738__A1 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1725_ _0142_ _0774_ _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1656_ freeRunCntr\[13\] _0318_ _0373_ freeRunCntr\[14\] _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2163__A1 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1910__A1 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2466__A2 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3188_ freeRunCntr\[27\] freeRunCntr\[28\] _0728_ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_26_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2208_ _1235_ _1245_ _1255_ _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_2139_ _1118_ _1186_ _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_4
XANTENNA__2218__A2 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1977__A1 _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2926__B1 freeRunCntr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2154__B2 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2154__A1 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1901__A1 freeRunCntr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1665__B1 _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1968__A1 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3202__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2490_ _1558_ _1559_ _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_4_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3111_ _0666_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3042_ _0596_ _0599_ _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1656__B1 _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1959__A1 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2826_ _0363_ _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_31_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2757_ _0248_ _0267_ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2384__A1 _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2688_ _1431_ _0210_ _0211_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1708_ _0730_ _0738_ _0757_ _0571_ _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1639_ _0175_ _0153_ _0186_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_48_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2439__A2 _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3225__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2375__A1 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2127__A1 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1990_ _0787_ _0754_ _1038_ _1521_ _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_13_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2611_ _0122_ _0125_ _0126_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2542_ _0049_ _0050_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2473_ _1175_ _1289_ _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2118__A1 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3025_ freeRunCntr\[13\] _0581_ _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1979__C _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2054__B1 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2809_ _0343_ _0344_ _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2357__A1 _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1889__C _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3085__A2 _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2832__A2 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2045__B1 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2596__A1 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2596__B2 _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2348__B2 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2348__A1 _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1874__A3 _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1973_ _0764_ _0827_ _0867_ _0934_ _0285_ _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__2339__A1 _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2525_ _1379_ _1591_ _1589_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2456_ _1520_ _1522_ _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_68_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2511__A1 _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2387_ _1175_ _1377_ _1446_ _1173_ _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_28_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3008_ _0417_ _1189_ _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3231__RN net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1856__A3 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3058__A2 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2805__A2 _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1792__A2 _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2741__A1 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2310_ _1355_ _1361_ _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__3222__RN net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2241_ _1131_ _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_25_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2172_ _1163_ _1166_ _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1956_ _0896_ _1004_ _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2024__A3 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1783__A2 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2980__A1 _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1887_ _0175_ _0582_ _1598_ _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3213__RN net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2508_ _1500_ _1523_ _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__2732__A1 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2439_ _1078_ _1176_ _1502_ _1503_ _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2015__A3 _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1675__S _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1774__A2 _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3204__RN net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1829__A3 _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1810_ _0670_ _0850_ _0571_ _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2790_ _0812_ _1317_ _1318_ _0794_ _0373_ _1252_ _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_4
X_1741_ _0784_ _0786_ _0788_ _0790_ _1400_ _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_1672_ freeRunCntr\[9\] _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2190__A2 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2224_ _1259_ _1271_ _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_38_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2155_ _1198_ _1201_ _1202_ _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_38_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2086_ _1132_ _1133_ _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2988_ _0528_ _0541_ _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_21_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1939_ _1587_ _0774_ _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2953__A1 freeRunCntr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2705__A1 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2705__B2 _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2181__A2 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2339__B _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1692__A1 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2074__B _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2944__A1 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1747__A2 _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3121__A1 freeRunCntr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2911_ _0200_ _0202_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_31_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1986__A2 _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2842_ _0316_ _0327_ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2773_ _0299_ _0304_ _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1738__A2 _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1724_ _1466_ _1411_ _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_1655_ _1356_ _0362_ _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_4
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2163__A2 _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1910__A2 _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2207_ _1165_ _1250_ _1254_ _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_54_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3187_ _0732_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2138_ _1115_ sigRom.address\[0\] _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2069_ sigRom.address\[1\] _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__1977__A2 _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2926__A1 freeRunCntr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2154__A2 _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1901__A2 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1665__B2 freeRunCntr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1665__A1 freeRunCntr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1701__B _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2090__A1 _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1968__A2 _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1662__I _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3110_ _0662_ _0665_ _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_67_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3041_ freeRunCntr\[1\] _0598_ _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_36_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1656__B2 freeRunCntr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1656__A1 freeRunCntr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1959__A2 _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2081__A1 _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2825_ _0360_ _0361_ _0326_ _0325_ _0320_ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_2756_ _0250_ _0266_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2687_ _1486_ _1529_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1707_ _1543_ _1444_ _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_1638_ _0142_ _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_58_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1895__A1 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout10 net11 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_10_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2072__A1 _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2375__A2 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2127__A2 _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1810__A1 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1657__I _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2610_ _0082_ _0093_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2541_ _1555_ _1560_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2771__C1 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2472_ _0749_ _1539_ _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2118__A2 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1877__A1 freeRunCntr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3024_ _0580_ _0572_ _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1629__A1 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2054__B2 _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1801__A1 _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2808_ _0275_ _0276_ _0272_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2739_ _0248_ _0267_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_3_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1868__A1 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2293__A1 _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2045__A1 _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2045__B2 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2348__A2 _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1859__A1 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2284__A1 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2036__A1 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1972_ _0689_ _0894_ _0779_ _0998_ _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2339__A2 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2524_ _1596_ _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3215__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2455_ _1471_ _1472_ _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_68_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2386_ _1017_ _1445_ _1267_ _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3007_ _0533_ _0534_ _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2027__A1 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2266__A1 _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2018__A1 _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1792__A3 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2240_ _0955_ _0968_ _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_65_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2171_ _1210_ _1218_ _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_38_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2009__A1 _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1955_ _0915_ _0759_ _0801_ _0827_ _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1886_ _0933_ _0935_ _0439_ _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2980__A2 _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2507_ _1549_ _1577_ _1578_ _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__2732__A2 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1940__B1 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2438_ _1156_ _1214_ _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2369_ _1425_ _1426_ _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_56_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2015__A4 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2420__A1 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1774__A3 _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1931__B1 _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1704__B _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2487__A1 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2239__A1 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1740_ _0764_ _0789_ _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1671_ _0483_ _0527_ _0538_ _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_7_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2223_ _1262_ _1270_ _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2154_ _0884_ _1187_ _1189_ _0900_ _1193_ _1154_ _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_38_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2085_ _1045_ _1126_ _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2987_ _0539_ _0540_ _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1938_ _0986_ _0757_ _0698_ _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1869_ _0916_ _0918_ _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2705__A2 _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2469__A1 _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1692__A2 _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3197__A2 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2944__A2 _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3121__A2 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2632__A1 _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2910_ _0194_ _0196_ _0198_ _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2841_ _0316_ _0327_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2772_ _0302_ _0303_ _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1723_ _1554_ _1587_ _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_7_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1654_ _1400_ _0274_ _0340_ _0351_ _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2206_ _1154_ _1187_ _1189_ _1194_ _1253_ _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3186_ freeRunCntr\[28\] _0731_ _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2137_ _1184_ _1160_ _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2068_ _1115_ _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__2623__A1 _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1665__A2 _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1701__C _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3040_ net2 _0597_ net3 net4 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__2302__B1 _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2853__A1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1656__A2 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2081__A2 _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2824_ _0317_ _0319_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2442__C _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2755_ _0221_ _0247_ _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2686_ _1483_ _1484_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1706_ _0750_ _0752_ _0755_ _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1637_ _1477_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1895__A2 _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3169_ csTable.address\[3\] _1411_ csTable.address\[4\] _0711_ _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__1802__B _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout11 net12 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2072__A2 _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3021__A1 freeRunCntr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2540_ _0046_ _0047_ _0048_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1673__I _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2771__C2 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2771__B1 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2471_ _0945_ _1142_ _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1877__A2 _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3079__A1 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3023_ _0556_ _0558_ _0559_ _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_48_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1629__A2 csTable.address\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2807_ _1329_ _1369_ _0342_ _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2738_ _0250_ _0266_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2669_ _0161_ _0177_ _0179_ _0181_ _0190_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__1868__A2 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2045__A2 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1859__A2 _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2036__A2 _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1971_ _1477_ _1422_ _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2595__I0 _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2523_ _1045_ _1541_ _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2454_ _1501_ _1518_ _1519_ _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2385_ _1017_ _1171_ _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput1 divSel[0] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3006_ _0972_ _1151_ _0536_ _0561_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1786__A1 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1710__A1 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2266__A2 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2018__A2 _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_0_clk_I clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1701__A1 _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2170_ _1216_ _1217_ _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_65_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1954_ _0778_ _0824_ _0765_ _0750_ _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1885_ _0902_ _0754_ _0934_ _0764_ _0779_ _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__2193__A1 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2506_ _1574_ _1575_ _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1940__B2 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2437_ _1157_ _1237_ _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1940__A1 _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2368_ _1183_ _1274_ _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2299_ _1348_ _1349_ _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2248__A2 _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1810__B _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1759__A1 _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3028__I freeRunCntr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1931__A1 _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1931__B2 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2487__A2 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2239__A2 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1998__A1 _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3205__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1670_ freeRunCntr\[13\] _0318_ _0384_ _0494_ _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2175__A1 _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1922__A1 _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1681__I _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2222_ _1263_ _1269_ _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2153_ _1199_ _1200_ _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2084_ _1035_ _1131_ _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__1989__A1 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2986_ _0529_ _0537_ _0530_ _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA_fanout11_I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1937_ _1554_ _0142_ _0153_ _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1868_ _0571_ _0821_ _0751_ _0917_ _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_1_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2166__A1 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1799_ _0054_ _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__1913__A1 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3228__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1715__B _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2840_ _0359_ _0378_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2632__A2 _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1676__I _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2771_ _0794_ _1317_ _1318_ _0770_ _1252_ _0318_ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_4
XANTENNA__2396__A1 _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1722_ freeRunCntr\[10\] _0770_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1653_ _0285_ _0208_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2205_ _0848_ _1252_ _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2856__C1 _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3185_ freeRunCntr\[27\] _0728_ _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2136_ _0792_ _0793_ _1158_ _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__3131__I freeRunCntr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2067_ sigRom.address\[2\] _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__2623__A2 _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2969_ _0416_ _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2387__B2 _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2387__A1 _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2139__A1 _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1898__B1 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3197__B _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1889__B1 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2302__A1 _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2853__A2 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2302__B2 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2823_ _0359_ _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2754_ _0227_ _0282_ _0283_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1705_ _0753_ _0754_ _0602_ _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2685_ _1584_ _0070_ _0072_ _0207_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1636_ _1477_ _0142_ _0153_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2030__I _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2541__A1 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3168_ _0717_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2119_ _1163_ _1166_ _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_54_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3099_ _0653_ _0654_ _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout12 net5 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3021__A2 freeRunCntr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2532__A1 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2599__A1 _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2771__A1 _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2771__B2 _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2470_ _1078_ _1534_ _1132_ _1537_ _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2523__A1 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3022_ freeRunCntr\[12\] _0550_ _0578_ _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3003__A2 _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2806_ _1332_ _1368_ _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2737_ _0257_ _0265_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2668_ _0172_ _0173_ _0189_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1619_ _1334_ _1466_ _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_4
X_2599_ _1432_ _0113_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1970_ _0641_ _0715_ _1009_ _1018_ _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2522_ _1589_ _1592_ _1594_ _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3225__RN net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2453_ _1516_ _1517_ _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2384_ _1129_ _1383_ _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_68_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput2 divSel[1] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3005_ _0425_ _0426_ _0535_ _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_36_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1786__A2 _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1808__B _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3216__RN net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1718__B _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2726__A1 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3207__RN net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1701__A2 _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1953_ _0796_ _0998_ _0999_ _1001_ _0857_ _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__2965__B2 freeRunCntr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1884_ _1554_ _0142_ _0054_ _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1628__B _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2505_ _1574_ _1575_ _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2193__A2 _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2436_ _1497_ _1498_ _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1940__A2 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3142__A1 freeRunCntr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2367_ _1401_ _1423_ _1424_ _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2298_ _1309_ _1321_ _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2194__B _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2956__A1 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2956__B2 freeRunCntr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2169__C1 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1931__A2 _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3044__I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1695__A1 _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1998__A2 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2947__A1 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2123__I _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2175__A2 _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2221_ _1264_ _1266_ _1268_ _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_66_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2883__B1 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2152_ _0794_ _0836_ _1197_ _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2083_ _1115_ _1130_ _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2985_ _0529_ _0530_ _0537_ _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1936_ _1323_ _0984_ _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__1610__A1 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1867_ _1554_ _1521_ _0329_ _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1798_ _0406_ _0847_ _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_4
XANTENNA__2166__A2 _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3115__A1 freeRunCntr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2419_ _1479_ _1480_ _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1677__A1 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1821__B _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3039__I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1668__A1 freeRunCntr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1840__A1 _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2770_ _0300_ _0301_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1721_ _0560_ _0749_ _0770_ freeRunCntr\[10\] _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2396__A2 _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1652_ _0131_ _0164_ _0329_ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_2_1__f_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3184_ _0729_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2204_ _1251_ _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_39_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2856__C2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2856__B1 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2135_ _1138_ _1181_ _1182_ _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2066_ _0974_ _0975_ _1114_ _0966_ net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_19_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2084__A1 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2968_ _0415_ _0411_ _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1919_ _0670_ _0351_ _0967_ _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2899_ _0414_ _0420_ _0443_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1816__B _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1898__B2 _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1777__I _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1822__A1 _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1726__B _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1889__B2 _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1889__A1 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2302__A2 _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1813__A1 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2822_ _0317_ _0319_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2753_ _0246_ _0281_ _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1704_ _1543_ _1576_ _1488_ _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_2684_ _0068_ _0069_ _0138_ _0204_ _0206_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__1636__B _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3218__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1635_ _1422_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3167_ csTable.address\[4\] _0716_ _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_64_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3098_ net2 _0597_ _0624_ _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_2118_ _1097_ _1164_ _1165_ _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2049_ freeRunCntr\[2\] _1079_ _1097_ freeRunCntr\[3\] _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__2057__A1 _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1804__A1 _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2048__A1 _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2332__S _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2220__A1 _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2771__A2 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3021_ freeRunCntr\[15\] freeRunCntr\[16\] _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2039__A1 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2805_ _1370_ _1373_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2736_ _0258_ _0264_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2211__A1 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2667_ _0113_ _0184_ _0188_ _0174_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1618_ _1521_ _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2598_ _1435_ _1289_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_59_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3219_ _0009_ net11 clknet_2_2__leaf_clk csTable.address\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_39_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2925__B _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1789__B1 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2886__I _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2521_ _1132_ _1593_ _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_5_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2452_ _1516_ _1517_ _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2383_ _1432_ _1436_ _1441_ _1440_ _1438_ _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3004_ _0465_ _0466_ _0412_ _0557_ _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
Xinput3 divSel[2] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_36_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2432__A1 _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1808__C _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2735__A2 _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2719_ _0242_ _0245_ _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1824__B _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2423__A1 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1734__B _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2662__A1 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1952_ _0991_ _0976_ _1000_ _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2965__A2 _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1883_ _0764_ _0775_ _0932_ _0802_ _0230_ _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__2520__S _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2504_ _1501_ _1518_ _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2435_ _1497_ _1498_ _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2366_ _1420_ _1421_ _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2297_ _1313_ _1320_ _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1819__B _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2169__B1 _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2169__C2 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1931__A3 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1695__A2 _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2644__A1 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2947__A2 _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2220_ _1017_ _1126_ _1267_ _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_23_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2883__A1 _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2883__B2 _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2151_ _0945_ _1184_ _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2082_ _1117_ _1118_ _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2984_ _0531_ _0536_ _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_21_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3060__A1 _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1935_ _0889_ _0976_ _0978_ _0983_ _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1866_ _0802_ _0789_ _0915_ _0743_ _0602_ _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__1610__A2 _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1797_ _0837_ _0840_ _0843_ _0846_ _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2418_ _1479_ _1480_ _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1677__A2 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2349_ _1190_ _1187_ _1189_ _1403_ _1193_ _0884_ _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1668__A2 _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2093__A2 _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1840__A2 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3042__A1 _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1720_ _0768_ _0769_ _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_11_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1651_ _1345_ csTable.address\[4\] _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_4
XFILLER_7_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2856__A1 _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3183_ freeRunCntr\[27\] _0728_ _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2203_ _1122_ _1192_ _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2856__B2 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2134_ _1170_ _1180_ _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2065_ _0997_ _1110_ _1113_ _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2608__A1 _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2084__A2 _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2967_ _0352_ _0358_ _0475_ _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2898_ _0436_ _0442_ _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1918_ _0857_ _0830_ _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1849_ _0888_ _0897_ _0417_ _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_69_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1822__A2 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2386__I0 _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1889__A2 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1742__B _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1813__A2 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2821_ _0355_ _0357_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2752_ _0246_ _0281_ _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1703_ _0175_ _0065_ _0186_ _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2683_ _1264_ _1585_ _1586_ _0205_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_1634_ _1444_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1652__B _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2829__A1 _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3166_ csTable.address\[3\] _1411_ _0711_ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2117_ _0373_ _1158_ _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3097_ _0601_ _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_39_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2057__A2 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2048_ _1323_ _1096_ _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__1804__A2 _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3006__A1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1827__B _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1740__A1 _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2048__A2 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2220__A2 _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1731__A1 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3020_ freeRunCntr\[14\] _0573_ _0576_ _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_48_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2039__A2 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1798__A1 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2804_ _0338_ _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2735_ _0261_ _0262_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2666_ _0185_ _0187_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1970__A1 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1617_ _1488_ _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2597_ _1159_ _0083_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1722__A1 freeRunCntr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3218_ _0008_ net11 clknet_2_2__leaf_clk freeRunCntr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_54_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3149_ _0702_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1789__A1 _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1789__B2 _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1961__A1 _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3208__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2520_ _1536_ _1078_ _1534_ _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1952__A1 _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2451_ _1464_ _1467_ _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2382_ _1438_ _1440_ _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_3003_ _0420_ _0557_ _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput4 divSel[3] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1930__B _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_2_1__f_clk clknet_0_clk clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_24_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2718_ _0243_ _0244_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2196__A1 _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1943__A1 _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2649_ _0166_ _0168_ _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_19_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1840__B _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2187__A1 _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1934__A1 _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1750__B _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2662__A2 _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1951_ _0764_ _0988_ _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1882_ _1565_ _0827_ _1532_ _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2503_ _1551_ _1572_ _1573_ _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2434_ _1121_ _1447_ _1448_ _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2365_ _1420_ _1421_ _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2350__A1 _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2296_ _1335_ _1346_ _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_71_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2169__B2 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2169__A1 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1916__A1 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2644__A2 _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1907__A1 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2883__A2 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2150_ _0812_ _1197_ _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2081_ _0996_ _1119_ _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_53_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2983_ _0532_ _0535_ _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_21_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2399__A1 _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1934_ _0285_ _0980_ _0981_ _0982_ _1389_ _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_1865_ _0043_ _1444_ _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1796_ _0844_ _0845_ _0428_ _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2417_ _1401_ _1423_ _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2348_ _1403_ _1187_ _1193_ _0900_ _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_2279_ _1286_ _1293_ _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2562__A1 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3004__C _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1825__B1 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1840__A3 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1650_ _1356_ _0307_ _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_4
XFILLER_7_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2305__A1 _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3182_ _0727_ _0724_ _0720_ _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2202_ _1247_ _1249_ _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2856__A2 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2133_ _1170_ _1180_ _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_66_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2064_ freeRunCntr\[12\] _0985_ _1112_ _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2966_ freeRunCntr\[10\] _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2897_ _0440_ _0441_ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1917_ freeRunCntr\[13\] _0962_ _0965_ freeRunCntr\[14\] _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1848_ _0417_ _0888_ _0897_ _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1779_ _0783_ _0828_ _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3156__I _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2544__A1 _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1813__A3 _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2820_ _0313_ _0356_ _0336_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2751_ _0268_ _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1702_ _0571_ _1598_ _0751_ _0230_ _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_8_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2682_ _1263_ _1525_ _1526_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_1633_ _0120_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1933__B _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2829__A2 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3165_ _0714_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3096_ _0652_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2116_ _1117_ _1144_ _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2047_ _0439_ _1091_ _1093_ _1095_ _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__3006__A2 _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2949_ freeRunCntr\[1\] _0492_ _0493_ freeRunCntr\[2\] _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__2765__A1 _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1827__C _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2004__B _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2517__A1 _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1740__A2 _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1731__A2 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2803_ _0312_ _0337_ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3228__RN net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2734_ _1157_ _1187_ _1189_ _1300_ _1212_ _1193_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_2665_ _0113_ _0184_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1970__A2 _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2596_ _0900_ _0108_ _0110_ _1385_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1616_ _1455_ _1499_ _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3172__A1 csTable.address\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1722__A2 _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3217_ _0007_ net9 clknet_2_0__leaf_clk freeRunCntr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3148_ freeRunCntr\[16\] _0701_ _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_27_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3079_ _0882_ _0626_ _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1789__A2 _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1838__B _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3219__RN net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1961__A2 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3163__A1 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1799__I _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1748__B _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2441__A3 _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2450_ _1513_ _1514_ _1515_ _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3154__A1 _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2901__A1 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2381_ _1439_ _1394_ _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_39_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3002_ _0468_ _0546_ _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput5 rst net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_64_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1640__A1 _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2717_ _0228_ _0240_ _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1943__A2 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2648_ _1402_ _0167_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3145__A1 freeRunCntr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2579_ _0045_ _0091_ _0047_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_59_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1631__A1 _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2187__A2 _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1698__A1 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1870__A1 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1950_ _0915_ _0743_ _0602_ _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1881_ freeRunCntr\[4\] _0865_ _0881_ _0882_ _0930_ _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__1622__A1 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2178__A2 _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2502_ _1570_ _1571_ _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2433_ _1491_ _1495_ _1496_ _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1689__A1 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2364_ _1229_ _1230_ _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_29_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2295_ _1338_ _1344_ _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_37_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1861__A1 _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1613__A1 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2169__A2 _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2341__A2 _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1852__A1 _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1907__A2 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1745__C _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2580__A2 _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1761__B _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2080_ _1121_ _1127_ _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1843__A1 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2982_ _0533_ _0534_ _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1933_ _0065_ _0773_ _0806_ _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1864_ freeRunCntr\[2\] _0913_ _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1795_ _0120_ _0054_ _1543_ _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2020__A1 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2308__C1 _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2416_ _1454_ _1476_ _1478_ _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2347_ _1367_ _0925_ _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_2278_ _1276_ _1326_ _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2087__A1 _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2011__A1 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2562__A2 _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1825__B2 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1825__A1 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1756__B _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2002__A1 _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2305__A2 _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3181_ freeRunCntr\[26\] _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2201_ _0318_ _0749_ _1248_ _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2132_ _1172_ _1179_ _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2063_ _0970_ _1111_ _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1816__A1 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2965_ _0488_ _0509_ _0514_ freeRunCntr\[8\] _0515_ _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_2896_ _0408_ _0407_ _0435_ _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1916_ _0955_ _0964_ _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_1847_ _0889_ _0891_ _0892_ _0895_ _0896_ _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_1778_ _0763_ _0827_ _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2544__A2 _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2471__A1 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2750_ _0269_ _0279_ _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2223__A1 _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1701_ _1565_ _1598_ _0689_ _0131_ _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2681_ _0133_ _0139_ _0199_ _0203_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1982__B1 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1632_ _1345_ csTable.address\[3\] _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_4
XTAP_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3233_ _0025_ net11 clknet_2_3__leaf_clk sigRom.address\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_66_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3164_ csTable.address\[3\] _0713_ _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_54_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3095_ _0647_ _0650_ _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2115_ _1056_ _1150_ _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_54_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2046_ _0439_ _1094_ _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2462__A1 _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2948_ _0210_ _0497_ _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2879_ _0366_ _0367_ _0402_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__1973__B1 _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2517__A2 _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2205__A1 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1731__A3 _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2444__A1 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2802_ _0313_ _0336_ _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2733_ _0259_ _0260_ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1955__B1 _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2664_ _0162_ _0165_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_8_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2595_ _0913_ _0108_ _1506_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1615_ _1477_ _1422_ _1488_ _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__3231__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3216_ _0006_ net10 clknet_2_3__leaf_clk freeRunCntr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_67_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2267__S _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3147_ _0699_ _0695_ _0700_ _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2683__A1 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1730__I0 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3078_ _0882_ _0626_ _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2029_ _1077_ _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_35_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3163__A2 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2426__A1 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2380_ _1077_ _1303_ _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3001_ _0436_ _0555_ _0545_ _0441_ _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3090__A1 freeRunCntr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1640__A2 _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2716_ _0223_ _0225_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2647_ _1556_ _0926_ _0108_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2578_ _0040_ _0041_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2408__A1 _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1849__B _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1698__A2 _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1603__I _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1870__A2 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3072__A1 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1880_ _0883_ _0884_ _0929_ _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1622__A2 _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2501_ _1570_ _1571_ _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2432_ _1492_ _1493_ _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1689__A2 _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2363_ _1417_ _1418_ _1419_ _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2294_ _1339_ _1343_ _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_49_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3063__A1 freeRunCntr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1613__A2 _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2271__C1 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3118__A2 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2012__C _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2629__A1 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1852__A2 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3054__A1 freeRunCntr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2868__A1 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3034__B _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1843__A2 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2981_ _1378_ _1317_ _1318_ _0472_ _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3045__A1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2399__A3 _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1932_ _0800_ _0754_ _0098_ _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1863_ _0911_ _0912_ _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_1794_ _0153_ _0142_ _0087_ _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2020__A2 _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2308__C2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2308__B1 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2415_ _1474_ _1475_ _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2346_ _0884_ _1142_ _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_2277_ _1278_ _1280_ _1325_ _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_72_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1834__A2 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3036__A1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2011__A2 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1770__A1 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1862__B _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2078__A2 _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1825__A2 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2002__A2 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1772__B _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1761__A1 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2200_ _1197_ _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_21_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3180_ _0726_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2710__B1 _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2131_ _1174_ _1178_ _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2062_ freeRunCntr\[13\] _0962_ _0975_ _0973_ _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_54_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1816__A2 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3018__A1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2964_ _0946_ _0487_ _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1915_ _0450_ _0963_ _0830_ _0959_ _0896_ _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_2895_ _0437_ _0438_ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1846_ _0428_ _0329_ _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1777_ _0186_ _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__1752__A1 _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1682__B _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2069__I sigRom.address\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2329_ _1121_ _1127_ _1381_ _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3009__A1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1857__B _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1991__A1 _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1991__B2 _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1743__A1 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2471__A2 _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1700_ _1400_ _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2680_ _0200_ _0202_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1982__A1 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1631_ _1532_ _0076_ _0098_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_8_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1734__A1 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3232_ _0024_ net11 clknet_2_3__leaf_clk sigRom.address\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3163_ _1411_ _0711_ _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input4_I divSel[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2114_ _0770_ _1155_ _1160_ _1161_ _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3094_ _0648_ _0643_ _0649_ _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2045_ _0230_ _0592_ _0754_ _0849_ _1063_ _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_50_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2462__A2 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1677__B _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2947_ _0460_ _0211_ _0496_ _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout9_I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2878_ _0403_ _0405_ _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1973__A1 _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1973__B2 _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1829_ _1367_ _0871_ _0878_ _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA__1725__A1 _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2150__A1 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2971__B _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2453__A2 _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2205__A2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1964__A1 _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1716__A1 _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1606__I _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2444__A2 _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2801_ _0332_ _0335_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2732_ _1025_ _1164_ _1143_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1955__B2 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1955__A1 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2900__I _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2663_ _0182_ _0183_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_8_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2594_ _0913_ _1248_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1614_ _1334_ csTable.address\[3\] _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__2380__A1 _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1960__B _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3215_ _0005_ net10 clknet_2_3__leaf_clk freeRunCntr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_67_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2132__A1 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3146_ freeRunCntr\[15\] _0697_ _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3077_ freeRunCntr\[6\] _0633_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1730__I1 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2028_ _0955_ _1076_ _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_35_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1946__A1 _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1854__C _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2371__A1 _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2257__I _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2426__A2 _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1937__A1 _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2362__A1 _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2114__A1 _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3000_ _0542_ _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_64_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3203__D _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3090__A2 _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1928__A1 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2715_ _0228_ _0240_ _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2050__B1 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2646_ _0162_ _0165_ _0163_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2577_ _0086_ _0088_ _0089_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3129_ _0586_ _0681_ _0683_ _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_27_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2026__B _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1919__A1 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2344__A1 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1759__C _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3221__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2583__A1 _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2500_ _1511_ _1512_ _1514_ _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_2431_ _1494_ _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2335__A1 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2362_ _1415_ _1416_ _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2293_ _1340_ _1342_ _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_56_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2271__B1 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2271__C2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2574__A1 _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2629_ _1078_ _1435_ _1289_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2326__A1 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2629__A2 _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2565__A1 _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2980_ _0969_ _1304_ _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3045__A2 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1931_ _0787_ _0979_ _0873_ _0807_ _0806_ _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_1862_ _0905_ _0910_ _1378_ _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1793_ _0826_ _0841_ _0842_ _0098_ _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2020__A3 _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2308__A1 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2308__B2 _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2414_ _1474_ _1475_ _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_69_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2345_ _1384_ _1398_ _1399_ _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2276_ _1295_ _1324_ _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_37_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3036__A2 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1770__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2538__A1 _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1761__A2 _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2710__A1 _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2710__B2 _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2130_ _1120_ _1177_ _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2061_ freeRunCntr\[11\] _0996_ _1007_ freeRunCntr\[10\] _1109_ _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_34_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3018__A2 _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2963_ _0512_ _0513_ _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1914_ _0340_ _0351_ _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2894_ _0421_ _0435_ _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1845_ _0893_ _0894_ _0757_ _0759_ _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1776_ _0054_ _0142_ _0774_ _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__1752__A2 _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1682__C _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2328_ _1121_ _1127_ _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_72_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2259_ _1035_ _1303_ _1306_ _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_65_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3009__A2 _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2768__A1 _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1743__A2 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2759__A1 _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1982__A2 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1630_ _0087_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__1734__A2 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3206__D _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3231_ _0023_ net10 clknet_2_3__leaf_clk sigRom.address\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3162_ _0712_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2113_ _0815_ _1142_ _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3093_ freeRunCntr\[7\] _0640_ _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2044_ _0582_ _0998_ _1092_ _0230_ _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__2998__A1 freeRunCntr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1670__A1 freeRunCntr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2462__A3 _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2946_ _1486_ _1529_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2877_ _0419_ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1973__A2 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1828_ _0857_ _0875_ _0877_ _0750_ _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__3175__A1 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1725__A2 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1759_ _0230_ _0803_ _0808_ _0439_ _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2150__A2 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1964__A2 _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3166__A1 csTable.address\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1716__A2 _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2913__B2 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1652__A1 _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2800_ _0286_ _0333_ _0334_ _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2731_ _1007_ _1151_ _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2662_ _1078_ _1289_ _0108_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3157__A1 _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2593_ _1159_ _0083_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1613_ _1334_ _1466_ _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_4
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2904__A1 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2380__A2 _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3214_ _0004_ net10 clknet_2_1__leaf_clk freeRunCntr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_67_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3145_ freeRunCntr\[15\] _0697_ _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3076_ _0601_ _0632_ _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1891__A1 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2027_ _0670_ _1071_ _1072_ _1075_ _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1688__B _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1643__A1 _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1643__B2 _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2929_ _0470_ _0476_ _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2199__A2 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3148__A1 freeRunCntr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1882__A1 _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1937__A2 _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3139__A1 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1617__I _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2362__A2 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2114__A2 _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1873__A1 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1625__A1 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1928__A2 _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2714_ _0233_ _0239_ _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2050__A1 freeRunCntr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2050__B2 freeRunCntr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2645_ _1506_ _0140_ _0163_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2576_ _0084_ _0085_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_59_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1864__A1 freeRunCntr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3128_ _0674_ _0677_ _0682_ _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_27_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3059_ net3 _0615_ _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1616__A1 _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2041__A1 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2042__B _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1775__C _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2032__A1 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2583__A2 _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2430_ _1492_ _1493_ _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2335__A2 _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2361_ _1384_ _1396_ _1397_ _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_2292_ _1288_ _1173_ _1341_ _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2099__A1 _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1846__A1 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1966__B _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2271__A1 _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2271__B2 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2023__A1 _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2574__A2 _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2628_ _0144_ _0145_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2326__A2 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2559_ _1583_ _1588_ _0068_ _0069_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1837__A1 _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2262__A1 _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2014__A1 _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1828__A1 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1630__I _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1930_ _1554_ _0054_ _1521_ _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1861_ _1378_ _0905_ _0910_ _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__2005__A1 _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1792_ _0120_ _0142_ _0761_ _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_6_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2308__A2 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2413_ _1417_ _1418_ _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2344_ _1396_ _1397_ _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_69_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2275_ _1298_ _1322_ _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1819__A1 _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2492__A1 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3036__A3 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2244__A1 _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3211__CLK clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2483__A1 _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2235__A1 _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2710__A2 _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2060_ _1107_ _1108_ _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2474__A1 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3018__A3 _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2962_ _0356_ _0511_ _0337_ _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1913_ _0955_ _0961_ _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_2893_ _0408_ _0407_ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1844_ _0175_ _0252_ _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1775_ _1499_ _0824_ _0631_ _0778_ _0779_ _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_69_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2327_ _1377_ _1380_ _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2258_ _1045_ _1304_ _1305_ _1025_ _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2189_ _0848_ _1197_ _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2217__A1 _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2768__A2 _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2940__A2 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1743__A3 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1900__B1 _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1783__C _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1734__A3 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3230_ _0021_ net10 clknet_2_3__leaf_clk sigRom.address\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XANTENNA__2695__A1 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3161_ _1411_ _0711_ _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2112_ _1156_ _1157_ _1159_ _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3092_ freeRunCntr\[7\] _0640_ _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2447__A1 _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2043_ _0763_ _0131_ _0827_ _0842_ _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__1670__A2 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2945_ freeRunCntr\[2\] freeRunCntr\[1\] _0492_ _0493_ _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_13_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2876_ _0416_ _0418_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1827_ _0876_ _0707_ _0715_ _1499_ _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1758_ _0263_ _0805_ _0806_ _0807_ _0098_ _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_1689_ _0689_ _0707_ _0715_ _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2438__A1 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1868__C _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1884__B _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3166__A2 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2429__A1 _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1652__A2 _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2730_ _0236_ _0237_ _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2601__A1 _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2661_ _1078_ _0108_ _1556_ _0162_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__1794__B _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1612_ csTable.address\[1\] _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2592_ _0080_ _0097_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3213_ _0003_ net12 clknet_2_1__leaf_clk freeRunCntr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_67_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3144_ _0693_ _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3075_ _0624_ _0630_ _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1891__A2 _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3093__A1 freeRunCntr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2026_ _1073_ _1074_ _0670_ _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2928_ _0352_ _0358_ _0475_ _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2859_ _0370_ _0374_ _0399_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3148__A2 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2659__A1 _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1882__A2 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3084__A1 _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3139__A2 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1633__I _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1625__A2 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2713_ _0234_ _0238_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2050__A2 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2644_ _0926_ _1506_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2575_ _1132_ _0074_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3127_ _0672_ _0673_ _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1864__A2 _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3058_ net2 net1 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1616__A2 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2009_ _0896_ _1057_ _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2041__A2 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1791__A1 _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2360_ _1415_ _1416_ _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2291_ _1129_ _1290_ _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2099__A2 _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1846__A2 _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3048__A1 freeRunCntr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2271__A2 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1782__A1 _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2627_ _1385_ _0110_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2558_ _1172_ _1579_ _1580_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2489_ _1155_ _1505_ _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1837__A2 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2037__C _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2262__A2 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2014__A2 _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1773__A1 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1892__B _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2253__A2 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1860_ _0651_ _0907_ _0908_ _0909_ _0450_ _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_1791_ _1521_ _1587_ _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2412_ _1471_ _1472_ _1473_ _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2343_ _1396_ _1397_ _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2274_ _1309_ _1321_ _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1819__A2 _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2244__A2 _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1989_ _1477_ _1576_ _0787_ _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1755__A1 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2704__B1 _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2483__A2 _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1994__A1 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1746__A1 _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1906__I _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2171__A1 _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2474__A2 _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2961_ _0356_ _0337_ _0511_ _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1912_ _0450_ _0958_ _0960_ _0956_ _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2892_ _0421_ _0435_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1843_ _0849_ _0827_ _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1774_ _1565_ _0065_ _1587_ _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__1737__A1 _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2326_ _1056_ _1305_ _1379_ _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2257_ _1126_ _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2188_ _1223_ _1225_ _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2217__A2 _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1976__A1 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2331__B _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2940__A3 _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1900__B2 freeRunCntr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1900__A1 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1719__A1 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2392__A1 _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2144__A1 sigRom.address\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3160_ _0708_ _0709_ _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2695__A2 _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2467__I _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3091_ _0645_ _0646_ _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2111_ _0941_ _0942_ _1158_ _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_2042_ _0790_ _1090_ _0602_ _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2447__A2 _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1958__A1 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2944_ _0460_ _0211_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2875_ _0409_ _0407_ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1974__C _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3201__CLK clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1826_ _1477_ _0142_ _0054_ _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2383__B2 _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2383__A1 _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1757_ _0153_ _0631_ _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1688_ _0252_ _1587_ _0098_ _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_57_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2309_ _1359_ _1360_ _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1894__B1 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2438__A2 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2326__B _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1949__A1 _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2045__C _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3166__A3 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2374__A1 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2126__A1 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1885__B1 _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3224__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2660_ _1078_ _0162_ _0180_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1611_ _1422_ _1444_ _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2591_ _0079_ _0102_ _0103_ _0104_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_5_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2117__A1 _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3212_ _0002_ net12 clknet_2_1__leaf_clk freeRunCntr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XANTENNA_input2_I divSel[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3143_ _0696_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3074_ net2 _0597_ _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_35_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2025_ _0778_ _0800_ _0651_ _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1891__A3 _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2927_ _0388_ _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2053__B1 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2858_ _0371_ _0372_ _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2789_ _0321_ _0322_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1809_ _0750_ _0263_ _0807_ _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_2_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3084__A2 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2347__A1 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1873__A3 _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1789__C _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2712_ _0236_ _0237_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2643_ _1590_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2574_ _0084_ _0085_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_59_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3126_ _0680_ _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_70_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3057_ _0614_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2008_ _0852_ _0876_ _1048_ _0252_ _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2329__A1 _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3230__RN net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2568__A1 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1791__A2 _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3221__RN net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1644__I _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2290_ _0972_ _1171_ _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_37_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2008__B1 _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1782__A2 _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1982__C _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2626_ _0143_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2731__A1 _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2557_ _1265_ _0066_ _0067_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3212__RN net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2488_ _1194_ _1556_ _1557_ _1159_ _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_28_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3109_ _0663_ _0656_ _0664_ _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1729__I _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2014__A3 _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3203__RN net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1790_ _0838_ _0839_ _1389_ _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2411_ _1469_ _1470_ _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2342_ _1120_ _1136_ _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2273_ _1313_ _1320_ _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_52_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1988_ _0867_ _0934_ _0087_ _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2952__A1 freeRunCntr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1755__A2 _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2609_ _0123_ _0124_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2704__A1 _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_2_2__f_clk clknet_0_clk clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__1691__A1 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1994__A2 _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2943__A1 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1746__A2 _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3120__A1 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1682__A1 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2960_ _0354_ _0485_ _0510_ _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2891_ _0423_ _0434_ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_63_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1911_ _0745_ _0959_ _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1842_ _0571_ _0849_ _0631_ _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1773_ _0778_ _0820_ _0822_ _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1737__A2 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2147__C1 _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1832__I freeRunCntr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2325_ _1065_ _1066_ _1289_ _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_27_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2256_ _1164_ _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_53_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1988__B _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2187_ _1216_ _1217_ _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1976__A2 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2153__A2 _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1900__A2 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1664__A1 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2208__A3 _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3169__A1 csTable.address\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2916__A1 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3090_ freeRunCntr\[8\] _0601_ _0594_ _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2110_ _1116_ sigRom.address\[0\] _1118_ _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_54_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2041_ _0783_ _0988_ _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1655__A1 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2943_ _0460_ _0211_ _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2874_ _0415_ _0411_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2080__A1 _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1825_ _0778_ _0797_ _0872_ _0873_ _0874_ _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_1756_ _1477_ _0043_ _0120_ _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_1687_ _0175_ _0186_ _0698_ _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2308_ _0848_ _1317_ _1318_ _0836_ _0770_ _1252_ _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_4
XANTENNA__1894__A1 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1894__B2 freeRunCntr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2239_ _1172_ _1268_ _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1646__A1 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1949__A2 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2071__A1 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2374__A2 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1885__B2 _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2062__A1 freeRunCntr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1647__I _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1610_ _1334_ _1433_ _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_2590_ _0100_ _0101_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2117__A2 _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3211_ _0001_ net12 clknet_2_1__leaf_clk freeRunCntr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
X_3142_ freeRunCntr\[15\] _0693_ _0695_ _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1876__A1 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3073_ _0629_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1628__A1 _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2024_ _0571_ _0876_ _0757_ _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_62_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2926_ freeRunCntr\[11\] _0444_ _0469_ freeRunCntr\[10\] _0473_ _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2053__B2 freeRunCntr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2053__A1 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2857_ _0396_ _0397_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1800__A1 _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1808_ _0851_ _0853_ _0856_ _0857_ _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_40_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2788_ _0996_ _1304_ _1224_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1739_ _0175_ _0065_ _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_49_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1867__A1 _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1619__A1 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2292__A1 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2044__A1 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2347__A2 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2035__A1 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2035__B2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2711_ _0749_ _1317_ _1318_ _0848_ _1252_ _0794_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_4
X_2642_ _0155_ _0157_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2573_ _1539_ _0044_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_19_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3125_ _0624_ _0653_ _0625_ _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3056_ _0885_ _0610_ _0613_ _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2007_ _0395_ _1055_ _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_23_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2909_ _0136_ _0103_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2734__C1 _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2112__S _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3214__CLK clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2008__A1 _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2008__B2 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2625_ _0913_ _0140_ _0141_ _1402_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__1835__I freeRunCntr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2556_ _0063_ _0064_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2731__A2 _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2487_ _0926_ _0881_ _1248_ _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3108_ _0560_ _0653_ _0654_ _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_28_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3039_ net1 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_23_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1758__B1 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2486__A1 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2410_ _1451_ _1452_ _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_42_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2341_ _1152_ _1388_ _1392_ _1393_ _1395_ _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__1921__B1 _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2272_ _1316_ _1319_ _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2477__A1 _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2229__A1 _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1987_ _1521_ _0915_ _0641_ _1020_ _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2608_ _0119_ _0121_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2539_ _0040_ _0045_ _0041_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2468__A1 _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1994__A3 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2943__A2 _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1682__A2 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2890_ _0429_ _0433_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1910_ _0783_ _0164_ _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2631__A1 _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1841_ _0738_ _0873_ _0890_ _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1772_ _1532_ _0821_ _0779_ _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2147__C2 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2147__B1 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2324_ _1025_ _1171_ _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2255_ _1148_ _1149_ _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2186_ _1219_ _1227_ _1233_ _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2165__B _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2689__A1 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3169__A2 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2377__B1 _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2129__B1 _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2040_ freeRunCntr\[2\] _1079_ _1088_ freeRunCntr\[1\] _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2942_ _1375_ _0490_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_15_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2873_ _0386_ _0383_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1824_ _1422_ _1587_ _1521_ _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1755_ _0582_ _0804_ _0252_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1686_ _0120_ _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_2307_ _1357_ _1358_ _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1894__A2 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2238_ _1284_ _1244_ _1285_ _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2169_ _1194_ _1187_ _1193_ _0945_ _1189_ _0884_ _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2071__A2 _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3020__A1 freeRunCntr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1885__A2 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3087__A1 _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2834__A1 _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2062__A2 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2533__B _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3210_ _0032_ net12 clknet_2_1__leaf_clk freeRunCntr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_67_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3141_ _0687_ _0691_ _0694_ _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1876__A2 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3072_ _0882_ _0626_ _0628_ _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__3078__A1 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1628__A2 _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2023_ _0274_ _0612_ _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2925_ _0470_ _0471_ _0414_ _0416_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2053__A2 _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2856_ _0373_ _1317_ _1318_ _0318_ _1378_ _1252_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_4
XANTENNA__1800__A2 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1807_ _0779_ _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2787_ _0985_ _1151_ _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1738_ _0779_ _0787_ _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1669_ freeRunCntr\[16\] _1378_ _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_49_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2108__A3 _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1867__A2 _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1619__A2 _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2292__A2 _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1858__A2 _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2528__B _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2035__A2 _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2710_ _0235_ _1248_ _1304_ _1017_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__1794__A1 _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2641_ _0123_ _0124_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2572_ _0900_ _0042_ _0083_ _1159_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2338__A3 _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1849__A2 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3124_ _0678_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3055_ _0605_ _0607_ _0611_ _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_27_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2006_ _0750_ _1050_ _1054_ _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_63_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2173__B _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2908_ _0136_ _0103_ _0453_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__1785__A1 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2839_ _0364_ _0377_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2734__B1 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2734__C2 _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_6_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1776__A1 _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3089__B freeRunCntr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2008__A2 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1767__A1 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2624_ _0108_ _1556_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2555_ _0063_ _0064_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2192__A1 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2486_ _0926_ _1248_ _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3107_ _0653_ _0654_ _0560_ _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3038_ freeRunCntr\[0\] _0595_ _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1800__B _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1758__B2 _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2183__A1 _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1930__A1 _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2486__A2 _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1694__B1 _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1710__B _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1997__A1 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2174__A1 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2340_ _1078_ _1303_ _1394_ _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1921__B2 freeRunCntr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1921__A1 freeRunCntr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2271_ _0836_ _1317_ _1318_ _0943_ _0749_ _1252_ _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_4
XFILLER_28_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1988__A1 _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3204__CLK clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1986_ _1323_ _1034_ _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_20_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2401__A2 _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2607_ _1056_ _0113_ _0115_ _1535_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2538_ _1379_ _1591_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1912__A1 _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2469_ _1535_ _1536_ _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2468__A2 _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1994__A4 _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2156__A1 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1705__B _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3227__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1840_ _1565_ _0582_ _0827_ _0131_ _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_8_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1771_ _0065_ _1587_ _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__2395__A1 _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2147__A1 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1615__B _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2323_ _1276_ _1326_ _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_57_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2254_ _1165_ _1301_ _1247_ _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2185_ _1210_ _1218_ _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1969_ _0764_ _0937_ _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2200__I _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3169__A3 csTable.address\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2377__A1 _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2377__B2 _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2129__B2 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2129__A1 _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2301__A1 _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2941_ _1430_ _0489_ _0214_ _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2604__A2 _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2872_ _0352_ _0358_ _0413_ _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1823_ _1477_ _1576_ _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1754_ _1466_ _1433_ _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1685_ _1433_ _1411_ _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_2306_ _1314_ _0472_ _1184_ _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2237_ _1239_ _1243_ _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_65_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2168_ _1211_ _1215_ _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_65_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2099_ _1140_ _1118_ _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_21_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2071__A3 _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2531__A1 _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2834__A2 _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1702__C _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2306__S _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2598__A1 _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3140_ _0685_ _0686_ _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3071_ _0618_ _0621_ _0627_ _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2022_ _1068_ _1069_ _1070_ _0857_ _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_50_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2924_ _0415_ _0411_ _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2855_ _0393_ _0394_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1806_ _1499_ _0757_ _0854_ _0855_ _0750_ _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_2786_ _0302_ _0303_ _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1737_ _1433_ _1411_ _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_1668_ freeRunCntr\[16\] _1378_ _0505_ _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1599_ csTable.address\[7\] _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3069__A2 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1764__I freeRunCntr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3233__RN net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2440__B1 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2640_ _0154_ _0158_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1794__A2 _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2571_ _0865_ _0042_ _1506_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1674__I _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3224__RN net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3123_ _0674_ _0677_ _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3054_ freeRunCntr\[2\] _0604_ _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2005_ _1036_ _1051_ _1052_ _1053_ _1400_ _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_35_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2907_ _0105_ _0133_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2838_ _0368_ _0376_ _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2769_ _1007_ _1304_ _1165_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3215__RN net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2734__B2 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2734__A1 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2629__B _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2265__A3 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2973__A1 freeRunCntr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1776__A2 _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2973__B2 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1708__B _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2725__A1 _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3206__RN net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3150__A1 freeRunCntr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2964__A1 _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1767__A2 _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2623_ _1403_ _1142_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2554_ _1549_ _1577_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2192__A2 _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2485_ _1088_ _1305_ _1540_ _1553_ _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3106_ _0659_ _0661_ _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2495__A3 _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3037_ _0593_ _0594_ _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_36_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_2_0__f_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2912__B _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2707__A1 _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2183__A2 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1930__A2 _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1694__A1 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1694__B2 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1921__A2 _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2270_ _1147_ _1188_ _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_35_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1685__A1 _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1988__A2 _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1985_ _1028_ _1033_ _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2732__B _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2606_ _0119_ _0121_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2537_ _0040_ _0041_ _0045_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2468_ _1077_ _1289_ _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2399_ _1402_ _1404_ _1458_ _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1811__B _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2928__A1 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2156__A2 _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3105__A1 _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1770_ _0730_ _0738_ _0757_ _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2147__A2 _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2322_ _1327_ _1374_ _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2253_ _1139_ _1300_ _1142_ _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1658__A1 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2184_ _1229_ _1230_ _1231_ _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1631__B _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1830__A1 _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2462__B _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1968_ _0955_ _1016_ _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_1899_ freeRunCntr\[7\] _0836_ _0848_ freeRunCntr\[8\] _0948_ _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__2138__A2 sigRom.address\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1897__A1 freeRunCntr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1649__A1 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3169__A4 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2377__A2 _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2129__A2 _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1888__A1 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2301__A2 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2940_ _1485_ _0460_ _0211_ _1531_ _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2871_ _0412_ _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1822_ _1565_ _0582_ _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1753_ _1532_ _0800_ _0753_ _0801_ _0802_ _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_1684_ _0612_ _0660_ _0670_ _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2305_ _1378_ _1248_ _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2236_ _1236_ _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2167_ _1212_ _1213_ _1214_ _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2098_ _1077_ _1145_ _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2056__A1 freeRunCntr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1803__A1 _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3217__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2531__A2 _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2295__A1 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2047__A1 _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2598__A2 _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3070_ _0883_ _0601_ _0616_ _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2021_ _0796_ _0797_ _0805_ _0920_ _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_35_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2038__B2 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2038__A1 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2923_ _0465_ _0466_ _0388_ _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1797__B1 _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2854_ _0965_ _1151_ _1304_ _0962_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2785_ _0965_ _1305_ _1290_ _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1805_ _0763_ _1598_ _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1736_ _0230_ _0785_ _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1667_ _0384_ _0483_ _0494_ _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2966__I freeRunCntr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1721__B1 _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3199_ freeRunCntr\[0\] _0595_ _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2219_ _1025_ _1119_ _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_38_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2201__A1 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2440__A1 _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2440__B2 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2570_ _0081_ _0077_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_4_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3122_ _0675_ _0669_ _0676_ _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3053_ net3 _0601_ _0609_ _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__2259__A1 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2004_ _1047_ _0707_ _0779_ _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_48_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2906_ _1120_ _0071_ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2982__A2 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2837_ _0369_ _0375_ _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2768_ _0996_ _1151_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2699_ _0218_ _0222_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1719_ _0406_ _0756_ _0767_ _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA__2734__A2 _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1814__B _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1708__C _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2725__A2 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2489__A1 _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3150__A2 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2661__A1 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2622_ _0136_ _0103_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2553_ _0036_ _0061_ _0062_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__1924__B1 _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2484_ _1552_ _1246_ _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3105_ _0518_ _0624_ _0593_ _0603_ _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_3036_ net2 net1 net3 _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_51_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2652__A1 _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2404__A1 _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3132__A2 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1694__A2 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2882__A1 _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1685__A2 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1984_ _1400_ _1030_ _1031_ _1032_ _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_20_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2605_ _0086_ _0088_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2536_ _1194_ _0042_ _0044_ _1552_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2467_ _1534_ _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2398_ _1402_ _1404_ _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3019_ _0562_ _0566_ _0574_ _0575_ _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2625__A1 _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2625__B2 _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3041__A1 freeRunCntr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2321_ _1370_ _1373_ _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_33_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2252_ _0747_ _0748_ _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_65_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1658__A2 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2183_ _1207_ _1228_ _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2607__A1 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2607__B2 _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1830__A2 _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3032__A1 freeRunCntr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1967_ _1010_ _1012_ _1014_ _1015_ _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_1898_ _0931_ _0944_ _0945_ _0946_ _0947_ _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__1806__C _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2519_ _1379_ _1591_ _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1897__A2 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3099__A1 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2074__A2 sigRom.address\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1888__A2 _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1732__B _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2870_ _0388_ _0411_ _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_15_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1821_ _0866_ _0842_ _0439_ _0870_ _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_1752_ _0153_ _0186_ _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1683_ _1400_ _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_7_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2304_ _1316_ _1319_ _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2235_ _1263_ _1269_ _1282_ _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2166_ _0848_ _1158_ _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_38_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2029__I _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2097_ _1117_ _1144_ _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2056__A2 _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1803__A2 _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2999_ _0474_ _0478_ _0517_ _0526_ _0553_ _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_5_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1817__B _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2020_ _0797_ _0979_ _0807_ _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_62_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2922_ _0467_ _0419_ _0468_ _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_62_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2853_ _0972_ _1305_ _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2784_ _0300_ _0301_ _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1804_ _0065_ _0186_ _0698_ _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1735_ _1532_ _0631_ _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_7_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1666_ freeRunCntr\[16\] _1378_ _0472_ freeRunCntr\[15\] _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1721__A1 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1721__B2 freeRunCntr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3198_ _1144_ _0737_ _0740_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2218_ _1265_ _1177_ _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_26_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2149_ _1158_ _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_53_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1788__A1 _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2201__A2 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1960__A1 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1712__A1 _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1779__A1 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2440__A2 _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1951__A1 _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1703__A1 _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3121_ freeRunCntr\[11\] _0653_ _0667_ _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3052_ net2 net1 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2259__A2 _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2003_ _0252_ _0802_ _0773_ _0789_ _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_23_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3207__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2905_ _0205_ _0446_ _0448_ _0449_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_31_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2836_ _0370_ _0374_ _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_31_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2767_ _0261_ _0262_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2698_ _1339_ _1343_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1718_ _0756_ _0767_ _0417_ _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1649_ _1400_ _0241_ _0296_ _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1942__A1 _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1830__B _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1933__A1 _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2110__A1 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2621_ _0105_ _0133_ _0137_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2177__A1 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2552_ _0059_ _0060_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1924__A1 freeRunCntr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1924__B2 freeRunCntr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2483_ _0836_ _1248_ _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3104_ _0653_ _0658_ freeRunCntr\[10\] _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3035_ net4 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2101__A1 sigRom.address\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2819_ _0269_ _0279_ _0311_ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_11_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1915__A1 _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1915__B2 _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2340__A1 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1694__A3 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2882__A2 _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1983_ _0774_ _0832_ _0917_ _1389_ _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2398__A1 _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2604_ _0107_ _0111_ _0112_ _0116_ _0118_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_2535_ _1385_ _0881_ _0042_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2466_ _1045_ _1171_ _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_68_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2322__A1 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2397_ _0900_ _1457_ _1142_ _0945_ _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_68_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3018_ _0972_ _1304_ _0564_ _0563_ _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_36_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2561__A1 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3105__A3 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2616__A2 _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1675__I0 _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2320_ _1278_ _1371_ _1372_ _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2251_ _1240_ _1242_ _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2182_ _1138_ _1181_ _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_65_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1966_ _1532_ _0285_ _0800_ _1400_ _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1897_ freeRunCntr\[6\] _0943_ _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2518_ _1237_ _1590_ _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2449_ _1511_ _1512_ _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2059__B1 _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1806__B1 _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2074__A3 _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3023__A2 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2470__B1 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1820_ _0867_ _0868_ _0787_ _0869_ _0602_ _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_11_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1751_ _1488_ _0761_ _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1682_ _0622_ _0641_ _0651_ _1499_ _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2525__A1 _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2303_ _1351_ _1353_ _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2234_ _1266_ _1281_ _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1887__I0 _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2165_ _0810_ _0811_ _1141_ _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_53_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2096_ _1115_ _1123_ _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3005__A2 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2998_ freeRunCntr\[12\] _0550_ _0552_ _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1949_ _1565_ _0827_ _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2764__A1 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2516__A1 _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2921_ _0436_ _0442_ _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2852_ _0390_ _0376_ _0391_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2783_ _0298_ _0305_ _0315_ _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1803_ _0450_ _0852_ _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1734_ _0783_ _0730_ _0738_ _0208_ _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__3227__RN net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1665_ freeRunCntr\[14\] _0373_ _0472_ freeRunCntr\[15\] _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1721__A2 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2217_ _0985_ _1119_ _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_66_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3197_ _1124_ _0733_ _1118_ _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2148_ _1185_ _1195_ _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2079_ _1045_ _1119_ _1126_ _1067_ _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__1788__A2 _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3218__RN net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1712__A2 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1779__A2 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3209__RN net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1951__A2 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1703__A2 _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3120_ _0653_ _0667_ freeRunCntr\[11\] _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3051_ _0608_ _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2002_ _0763_ _0689_ _0285_ _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_63_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2967__A1 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2267__I0 _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2904_ _1264_ _1579_ _1580_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_2835_ _0371_ _0372_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2766_ _0294_ _0297_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2195__A2 _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2697_ _1340_ _0220_ _0221_ _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1717_ _0758_ _0760_ _0766_ _0670_ _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_1648_ _1400_ _0274_ _0285_ _1510_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__1942__A2 _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2958__A1 _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1933__A2 _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3135__A1 freeRunCntr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1697__A1 _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2110__A2 sigRom.address\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2949__A1 freeRunCntr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2620_ _0136_ _0103_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2551_ _0059_ _0060_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2177__A2 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1924__A2 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2482_ _1550_ _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1688__A1 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3103_ _0624_ _0603_ _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3034_ _0554_ _0588_ _0591_ net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1860__A1 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2818_ _0338_ _0354_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2749_ _0272_ _0277_ _0278_ _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2002__B _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1679__A1 _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2340__A2 _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3108__A1 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1842__A1 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1982_ _1499_ _0824_ _0622_ _0759_ _0715_ _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_20_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2603_ _0111_ _0117_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2534_ _0863_ _0864_ _1197_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_5_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2465_ _1431_ _1531_ _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2396_ _0911_ _0912_ _1251_ _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_68_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3017_ _0568_ _0570_ _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2086__A1 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2010__A1 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1824__A1 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1675__I1 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2001__B2 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2250_ _1245_ _1296_ _1297_ _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2181_ _1207_ _1228_ _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1965_ _0783_ _1013_ _0641_ _1455_ _0329_ _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__2240__A1 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1896_ freeRunCntr\[7\] _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_2517_ _1434_ _1289_ _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2448_ _1491_ _1494_ _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2487__B _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2379_ _1300_ _1237_ _1437_ _1184_ _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2059__B2 freeRunCntr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2059__A1 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1806__A1 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3023__A3 _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2241__I _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2534__A2 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2397__B _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2470__A1 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1750_ _1543_ _1576_ _1422_ _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__2222__A1 _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1681_ _0285_ _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_7_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2302_ _1175_ _1303_ _1145_ _1035_ _1352_ _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_57_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2289__A1 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2233_ _1264_ _1268_ _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1887__I1 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2164_ _0810_ _0811_ _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_26_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2095_ _1139_ _1142_ _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2997_ _0548_ _0551_ _0814_ _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2213__A1 _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1948_ freeRunCntr\[12\] _0985_ _0996_ freeRunCntr\[11\] _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2764__A2 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1879_ _0901_ _0928_ _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2516__A2 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2010__B _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3067__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_2_3__f_clk clknet_0_clk clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_62_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2920_ _0465_ _0466_ _0412_ _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2443__A1 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2443__B2 _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2851_ _0323_ _0324_ _0375_ _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2782_ _0299_ _0304_ _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1802_ _0153_ _1587_ _1521_ _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1733_ _0698_ _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_7_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1664_ _0417_ _0461_ _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2216_ _0962_ _1119_ _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
X_3196_ _0739_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2682__A1 _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2147_ _0900_ _1187_ _1189_ _1190_ _1193_ _1194_ _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_38_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2078_ _1122_ _1125_ _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__2434__A1 _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1788__A3 _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_2_3__f_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1828__C _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3230__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2167__S _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2425__A1 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1703__A3 _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3050_ _0605_ _0607_ _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_67_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2001_ _0822_ _1046_ _1049_ _0602_ _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_48_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output8_I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2903_ _1120_ _0071_ _0447_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_31_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2834_ _0985_ _1304_ _1241_ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2765_ _1263_ _0295_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2696_ _1340_ _1341_ _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1716_ _0762_ _0707_ _0765_ _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1647_ _0098_ _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3179_ freeRunCntr\[26\] _0725_ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2958__A2 _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1697__A2 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2110__A3 _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1749__B _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2550_ _1550_ _1572_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_56_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2481_ _1547_ _1548_ _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_49_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1688__A2 _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3102_ _0657_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3033_ _0589_ _0590_ _0578_ _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2535__S _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3062__A1 freeRunCntr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1999__I0 _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2817_ _0347_ _0353_ _0348_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2748_ _0275_ _0276_ _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2679_ _0079_ _0102_ _0201_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1679__A2 _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1851__A2 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3053__A1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3108__A2 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2167__I0 _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2095__A2 _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1842__A2 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1981_ _0131_ _0826_ _1029_ _0285_ _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_13_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2602_ _0107_ _0112_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2533_ _0039_ _1557_ _1159_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2464_ _1485_ _1530_ _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2395_ _1402_ _1404_ _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3016_ _0556_ _0558_ _0559_ _0572_ _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_24_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1824__A2 _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1760__A1 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2180_ _1219_ _1227_ _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2149__I _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1815__A2 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1964_ _0773_ _0775_ _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1937__B _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1895_ _0406_ _0835_ _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2516_ _1434_ _1237_ _1289_ _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2447_ _1511_ _1512_ _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1751__A1 _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2378_ _0749_ _1246_ _1214_ _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2059__A2 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1806__A2 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3008__A1 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1990__A1 _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1990__B2 _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1742__A1 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2397__C _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1601__I _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2470__A2 _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1981__A1 _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1680_ _0043_ _0631_ _0120_ _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2301_ _1007_ _1305_ _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2232_ _1257_ _1272_ _1279_ _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2163_ _0318_ _1158_ _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2094_ _1141_ _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2996_ _0414_ _0420_ _0443_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1947_ _0955_ _0995_ _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__1972__A1 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1878_ _0885_ _0900_ _0914_ _0927_ _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__2516__A3 _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1724__A1 _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2452__A2 _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1963__A1 _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1715__A1 _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2201__B _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2850_ _0368_ _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1801_ _0775_ _0850_ _0764_ _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2781_ _0294_ _0297_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1732_ _0777_ _0781_ _0439_ _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1663_ _0450_ _0340_ _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1954__A1 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1934__C _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1706__A1 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2111__B _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1950__B _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2215_ _0965_ _1171_ _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3195_ _1116_ _0737_ _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_26_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2146_ _0879_ _0880_ _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2077_ _1123_ _1124_ _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2979_ _0425_ _0426_ _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2005__C _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1945__A1 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1945__B2 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1881__B1 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2425__A2 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2189__A1 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1936__A1 _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1770__B _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2000_ _1047_ _0841_ _1048_ _1532_ _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2113__A1 _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2902_ _0063_ _0064_ _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_50_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2833_ _0962_ _1151_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2764_ _0962_ _1305_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1715_ _0763_ _0764_ _0230_ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1927__A1 _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2695_ _1288_ _1173_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1646_ _0252_ _0263_ _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2352__A1 _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1680__B _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2104__A1 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3178_ _0724_ _0720_ _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2129_ _1175_ _1131_ _1176_ _1035_ _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1918__A1 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1855__B _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2343__A1 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1697__A3 _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1909__A1 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2031__B1 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2480_ _1547_ _1548_ _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2334__A1 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3101_ _0560_ _0655_ _0656_ _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_3032_ freeRunCntr\[13\] _0581_ _0577_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1845__B1 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1999__I1 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2816_ _0341_ _0345_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3220__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2747_ _0275_ _0276_ _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2678_ _0106_ _0128_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1629_ _1345_ csTable.address\[4\] _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__2325__A1 _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2628__A2 _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3053__A2 _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2564__A1 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2167__I1 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1604__I _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1842__A3 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1980_ _0631_ _0689_ _0698_ _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2601_ _1534_ _0115_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2532_ _1159_ _0039_ _1557_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_5_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2307__A1 _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2463_ _1483_ _1484_ _1486_ _1529_ _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2394_ _1442_ _1443_ _1453_ _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3015_ _0568_ _0570_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_51_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2785__A1 _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1760__A2 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1963_ _0439_ _1011_ _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2776__A1 _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1894_ _0882_ _0881_ _0943_ freeRunCntr\[6\] _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2515_ _1264_ _1585_ _1586_ _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2446_ _1460_ _1461_ _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1751__A2 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2377_ _1434_ _1303_ _1176_ _1435_ _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_68_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2075__I _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3008__A2 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2519__A1 _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1990__A2 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3192__A1 _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1742__A2 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1981__A2 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2930__A1 freeRunCntr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2930__B2 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2300_ _1157_ _1310_ _1314_ _1315_ _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2231_ _1234_ _1256_ _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_65_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2162_ _1208_ _1209_ _1202_ _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_65_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2093_ _1115_ _1140_ _1123_ _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_38_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2995_ _0546_ _0547_ _0548_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1946_ _0450_ _0990_ _0994_ _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1877_ freeRunCntr\[2\] _0913_ _0926_ freeRunCntr\[1\] _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1972__A2 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1724__A2 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2429_ _1432_ _1436_ _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_29_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1660__A1 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1858__B _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1715__A2 _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2912__A1 _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2140__A2 _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1651__A1 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1800_ _0763_ _0849_ _1598_ _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2780_ _0284_ _0310_ _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1731_ _0778_ _0779_ _0780_ _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_11_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1662_ _0439_ _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__1954__A2 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2903__A1 _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3194_ _1117_ _0735_ _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2214_ _1220_ _1260_ _1261_ _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2145_ _1122_ _1192_ _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_4
XFILLER_19_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2076_ _1115_ sigRom.address\[0\] _1117_ _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1890__A1 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2978_ _0972_ _1151_ _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1929_ _0745_ _0977_ _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1860__C _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1881__A1 freeRunCntr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1881__B2 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2189__A2 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2361__A2 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2113__A2 _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1872__A1 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2901_ _1172_ _1581_ _1582_ _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_43_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2832_ _0318_ _1317_ _1318_ _0812_ _1252_ _0472_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_4
XFILLER_31_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2763_ _0259_ _0260_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1714_ _0252_ _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2694_ _1351_ _1353_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3129__A1 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1645_ _1554_ _0065_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_58_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3177_ _0955_ _1345_ _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1863__A1 _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2128_ _1122_ _1125_ _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2059_ _0560_ _1025_ _1007_ freeRunCntr\[10\] _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1615__A1 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2040__A1 freeRunCntr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2032__B _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1871__B _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1854__A1 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2031__A1 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2031__B2 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2334__A2 _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3100_ _0647_ _0650_ _0646_ _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3031_ freeRunCntr\[14\] _0584_ _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3204__D _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2098__A1 _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2815_ _1533_ _0217_ _0339_ _0350_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_31_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2746_ _0243_ _0244_ _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2022__B2 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2677_ _0129_ _0134_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1628_ _1565_ _1598_ _0065_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2325__A2 _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3229_ _0020_ net11 clknet_2_2__leaf_clk freeRunCntr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__1836__A1 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2013__A1 _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1827__A1 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1776__B _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2600_ _1056_ _0113_ _0114_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2531_ _1403_ _1385_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1763__B1 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2462_ _0965_ _1171_ _1527_ _1528_ _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_2393_ _1451_ _1452_ _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3014_ _0543_ _0542_ _0569_ _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1818__A1 _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2626__I _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2243__A1 _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2729_ _0251_ _0256_ _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_59_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1809__A1 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2785__A2 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1745__B1 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2220__B _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1760__A3 _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3210__CLK clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2473__A1 _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1962_ _0787_ _0979_ _0806_ _0800_ _0098_ _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_1893_ _0941_ _0942_ _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_5_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2514_ _1579_ _1580_ _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2445_ _1504_ _1508_ _1509_ _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2376_ _0395_ _1096_ _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_71_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2216__A1 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2767__A2 _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3233__CLK clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2040__B _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2207__A1 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3097__I _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2230_ _1259_ _1271_ _1277_ _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2161_ _1199_ _1200_ _1198_ _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2092_ sigRom.address\[0\] _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_65_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2994_ _0467_ _0419_ _0468_ _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1945_ _0745_ _0992_ _0993_ _1499_ _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1876_ _0417_ _0925_ _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_2428_ _0770_ _1214_ _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2359_ _1204_ _1205_ _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2437__A1 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1660__A2 csTable.address\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1948__B1 _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1874__B _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2428__A1 _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2979__A2 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1651__A2 csTable.address\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2600__A1 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1730_ _1422_ _0761_ _1444_ _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1661_ _0428_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3207__D _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3193_ _0736_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2213_ _1222_ _1226_ _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2144_ sigRom.address\[0\] _1191_ _1123_ _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2419__A1 _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2075_ _1118_ _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__1959__B _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3092__A1 freeRunCntr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2977_ _0431_ _0429_ _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2198__A3 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1928_ _0849_ _0841_ _0842_ _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1859_ _0651_ _0707_ _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1713__I _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3083__A1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1872__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3074__A1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2900_ _1533_ _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2831_ _0323_ _0324_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2762_ _0258_ _0264_ _0292_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1713_ _1477_ _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2693_ _0209_ _0212_ _0216_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1644_ _1521_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3176_ _0417_ _0720_ _0723_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1863__A2 _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2127_ _0395_ _1016_ _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__1689__B _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2058_ freeRunCntr\[8\] _1017_ _1025_ _0560_ _1106_ _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2112__I0 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1615__A2 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2040__A2 _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2032__C _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1871__C _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1854__A2 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2031__A2 _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1618__I _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1781__C _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3030_ _0577_ _0579_ _0583_ _0587_ _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__2098__A2 _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1845__A2 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3047__A1 freeRunCntr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output6_I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2814_ _0346_ _0349_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2745_ _1350_ _1365_ _0273_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_11_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2676_ _0194_ _0196_ _0198_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__1781__A1 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1972__B _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1627_ _0054_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__2325__A3 _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3228_ _0019_ net11 clknet_2_2__leaf_clk freeRunCntr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_39_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3159_ _0710_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2094__I _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1866__C _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2013__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1772__A1 _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1882__B _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1827__A2 _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3029__A1 freeRunCntr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3029__B2 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2004__A2 _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2530_ _1121_ _0037_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1763__A1 freeRunCntr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1763__B2 freeRunCntr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2461_ _1525_ _1526_ _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2392_ _1442_ _1443_ _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_3013_ _0528_ _0541_ _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_36_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1818__A2 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2243__A2 _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2728_ _0254_ _0255_ _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1754__A1 _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2659_ _1432_ _0171_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_59_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1877__B _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1993__A1 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1745__B2 _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1745__A1 _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2170__A1 _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2473__A2 _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1961_ _0764_ _0988_ _1009_ _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1892_ _0936_ _0940_ _1367_ _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__1984__A1 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1736__A1 _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2513_ _1579_ _1580_ _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2444_ _1159_ _1458_ _1505_ _1507_ _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_2375_ _0955_ _1087_ _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2216__A2 _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1975__A1 _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1727__A1 _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2040__C freeRunCntr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2152__A1 _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1966__A1 _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2391__A1 _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2694__A2 _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2160_ _1198_ _1199_ _1200_ _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2091_ _0417_ _0307_ _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1654__B1 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2993_ _0441_ _0546_ _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_9_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1944_ _0902_ _0889_ _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1957__A1 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1875_ _0670_ _0919_ _0923_ _0924_ _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__1709__A1 _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2382__A1 _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1980__B _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2427_ _1487_ _1490_ _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_69_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2134__A1 _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2358_ _1412_ _1413_ _1414_ _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2289_ _1290_ _1292_ _1291_ _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2437__A2 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1948__B2 freeRunCntr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1948__A1 freeRunCntr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2125__A1 _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2428__A2 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1939__A1 _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2061__B1 _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1660_ _1345_ csTable.address\[5\] _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2116__A1 _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3192_ _1117_ _0735_ _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2212_ _1222_ _1226_ _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2143_ _1115_ _1117_ _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2074_ _1115_ sigRom.address\[0\] _1117_ _1118_ _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_34_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2136__B _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3223__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2976_ _0424_ _0427_ _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout10_I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2052__B1 _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1927_ _0131_ _0902_ _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1858_ _0263_ _0742_ _0571_ _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1789_ _0153_ _0142_ _0631_ _1521_ _0087_ _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__2355__A1 _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1866__B1 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3083__A2 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2594__A1 _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2346__A1 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3074__A2 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2830_ _0366_ _0367_ _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_31_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2761_ _0257_ _0265_ _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2692_ _0213_ _0215_ _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1712_ _1598_ _0761_ _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1643_ _1510_ _0109_ _0219_ _0230_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_6_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2888__A2 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3175_ _0955_ _0720_ _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2126_ _1132_ _1133_ _1173_ _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2057_ _0946_ _1035_ _1104_ _1105_ _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2112__I1 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2959_ _0312_ _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2576__A1 _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2328__A1 _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2500__A1 _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2567__A1 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3220__RN net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2813_ _0347_ _0348_ _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_31_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2558__A1 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2744_ _1347_ _1366_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2675_ _0159_ _0160_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1626_ _0043_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__3211__RN net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3227_ _0018_ net11 clknet_2_2__leaf_clk freeRunCntr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_39_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3158_ _0708_ _0709_ _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2109_ _0768_ _0769_ _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_54_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3089_ _0601_ _0594_ freeRunCntr\[8\] _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2013__A3 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1772__A2 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3202__RN net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2485__B1 _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2788__A1 _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1763__A2 _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2460_ _1525_ _1526_ _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_5_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2391_ _1121_ _1449_ _1450_ _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3012_ _0539_ _0567_ _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2243__A3 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1983__B _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2727_ _0235_ _1357_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1754__A2 _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2658_ _0178_ _0177_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1609_ csTable.address\[0\] _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2589_ _0036_ _0059_ _0060_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XANTENNA__2306__I1 _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1809__A3 _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1690__A1 _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1877__C freeRunCntr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3195__A1 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1745__A2 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2170__A2 _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1787__C _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1960_ _0252_ _1008_ _0329_ _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1891_ _1367_ _0936_ _0940_ _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_41_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2512_ _1172_ _1581_ _1582_ _1583_ _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_2443_ _1159_ _1505_ _1507_ _1458_ _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2374_ _1056_ _1171_ _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_68_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2161__A2 _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3177__A1 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1727__A2 _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2152__A2 _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3101__A1 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1663__A1 _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1888__B _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2207__A3 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1966__A2 _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2143__A2 _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1642__I _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2090_ _1120_ _1136_ _1137_ _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1654__A1 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2992_ _0545_ _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1943_ _0800_ _0754_ _0991_ _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1874_ _0651_ _0867_ _0775_ _0750_ _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__1709__A2 _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2906__A1 _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2426_ _1132_ _1489_ _1487_ _1445_ _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2357_ _1409_ _1410_ _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2288_ _1299_ _1308_ _1337_ _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1645__A1 _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1948__A2 _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1890__C _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2125__A2 _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1884__A1 _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1636__A1 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1939__A2 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2061__A1 freeRunCntr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2061__B2 freeRunCntr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1637__I _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2349__C1 _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2116__A2 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3191_ _1140_ _0733_ _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2211_ _1172_ _1179_ _1258_ _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2142_ _0911_ _0912_ _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__1875__A1 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2073_ _1007_ _1119_ _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_19_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2975_ _0432_ _0429_ _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2931__I freeRunCntr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2052__A1 freeRunCntr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1926_ freeRunCntr\[16\] _0972_ _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2052__B2 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2152__B _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1857_ _0805_ _0906_ _0775_ _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1788_ _0120_ _0054_ _0804_ _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2107__A2 _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2409_ _1469_ _1470_ _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1866__A1 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1866__B2 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2291__A1 _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1885__C _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2043__A1 _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2594__A2 _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2997__B _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2346__A2 _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2034__A1 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2760_ _0254_ _0255_ _0290_ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2691_ _1374_ _0214_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1711_ _1466_ _1411_ _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_1642_ _0098_ _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1848__A1 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3174_ _0721_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2125_ _0996_ _1119_ _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2056_ freeRunCntr\[8\] _1017_ _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2273__A1 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2958_ _0479_ _0484_ _0504_ _0507_ _0508_ _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__2025__A1 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1909_ _0857_ _0219_ _0957_ _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2576__A2 _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2889_ _0431_ _0432_ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1839__A1 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2500__A2 _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2016__A1 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1775__B1 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3213__CLK clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2007__A1 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2812_ _0269_ _0279_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2743_ _0271_ _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2674_ _0126_ _0195_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1625_ _1334_ _1411_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3226_ _0017_ net10 clknet_2_2__leaf_clk csTable.address\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3157_ _1433_ freeRunCntr\[17\] _0703_ _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2494__A1 _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2108_ _0768_ _0769_ _1141_ _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_3088_ _0644_ _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2039_ _0395_ _1087_ _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_35_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2485__A1 _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2237__A1 _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2788__A2 _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2390_ _1447_ _1448_ _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3011_ _0562_ _0566_ _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_67_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2476__A1 _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1987__B1 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1983__C _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2726_ _1172_ _0253_ _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2657_ _0176_ _0169_ _0174_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1608_ _1334_ _1411_ _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_4
X_2588_ _0100_ _0101_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_47_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3209_ _0031_ net9 clknet_2_1__leaf_clk freeRunCntr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1690__A2 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2219__A1 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2630__A1 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1890_ _0851_ _0938_ _0939_ _0750_ _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_2511_ _1263_ _1525_ _1526_ _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2442_ _0836_ _1248_ _1252_ _0913_ _1506_ _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_2373_ _1375_ _1430_ _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2697__A1 _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2449__A1 _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3177__A2 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1727__A3 _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2709_ _0799_ _0809_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1663__A2 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1966__A3 _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1654__A2 _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2991_ _0542_ _0544_ _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_61_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2603__A1 _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1942_ _0131_ _0804_ _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1873_ _0651_ _0921_ _0922_ _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_6_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1833__I freeRunCntr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2425_ _1097_ _1171_ _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2356_ _1395_ _1393_ _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2287_ _1302_ _1336_ _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1989__B _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1645__A2 _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1884__A2 _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2833__A1 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1636__A2 _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2061__A2 _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2349__B1 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2349__C2 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2210_ _1174_ _1178_ _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3190_ _0734_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2141_ _1147_ _1188_ _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_4
XANTENNA__1875__A2 _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2072_ _0985_ _1119_ _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__3077__A1 freeRunCntr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2974_ _0474_ _0524_ _0525_ _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1925_ _0966_ _0970_ _0973_ _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2052__A2 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1856_ _0698_ _0065_ _0631_ _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1787_ _0698_ _0780_ _0800_ _0806_ _0087_ _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__1991__C _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2408_ _1409_ _1410_ _1413_ _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__1866__A2 _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2595__S _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2339_ _1088_ _1164_ _1213_ _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3068__A1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2815__A1 _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2291__A2 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2043__A2 _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3059__A1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2034__A2 _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2253__B _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2690_ _1376_ _1429_ _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1710_ _0631_ _0759_ _0651_ _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1641_ _0131_ _0164_ _0197_ _0208_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__1793__A1 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input5_I rst vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3173_ _1345_ _0720_ _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2124_ _0962_ _1171_ _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_39_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2055_ freeRunCntr\[6\] _1045_ _1103_ _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2957_ _0882_ _0506_ _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2025__A2 _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2888_ _0398_ _0400_ _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1908_ _0956_ _0351_ _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1784__A1 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2981__B1 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1839_ _0428_ _0285_ _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1839__A2 _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1775__B2 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1775__A1 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2007__A2 _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2811_ _0343_ _0344_ _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2742_ _1335_ _1346_ _0270_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1766__A1 freeRunCntr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2673_ _0122_ _0125_ _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1624_ _1587_ _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2191__A1 _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3225_ _0016_ net11 clknet_2_2__leaf_clk csTable.address\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3156_ _1466_ _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3087_ _0946_ _0640_ _0643_ _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_27_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2107_ _1154_ _1142_ _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2038_ _0670_ _1082_ _1084_ _0745_ _1086_ _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_54_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1757__A1 _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2485__A2 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1996__A1 _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1748__A1 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2173__A1 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1920__A1 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1661__I _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3010_ _0563_ _0564_ _0565_ _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_36_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1987__A1 _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1739__A1 _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2725_ _0985_ _1305_ _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2656_ _0169_ _0174_ _0176_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1607_ csTable.address\[2\] _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_2587_ _0038_ _0057_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1911__A1 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3208_ _0030_ net10 clknet_2_3__leaf_clk freeRunCntr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_3139_ _0593_ _0639_ _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_27_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1690__A3 _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2219__A2 _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1978__A1 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3203__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1666__B1 _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1969__A1 _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2630__A2 _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2510_ _1579_ _1580_ _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2394__A1 _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2441_ _0898_ _0899_ _1142_ _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_45_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2372_ _1376_ _1429_ _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2449__A2 _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3226__CLK clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2708_ _1359_ _1360_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2385__A1 _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2639_ _0155_ _0157_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2137__A1 _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2860__A2 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1820__B1 _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2376__A1 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2915__A3 _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2300__A1 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2990_ _0421_ _0435_ _0543_ _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1941_ _0602_ _0891_ _0987_ _0989_ _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1872_ _0730_ _0738_ _0757_ _0854_ _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_9_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2424_ _1435_ _1035_ _1289_ _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2355_ _1409_ _1410_ _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2286_ _1307_ _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_49_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3095__A2 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2530__A1 _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2833__A2 _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2597__A1 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2349__B2 _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3010__A2 _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2521__A1 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2140_ _1115_ _1117_ _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2071_ _1116_ _1117_ _1118_ _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_38_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2973_ freeRunCntr\[8\] _0512_ _0513_ _0477_ _0560_ _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__2037__B1 _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1924_ freeRunCntr\[16\] _0972_ _0969_ freeRunCntr\[15\] _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1855_ _0903_ _0904_ _0670_ _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1786_ _1367_ _0835_ _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_4
XFILLER_69_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2512__A1 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2407_ _1464_ _1467_ _1468_ _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2338_ _1390_ _1391_ _1388_ _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_57_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2269_ _1123_ _1186_ _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_4
XFILLER_29_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3068__A2 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2815__A2 _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2043__A3 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3232__RN net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2534__B _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1793__A2 _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1640_ _1554_ _0054_ _0120_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__3223__RN net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3172_ csTable.address\[5\] _0718_ _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2123_ _1119_ _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__1848__A3 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2054_ _1101_ _1102_ _1035_ _0946_ _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2258__B1 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2956_ _0882_ _0506_ _0491_ freeRunCntr\[4\] _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2887_ _0396_ _0430_ _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1907_ _0783_ _0849_ _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2981__A1 _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2981__B2 _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1838_ _0886_ _0887_ _0450_ _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1769_ _0771_ _0772_ _0818_ _0816_ _0813_ _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__3214__RN net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1775__A2 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2972__A1 _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput6 net6 qcomplex vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2724__A1 _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3205__RN net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1659__I _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2810_ _0341_ _0345_ _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2741_ _1338_ _1344_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1766__A2 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2672_ _0159_ _0160_ _0191_ _0193_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1623_ _1576_ _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__2191__A2 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3224_ _0015_ net11 clknet_2_2__leaf_clk csTable.address\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
.ends

